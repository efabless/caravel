magic
tech sky130A
magscale 1 2
timestamp 1666028836
<< viali >>
rect 3525 13481 3559 13515
rect 7205 13481 7239 13515
rect 6101 13413 6135 13447
rect 7665 13413 7699 13447
rect 8677 13413 8711 13447
rect 9137 13413 9171 13447
rect 6929 13345 6963 13379
rect 9505 13345 9539 13379
rect 11529 13345 11563 13379
rect 12725 13345 12759 13379
rect 1869 13277 1903 13311
rect 2237 13277 2271 13311
rect 3157 13277 3191 13311
rect 3433 13277 3467 13311
rect 4353 13277 4387 13311
rect 4905 13277 4939 13311
rect 5089 13277 5123 13311
rect 5549 13277 5583 13311
rect 6469 13277 6503 13311
rect 7021 13277 7055 13311
rect 7481 13277 7515 13311
rect 7797 13277 7831 13311
rect 8217 13277 8251 13311
rect 8309 13277 8343 13311
rect 8769 13277 8803 13311
rect 8953 13277 8987 13311
rect 9413 13277 9447 13311
rect 9597 13277 9631 13311
rect 10057 13277 10091 13311
rect 10609 13277 10643 13311
rect 10793 13277 10827 13311
rect 11345 13277 11379 13311
rect 12081 13277 12115 13311
rect 12173 13277 12207 13311
rect 12817 13277 12851 13311
rect 13369 13277 13403 13311
rect 1593 13209 1627 13243
rect 2053 13209 2087 13243
rect 2697 13209 2731 13243
rect 2789 13209 2823 13243
rect 2973 13209 3007 13243
rect 4077 13209 4111 13243
rect 4445 13209 4479 13243
rect 5641 13209 5675 13243
rect 6653 13209 6687 13243
rect 7297 13209 7331 13243
rect 7941 13209 7975 13243
rect 8033 13209 8067 13243
rect 10333 13209 10367 13243
rect 10885 13209 10919 13243
rect 11621 13209 11655 13243
rect 12633 13209 12667 13243
rect 13277 13209 13311 13243
rect 1409 13141 1443 13175
rect 1685 13141 1719 13175
rect 3341 13141 3375 13175
rect 4169 13141 4203 13175
rect 8493 13141 8527 13175
rect 9321 13141 9355 13175
rect 10425 13141 10459 13175
rect 13553 13141 13587 13175
rect 1593 12937 1627 12971
rect 11161 12937 11195 12971
rect 13369 12937 13403 12971
rect 4445 12869 4479 12903
rect 6193 12869 6227 12903
rect 8401 12869 8435 12903
rect 10057 12869 10091 12903
rect 10425 12869 10459 12903
rect 13093 12869 13127 12903
rect 13277 12869 13311 12903
rect 1685 12801 1719 12835
rect 2605 12801 2639 12835
rect 2789 12801 2823 12835
rect 3709 12801 3743 12835
rect 4629 12801 4663 12835
rect 5549 12801 5583 12835
rect 6377 12801 6411 12835
rect 7573 12801 7607 12835
rect 8217 12801 8251 12835
rect 8493 12801 8527 12835
rect 9413 12801 9447 12835
rect 10149 12801 10183 12835
rect 11069 12801 11103 12835
rect 11345 12801 11379 12835
rect 11529 12801 11563 12835
rect 12449 12801 12483 12835
rect 1777 12733 1811 12767
rect 2329 12733 2363 12767
rect 2237 12665 2271 12699
rect 2421 12665 2455 12699
rect 4261 12665 4295 12699
rect 7665 12665 7699 12699
rect 4077 12393 4111 12427
rect 5273 12393 5307 12427
rect 8769 12393 8803 12427
rect 10517 12393 10551 12427
rect 2789 12325 2823 12359
rect 3433 12325 3467 12359
rect 6837 12325 6871 12359
rect 9045 12325 9079 12359
rect 10149 12325 10183 12359
rect 6929 12257 6963 12291
rect 8585 12257 8619 12291
rect 9689 12257 9723 12291
rect 10241 12257 10275 12291
rect 1501 12189 1535 12223
rect 2605 12189 2639 12223
rect 3249 12189 3283 12223
rect 3893 12189 3927 12223
rect 4169 12189 4203 12223
rect 4813 12189 4847 12223
rect 5181 12189 5215 12223
rect 6377 12189 6411 12223
rect 7021 12189 7055 12223
rect 7941 12189 7975 12223
rect 8033 12189 8067 12223
rect 9224 12189 9258 12223
rect 9413 12189 9447 12223
rect 9597 12189 9631 12223
rect 10333 12189 10367 12223
rect 10517 12189 10551 12223
rect 10977 12189 11011 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 11989 12189 12023 12223
rect 12541 12189 12575 12223
rect 13185 12189 13219 12223
rect 5089 12121 5123 12155
rect 5457 12121 5491 12155
rect 5641 12121 5675 12155
rect 5825 12121 5859 12155
rect 5917 12121 5951 12155
rect 6101 12121 6135 12155
rect 6285 12121 6319 12155
rect 7297 12121 7331 12155
rect 8493 12121 8527 12155
rect 9321 12121 9355 12155
rect 12357 12121 12391 12155
rect 13461 12121 13495 12155
rect 3617 12053 3651 12087
rect 10701 12053 10735 12087
rect 12173 12053 12207 12087
rect 6469 11849 6503 11883
rect 7389 11849 7423 11883
rect 8125 11849 8159 11883
rect 10885 11849 10919 11883
rect 2237 11781 2271 11815
rect 2513 11781 2547 11815
rect 2605 11781 2639 11815
rect 4629 11781 4663 11815
rect 6009 11781 6043 11815
rect 10241 11781 10275 11815
rect 1593 11713 1627 11747
rect 2789 11713 2823 11747
rect 3065 11713 3099 11747
rect 3893 11713 3927 11747
rect 3985 11713 4019 11747
rect 4485 11713 4519 11747
rect 4721 11713 4755 11747
rect 4905 11713 4939 11747
rect 5268 11713 5302 11747
rect 5365 11713 5399 11747
rect 5457 11713 5491 11747
rect 5641 11713 5675 11747
rect 6193 11713 6227 11747
rect 6653 11713 6687 11747
rect 6837 11713 6871 11747
rect 6929 11713 6963 11747
rect 7073 11713 7107 11747
rect 7757 11713 7791 11747
rect 8013 11713 8047 11747
rect 8493 11713 8527 11747
rect 9229 11713 9263 11747
rect 9413 11713 9447 11747
rect 9505 11713 9539 11747
rect 9781 11713 9815 11747
rect 10057 11713 10091 11747
rect 10517 11713 10551 11747
rect 10773 11713 10807 11747
rect 11345 11713 11379 11747
rect 11713 11713 11747 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 13461 11713 13495 11747
rect 3525 11645 3559 11679
rect 3617 11645 3651 11679
rect 4077 11645 4111 11679
rect 8217 11645 8251 11679
rect 8309 11645 8343 11679
rect 8953 11645 8987 11679
rect 9321 11645 9355 11679
rect 10977 11645 11011 11679
rect 11069 11645 11103 11679
rect 1409 11577 1443 11611
rect 4353 11577 4387 11611
rect 10333 11577 10367 11611
rect 13277 11577 13311 11611
rect 3709 11509 3743 11543
rect 5089 11509 5123 11543
rect 5917 11509 5951 11543
rect 7205 11509 7239 11543
rect 7573 11509 7607 11543
rect 8585 11509 8619 11543
rect 9965 11509 9999 11543
rect 11253 11509 11287 11543
rect 11621 11509 11655 11543
rect 4905 11305 4939 11339
rect 5549 11305 5583 11339
rect 6469 11305 6503 11339
rect 7481 11305 7515 11339
rect 7665 11305 7699 11339
rect 9137 11305 9171 11339
rect 10793 11305 10827 11339
rect 11529 11305 11563 11339
rect 1869 11237 1903 11271
rect 5733 11237 5767 11271
rect 7297 11237 7331 11271
rect 12449 11237 12483 11271
rect 3065 11169 3099 11203
rect 3617 11169 3651 11203
rect 8677 11169 8711 11203
rect 11345 11169 11379 11203
rect 2329 11101 2363 11135
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 3525 11101 3559 11135
rect 3985 11101 4019 11135
rect 4721 11101 4755 11135
rect 4997 11101 5031 11135
rect 5370 11101 5404 11135
rect 5917 11101 5951 11135
rect 6290 11101 6324 11135
rect 6653 11101 6687 11135
rect 6837 11101 6871 11135
rect 6954 11079 6988 11113
rect 7055 11079 7089 11113
rect 7832 11101 7866 11135
rect 7981 11101 8015 11135
rect 8125 11101 8159 11135
rect 8401 11101 8435 11135
rect 9413 11101 9447 11135
rect 10241 11101 10275 11135
rect 10517 11101 10551 11135
rect 11049 11101 11083 11135
rect 11897 11101 11931 11135
rect 12173 11101 12207 11135
rect 12317 11101 12351 11135
rect 12633 11101 12667 11135
rect 13369 11101 13403 11135
rect 1593 11033 1627 11067
rect 1777 11033 1811 11067
rect 2881 11033 2915 11067
rect 3801 11033 3835 11067
rect 5181 11033 5215 11067
rect 5273 11033 5307 11067
rect 6101 11033 6135 11067
rect 6193 11033 6227 11067
rect 8217 11033 8251 11067
rect 8769 11033 8803 11067
rect 8953 11033 8987 11067
rect 9505 11033 9539 11067
rect 9689 11033 9723 11067
rect 9873 11033 9907 11067
rect 10057 11033 10091 11067
rect 10793 11033 10827 11067
rect 11621 11033 11655 11067
rect 11805 11033 11839 11067
rect 12081 11033 12115 11067
rect 13093 11033 13127 11067
rect 13185 11033 13219 11067
rect 1685 10965 1719 10999
rect 2513 10965 2547 10999
rect 9137 10965 9171 10999
rect 10425 10965 10459 10999
rect 11161 10965 11195 10999
rect 11253 10965 11287 10999
rect 13461 10965 13495 10999
rect 6561 10761 6595 10795
rect 8401 10761 8435 10795
rect 10149 10761 10183 10795
rect 3433 10693 3467 10727
rect 4261 10693 4295 10727
rect 5273 10693 5307 10727
rect 7205 10693 7239 10727
rect 9953 10693 9987 10727
rect 10977 10693 11011 10727
rect 1409 10625 1443 10659
rect 2697 10625 2731 10659
rect 3336 10625 3370 10659
rect 3525 10625 3559 10659
rect 3709 10625 3743 10659
rect 3985 10625 4019 10659
rect 4537 10625 4571 10659
rect 5181 10625 5215 10659
rect 5825 10625 5859 10659
rect 6193 10625 6227 10659
rect 6673 10625 6707 10659
rect 6929 10625 6963 10659
rect 7113 10625 7147 10659
rect 7849 10625 7883 10659
rect 7941 10625 7975 10659
rect 8567 10625 8601 10659
rect 8677 10625 8711 10659
rect 9137 10625 9171 10659
rect 9320 10625 9354 10659
rect 9689 10625 9723 10659
rect 10741 10625 10775 10659
rect 10885 10625 10919 10659
rect 11161 10625 11195 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 13369 10625 13403 10659
rect 5365 10557 5399 10591
rect 6377 10557 6411 10591
rect 6469 10557 6503 10591
rect 8217 10557 8251 10591
rect 8953 10557 8987 10591
rect 9413 10557 9447 10591
rect 9505 10557 9539 10591
rect 2697 10489 2731 10523
rect 3801 10489 3835 10523
rect 4169 10489 4203 10523
rect 8125 10489 8159 10523
rect 9873 10489 9907 10523
rect 10609 10489 10643 10523
rect 11253 10489 11287 10523
rect 13277 10489 13311 10523
rect 3157 10421 3191 10455
rect 6009 10421 6043 10455
rect 7297 10421 7331 10455
rect 7665 10421 7699 10455
rect 8861 10421 8895 10455
rect 10149 10421 10183 10455
rect 10333 10421 10367 10455
rect 11621 10421 11655 10455
rect 6469 10217 6503 10251
rect 9505 10217 9539 10251
rect 9873 10217 9907 10251
rect 13277 10217 13311 10251
rect 5089 10149 5123 10183
rect 5733 10149 5767 10183
rect 9045 10149 9079 10183
rect 11253 10149 11287 10183
rect 12541 10081 12575 10115
rect 13093 10081 13127 10115
rect 1501 10013 1535 10047
rect 1777 10013 1811 10047
rect 2697 10013 2731 10047
rect 2789 10013 2823 10047
rect 3341 10013 3375 10047
rect 3525 10013 3559 10047
rect 3801 10013 3835 10047
rect 4905 10013 4939 10047
rect 5641 10013 5675 10047
rect 5917 10013 5951 10047
rect 6193 10013 6227 10047
rect 6745 10013 6779 10047
rect 6929 10013 6963 10047
rect 7022 9991 7056 10025
rect 7147 10013 7181 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 8217 10013 8251 10047
rect 8401 10013 8435 10047
rect 8493 10013 8527 10047
rect 8585 10013 8619 10047
rect 8953 10013 8987 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 9965 10013 9999 10047
rect 10333 10013 10367 10047
rect 10701 10013 10735 10047
rect 10885 10013 10919 10047
rect 11121 10013 11155 10047
rect 11713 10013 11747 10047
rect 12449 10013 12483 10047
rect 13185 10013 13219 10047
rect 13369 10013 13403 10047
rect 1961 9945 1995 9979
rect 3065 9945 3099 9979
rect 6101 9945 6135 9979
rect 6469 9945 6503 9979
rect 6653 9945 6687 9979
rect 7389 9945 7423 9979
rect 8033 9945 8067 9979
rect 10149 9945 10183 9979
rect 10609 9945 10643 9979
rect 10977 9945 11011 9979
rect 11529 9945 11563 9979
rect 12633 9945 12667 9979
rect 1685 9877 1719 9911
rect 2973 9877 3007 9911
rect 3157 9877 3191 9911
rect 5457 9877 5491 9911
rect 7573 9877 7607 9911
rect 8769 9877 8803 9911
rect 10517 9877 10551 9911
rect 4629 9673 4663 9707
rect 4905 9673 4939 9707
rect 6009 9673 6043 9707
rect 7665 9673 7699 9707
rect 8125 9673 8159 9707
rect 8585 9673 8619 9707
rect 10057 9673 10091 9707
rect 1869 9605 1903 9639
rect 1961 9605 1995 9639
rect 3157 9605 3191 9639
rect 3801 9605 3835 9639
rect 4445 9605 4479 9639
rect 5181 9605 5215 9639
rect 6377 9605 6411 9639
rect 7297 9605 7331 9639
rect 7481 9605 7515 9639
rect 8309 9605 8343 9639
rect 9229 9605 9263 9639
rect 10885 9605 10919 9639
rect 11529 9605 11563 9639
rect 12357 9605 12391 9639
rect 1777 9537 1811 9571
rect 2513 9537 2547 9571
rect 2605 9537 2639 9571
rect 3341 9537 3375 9571
rect 3985 9537 4019 9571
rect 4997 9537 5031 9571
rect 5733 9537 5767 9571
rect 6193 9537 6227 9571
rect 6561 9537 6595 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 6963 9537 6997 9571
rect 7849 9537 7883 9571
rect 8401 9537 8435 9571
rect 8953 9537 8987 9571
rect 9321 9537 9355 9571
rect 9597 9537 9631 9571
rect 9827 9537 9861 9571
rect 9941 9537 9975 9571
rect 10241 9537 10275 9571
rect 10425 9537 10459 9571
rect 10701 9537 10735 9571
rect 11345 9537 11379 9571
rect 12081 9537 12115 9571
rect 12173 9537 12207 9571
rect 13369 9537 13403 9571
rect 1685 9469 1719 9503
rect 2421 9469 2455 9503
rect 3065 9469 3099 9503
rect 4537 9469 4571 9503
rect 9045 9469 9079 9503
rect 10149 9469 10183 9503
rect 12725 9469 12759 9503
rect 13277 9469 13311 9503
rect 3617 9401 3651 9435
rect 5273 9401 5307 9435
rect 7205 9401 7239 9435
rect 10333 9401 10367 9435
rect 11069 9401 11103 9435
rect 11621 9401 11655 9435
rect 13185 9401 13219 9435
rect 7481 9333 7515 9367
rect 8128 9333 8162 9367
rect 9413 9333 9447 9367
rect 11253 9333 11287 9367
rect 12449 9333 12483 9367
rect 13461 9333 13495 9367
rect 3617 9129 3651 9163
rect 6193 9129 6227 9163
rect 6469 9129 6503 9163
rect 7757 9129 7791 9163
rect 7941 9129 7975 9163
rect 9965 9129 9999 9163
rect 10241 9129 10275 9163
rect 12817 9129 12851 9163
rect 3893 9061 3927 9095
rect 6653 9061 6687 9095
rect 7021 9061 7055 9095
rect 9597 9061 9631 9095
rect 10701 9061 10735 9095
rect 11161 9061 11195 9095
rect 3801 8993 3835 9027
rect 4353 8993 4387 9027
rect 8493 8993 8527 9027
rect 13369 8993 13403 9027
rect 1777 8925 1811 8959
rect 1869 8925 1903 8959
rect 3341 8925 3375 8959
rect 4445 8925 4479 8959
rect 5089 8925 5123 8959
rect 6009 8925 6043 8959
rect 6285 8925 6319 8959
rect 7481 8925 7515 8959
rect 7941 8925 7975 8959
rect 8125 8925 8159 8959
rect 8401 8925 8435 8959
rect 8677 8925 8711 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9230 8925 9264 8959
rect 9338 8925 9372 8959
rect 9873 8925 9907 8959
rect 10057 8925 10091 8959
rect 10333 8925 10367 8959
rect 10793 8925 10827 8959
rect 10977 8925 11011 8959
rect 11345 8925 11379 8959
rect 12633 8925 12667 8959
rect 13001 8925 13035 8959
rect 3433 8857 3467 8891
rect 4905 8857 4939 8891
rect 4997 8857 5031 8891
rect 5273 8857 5307 8891
rect 6929 8857 6963 8891
rect 7205 8857 7239 8891
rect 7389 8857 7423 8891
rect 8769 8857 8803 8891
rect 10517 8857 10551 8891
rect 13277 8857 13311 8891
rect 1593 8789 1627 8823
rect 13185 8789 13219 8823
rect 2697 8585 2731 8619
rect 6561 8585 6595 8619
rect 7205 8585 7239 8619
rect 8493 8585 8527 8619
rect 9045 8585 9079 8619
rect 9781 8585 9815 8619
rect 10885 8585 10919 8619
rect 11253 8585 11287 8619
rect 2881 8517 2915 8551
rect 12311 8517 12345 8551
rect 1593 8449 1627 8483
rect 2789 8449 2823 8483
rect 3065 8449 3099 8483
rect 3801 8449 3835 8483
rect 4077 8449 4111 8483
rect 5549 8449 5583 8483
rect 5825 8449 5859 8483
rect 6009 8449 6043 8483
rect 6377 8449 6411 8483
rect 6745 8449 6779 8483
rect 7389 8449 7423 8483
rect 7665 8449 7699 8483
rect 7849 8449 7883 8483
rect 7941 8449 7975 8483
rect 8217 8449 8251 8483
rect 8309 8449 8343 8483
rect 8585 8449 8619 8483
rect 8769 8449 8803 8483
rect 9229 8449 9263 8483
rect 9321 8449 9355 8483
rect 9505 8449 9539 8483
rect 9597 8449 9631 8483
rect 10149 8449 10183 8483
rect 10695 8449 10729 8483
rect 10977 8449 11011 8483
rect 11069 8449 11103 8483
rect 11529 8449 11563 8483
rect 11897 8449 11931 8483
rect 12541 8449 12575 8483
rect 12633 8449 12667 8483
rect 13277 8449 13311 8483
rect 13553 8449 13587 8483
rect 1409 8381 1443 8415
rect 10057 8381 10091 8415
rect 10609 8381 10643 8415
rect 5365 8313 5399 8347
rect 6929 8313 6963 8347
rect 7757 8313 7791 8347
rect 11713 8313 11747 8347
rect 3893 8245 3927 8279
rect 10149 8245 10183 8279
rect 10333 8245 10367 8279
rect 10517 8245 10551 8279
rect 12265 8245 12299 8279
rect 3433 8041 3467 8075
rect 4353 8041 4387 8075
rect 7481 8041 7515 8075
rect 9413 8041 9447 8075
rect 9873 8041 9907 8075
rect 1685 7973 1719 8007
rect 8309 7973 8343 8007
rect 9045 7973 9079 8007
rect 11253 7973 11287 8007
rect 12173 7973 12207 8007
rect 7573 7905 7607 7939
rect 10241 7905 10275 7939
rect 11897 7905 11931 7939
rect 1593 7837 1627 7871
rect 1685 7837 1719 7871
rect 1961 7837 1995 7871
rect 2145 7837 2179 7871
rect 2329 7837 2363 7871
rect 2513 7837 2547 7871
rect 2973 7837 3007 7871
rect 3157 7837 3191 7871
rect 3249 7837 3283 7871
rect 3893 7837 3927 7871
rect 4077 7837 4111 7871
rect 4537 7837 4571 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 5457 7837 5491 7871
rect 5641 7837 5675 7871
rect 6101 7837 6135 7871
rect 6469 7837 6503 7871
rect 6929 7837 6963 7871
rect 8125 7837 8159 7871
rect 8401 7837 8435 7871
rect 8493 7837 8527 7871
rect 9229 7837 9263 7871
rect 9505 7837 9539 7871
rect 9597 7837 9631 7871
rect 9781 7837 9815 7871
rect 9873 7837 9907 7871
rect 10425 7837 10459 7871
rect 10793 7837 10827 7871
rect 10885 7837 10919 7871
rect 11713 7837 11747 7871
rect 12725 7837 12759 7871
rect 13001 7837 13035 7871
rect 1869 7769 1903 7803
rect 2789 7769 2823 7803
rect 4721 7769 4755 7803
rect 5733 7769 5767 7803
rect 7757 7769 7791 7803
rect 7941 7769 7975 7803
rect 11345 7769 11379 7803
rect 11989 7769 12023 7803
rect 12081 7769 12115 7803
rect 2605 7701 2639 7735
rect 4077 7701 4111 7735
rect 5181 7701 5215 7735
rect 5917 7701 5951 7735
rect 7297 7701 7331 7735
rect 8677 7701 8711 7735
rect 10057 7701 10091 7735
rect 10425 7701 10459 7735
rect 11253 7701 11287 7735
rect 13461 7701 13495 7735
rect 1777 7497 1811 7531
rect 2513 7497 2547 7531
rect 8861 7497 8895 7531
rect 9229 7497 9263 7531
rect 12265 7497 12299 7531
rect 1685 7429 1719 7463
rect 7941 7429 7975 7463
rect 9321 7429 9355 7463
rect 10977 7429 11011 7463
rect 4629 7361 4663 7395
rect 4905 7361 4939 7395
rect 5917 7361 5951 7395
rect 8493 7361 8527 7395
rect 8749 7361 8783 7395
rect 8953 7361 8987 7395
rect 9563 7361 9597 7395
rect 9689 7361 9723 7395
rect 9781 7361 9815 7395
rect 9965 7361 9999 7395
rect 10057 7361 10091 7395
rect 10333 7361 10367 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 11161 7361 11195 7395
rect 11345 7361 11379 7395
rect 11805 7361 11839 7395
rect 11897 7361 11931 7395
rect 12173 7361 12207 7395
rect 12909 7361 12943 7395
rect 1777 7293 1811 7327
rect 2697 7293 2731 7327
rect 2973 7293 3007 7327
rect 5181 7293 5215 7327
rect 8217 7293 8251 7327
rect 9045 7293 9079 7327
rect 12081 7293 12115 7327
rect 13001 7293 13035 7327
rect 4905 7225 4939 7259
rect 6469 7225 6503 7259
rect 10429 7225 10463 7259
rect 2237 7157 2271 7191
rect 4445 7157 4479 7191
rect 8309 7157 8343 7191
rect 11621 7157 11655 7191
rect 13553 7157 13587 7191
rect 1501 6953 1535 6987
rect 3525 6953 3559 6987
rect 12093 6953 12127 6987
rect 12633 6953 12667 6987
rect 3249 6817 3283 6851
rect 3985 6817 4019 6851
rect 6469 6817 6503 6851
rect 10609 6817 10643 6851
rect 12357 6817 12391 6851
rect 13185 6817 13219 6851
rect 3341 6749 3375 6783
rect 3801 6749 3835 6783
rect 6193 6749 6227 6783
rect 6377 6749 6411 6783
rect 9229 6749 9263 6783
rect 9689 6749 9723 6783
rect 10149 6749 10183 6783
rect 12633 6749 12667 6783
rect 12863 6749 12897 6783
rect 13461 6749 13495 6783
rect 2973 6681 3007 6715
rect 4261 6681 4295 6715
rect 6009 6681 6043 6715
rect 6745 6681 6779 6715
rect 5733 6613 5767 6647
rect 8217 6613 8251 6647
rect 10057 6613 10091 6647
rect 10333 6613 10367 6647
rect 13001 6613 13035 6647
rect 13093 6613 13127 6647
rect 13277 6613 13311 6647
rect 2697 6409 2731 6443
rect 4445 6409 4479 6443
rect 7021 6409 7055 6443
rect 7297 6409 7331 6443
rect 8769 6409 8803 6443
rect 9321 6409 9355 6443
rect 10885 6409 10919 6443
rect 11253 6409 11287 6443
rect 12173 6409 12207 6443
rect 13461 6409 13495 6443
rect 1869 6341 1903 6375
rect 3893 6341 3927 6375
rect 9873 6341 9907 6375
rect 12081 6341 12115 6375
rect 1685 6273 1719 6307
rect 2145 6273 2179 6307
rect 2513 6273 2547 6307
rect 2973 6273 3007 6307
rect 3249 6273 3283 6307
rect 4905 6273 4939 6307
rect 5549 6273 5583 6307
rect 5733 6273 5767 6307
rect 5917 6273 5951 6307
rect 6745 6273 6779 6307
rect 7021 6273 7055 6307
rect 7205 6273 7239 6307
rect 7389 6273 7423 6307
rect 7941 6273 7975 6307
rect 9319 6273 9353 6307
rect 10115 6273 10149 6307
rect 10609 6273 10643 6307
rect 10885 6273 10919 6307
rect 11069 6273 11103 6307
rect 11529 6273 11563 6307
rect 11713 6273 11747 6307
rect 12265 6273 12299 6307
rect 12449 6273 12483 6307
rect 12909 6273 12943 6307
rect 13093 6273 13127 6307
rect 13277 6273 13311 6307
rect 1501 6205 1535 6239
rect 1961 6205 1995 6239
rect 3893 6205 3927 6239
rect 3985 6205 4019 6239
rect 4629 6205 4663 6239
rect 4813 6205 4847 6239
rect 6101 6205 6135 6239
rect 7849 6205 7883 6239
rect 9781 6205 9815 6239
rect 10425 6205 10459 6239
rect 10517 6205 10551 6239
rect 3157 6137 3191 6171
rect 3433 6137 3467 6171
rect 9137 6137 9171 6171
rect 9689 6137 9723 6171
rect 12909 6137 12943 6171
rect 2329 6069 2363 6103
rect 4169 6069 4203 6103
rect 5089 6069 5123 6103
rect 5273 6069 5307 6103
rect 11805 6069 11839 6103
rect 12633 6069 12667 6103
rect 3341 5865 3375 5899
rect 7205 5865 7239 5899
rect 10774 5865 10808 5899
rect 8677 5797 8711 5831
rect 9045 5797 9079 5831
rect 1777 5729 1811 5763
rect 2789 5729 2823 5763
rect 4261 5729 4295 5763
rect 9505 5729 9539 5763
rect 13277 5729 13311 5763
rect 1501 5661 1535 5695
rect 1593 5661 1627 5695
rect 1961 5661 1995 5695
rect 2145 5661 2179 5695
rect 2237 5661 2271 5695
rect 2330 5661 2364 5695
rect 2697 5661 2731 5695
rect 2973 5661 3007 5695
rect 3525 5661 3559 5695
rect 4077 5661 4111 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 4905 5661 4939 5695
rect 4997 5661 5031 5695
rect 5090 5671 5124 5705
rect 5457 5661 5491 5695
rect 7389 5661 7423 5695
rect 7757 5661 7791 5695
rect 7941 5661 7975 5695
rect 8585 5661 8619 5695
rect 8769 5661 8803 5695
rect 9229 5661 9263 5695
rect 9781 5661 9815 5695
rect 10517 5661 10551 5695
rect 2605 5593 2639 5627
rect 5365 5593 5399 5627
rect 5733 5593 5767 5627
rect 8125 5593 8159 5627
rect 12449 5593 12483 5627
rect 3157 5525 3191 5559
rect 3893 5525 3927 5559
rect 4445 5525 4479 5559
rect 7573 5525 7607 5559
rect 10425 5525 10459 5559
rect 12265 5525 12299 5559
rect 1501 5321 1535 5355
rect 3157 5321 3191 5355
rect 3617 5321 3651 5355
rect 3709 5321 3743 5355
rect 9873 5321 9907 5355
rect 11603 5321 11637 5355
rect 12081 5321 12115 5355
rect 13461 5321 13495 5355
rect 1593 5253 1627 5287
rect 1961 5253 1995 5287
rect 3893 5253 3927 5287
rect 6561 5253 6595 5287
rect 9597 5253 9631 5287
rect 10701 5253 10735 5287
rect 12173 5253 12207 5287
rect 1777 5185 1811 5219
rect 2421 5185 2455 5219
rect 2973 5185 3007 5219
rect 3249 5185 3283 5219
rect 3525 5185 3559 5219
rect 5825 5185 5859 5219
rect 5917 5185 5951 5219
rect 6745 5185 6779 5219
rect 6929 5185 6963 5219
rect 9137 5185 9171 5219
rect 9505 5185 9539 5219
rect 9689 5185 9723 5219
rect 10517 5185 10551 5219
rect 10609 5185 10643 5219
rect 10885 5185 10919 5219
rect 11069 5185 11103 5219
rect 11897 5185 11931 5219
rect 12863 5185 12897 5219
rect 13001 5185 13035 5219
rect 13277 5185 13311 5219
rect 2053 5117 2087 5151
rect 2605 5117 2639 5151
rect 2789 5117 2823 5151
rect 5549 5117 5583 5151
rect 8861 5117 8895 5151
rect 10149 5117 10183 5151
rect 10333 5117 10367 5151
rect 12633 5117 12667 5151
rect 2145 5049 2179 5083
rect 3341 5049 3375 5083
rect 6101 5049 6135 5083
rect 9321 5049 9355 5083
rect 12725 5049 12759 5083
rect 4077 4981 4111 5015
rect 7389 4981 7423 5015
rect 1501 4777 1535 4811
rect 3341 4777 3375 4811
rect 5383 4777 5417 4811
rect 7573 4777 7607 4811
rect 9321 4777 9355 4811
rect 11253 4777 11287 4811
rect 2145 4709 2179 4743
rect 2973 4709 3007 4743
rect 7021 4709 7055 4743
rect 8033 4709 8067 4743
rect 12173 4709 12207 4743
rect 1869 4641 1903 4675
rect 4813 4641 4847 4675
rect 11621 4641 11655 4675
rect 1685 4573 1719 4607
rect 2145 4573 2179 4607
rect 2375 4573 2409 4607
rect 2697 4573 2731 4607
rect 2881 4573 2915 4607
rect 3065 4573 3099 4607
rect 3157 4573 3191 4607
rect 3801 4573 3835 4607
rect 4077 4573 4111 4607
rect 4445 4573 4479 4607
rect 5549 4573 5583 4607
rect 6377 4573 6411 4607
rect 6469 4573 6503 4607
rect 6653 4573 6687 4607
rect 7205 4573 7239 4607
rect 7389 4573 7423 4607
rect 7757 4573 7791 4607
rect 7941 4573 7975 4607
rect 8217 4573 8251 4607
rect 8401 4573 8435 4607
rect 9229 4573 9263 4607
rect 9321 4573 9355 4607
rect 9505 4573 9539 4607
rect 12817 4573 12851 4607
rect 13277 4573 13311 4607
rect 4353 4505 4387 4539
rect 4905 4505 4939 4539
rect 5089 4505 5123 4539
rect 5733 4505 5767 4539
rect 5917 4505 5951 4539
rect 6009 4505 6043 4539
rect 6193 4505 6227 4539
rect 8585 4505 8619 4539
rect 9781 4505 9815 4539
rect 11897 4505 11931 4539
rect 2513 4437 2547 4471
rect 2605 4437 2639 4471
rect 3617 4437 3651 4471
rect 4537 4437 4571 4471
rect 6561 4437 6595 4471
rect 11713 4437 11747 4471
rect 12449 4437 12483 4471
rect 2697 4233 2731 4267
rect 4629 4233 4663 4267
rect 6101 4233 6135 4267
rect 9321 4233 9355 4267
rect 9689 4233 9723 4267
rect 10517 4233 10551 4267
rect 11069 4233 11103 4267
rect 1501 4165 1535 4199
rect 7941 4165 7975 4199
rect 10333 4165 10367 4199
rect 1869 4097 1903 4131
rect 2145 4097 2179 4131
rect 2513 4097 2547 4131
rect 2789 4097 2823 4131
rect 3341 4097 3375 4131
rect 4169 4097 4203 4131
rect 4353 4097 4387 4131
rect 4629 4097 4663 4131
rect 4813 4097 4847 4131
rect 5273 4097 5307 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 8217 4097 8251 4131
rect 8769 4097 8803 4131
rect 9137 4097 9171 4131
rect 9873 4097 9907 4131
rect 10609 4097 10643 4131
rect 11069 4097 11103 4131
rect 11253 4097 11287 4131
rect 1961 4029 1995 4063
rect 2605 4029 2639 4063
rect 2881 4029 2915 4063
rect 5457 4029 5491 4063
rect 6193 4029 6227 4063
rect 8677 4029 8711 4063
rect 11529 4029 11563 4063
rect 11805 4029 11839 4063
rect 3157 3961 3191 3995
rect 6469 3961 6503 3995
rect 10057 3961 10091 3995
rect 13277 3961 13311 3995
rect 2973 3893 3007 3927
rect 5089 3893 5123 3927
rect 9137 3893 9171 3927
rect 1869 3689 1903 3723
rect 2053 3689 2087 3723
rect 3249 3689 3283 3723
rect 3525 3689 3559 3723
rect 3985 3689 4019 3723
rect 5089 3689 5123 3723
rect 5273 3689 5307 3723
rect 6377 3689 6411 3723
rect 9965 3689 9999 3723
rect 10149 3689 10183 3723
rect 12541 3689 12575 3723
rect 2329 3621 2363 3655
rect 5917 3621 5951 3655
rect 6193 3621 6227 3655
rect 9045 3621 9079 3655
rect 13185 3621 13219 3655
rect 1593 3553 1627 3587
rect 2881 3553 2915 3587
rect 5457 3553 5491 3587
rect 6929 3553 6963 3587
rect 10517 3553 10551 3587
rect 1685 3485 1719 3519
rect 1869 3485 1903 3519
rect 2513 3485 2547 3519
rect 2789 3485 2823 3519
rect 3249 3485 3283 3519
rect 4169 3485 4203 3519
rect 4261 3485 4295 3519
rect 4445 3485 4479 3519
rect 4537 3485 4571 3519
rect 4905 3485 4939 3519
rect 5641 3485 5675 3519
rect 6009 3485 6043 3519
rect 6653 3485 6687 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 7389 3485 7423 3519
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 9321 3485 9355 3519
rect 12909 3485 12943 3519
rect 13093 3485 13127 3519
rect 4629 3417 4663 3451
rect 6561 3417 6595 3451
rect 7573 3417 7607 3451
rect 7757 3417 7791 3451
rect 8769 3417 8803 3451
rect 9597 3417 9631 3451
rect 10149 3417 10183 3451
rect 10333 3417 10367 3451
rect 10793 3417 10827 3451
rect 12633 3417 12667 3451
rect 12817 3417 12851 3451
rect 2697 3349 2731 3383
rect 3065 3349 3099 3383
rect 4721 3349 4755 3383
rect 6377 3349 6411 3383
rect 7941 3349 7975 3383
rect 9505 3349 9539 3383
rect 12265 3349 12299 3383
rect 1869 3145 1903 3179
rect 3341 3145 3375 3179
rect 5089 3145 5123 3179
rect 6561 3145 6595 3179
rect 7389 3145 7423 3179
rect 9781 3145 9815 3179
rect 13461 3145 13495 3179
rect 2789 3077 2823 3111
rect 3801 3077 3835 3111
rect 7573 3077 7607 3111
rect 8309 3077 8343 3111
rect 10333 3077 10367 3111
rect 10517 3077 10551 3111
rect 11161 3077 11195 3111
rect 11897 3077 11931 3111
rect 12081 3077 12115 3111
rect 1593 3009 1627 3043
rect 1685 3009 1719 3043
rect 2329 3009 2363 3043
rect 2421 3009 2455 3043
rect 2973 3009 3007 3043
rect 3157 3009 3191 3043
rect 3525 3009 3559 3043
rect 4629 3009 4663 3043
rect 4813 3009 4847 3043
rect 5089 3009 5123 3043
rect 5181 3009 5215 3043
rect 5457 3009 5491 3043
rect 5733 3009 5767 3043
rect 6009 3009 6043 3043
rect 6561 3009 6595 3043
rect 6929 3009 6963 3043
rect 7113 3009 7147 3043
rect 7205 3009 7239 3043
rect 7665 3009 7699 3043
rect 7849 3009 7883 3043
rect 10977 3009 11011 3043
rect 11529 3009 11563 3043
rect 11713 3009 11747 3043
rect 13277 3009 13311 3043
rect 2145 2941 2179 2975
rect 2697 2941 2731 2975
rect 3709 2941 3743 2975
rect 5641 2941 5675 2975
rect 6377 2941 6411 2975
rect 8033 2941 8067 2975
rect 10609 2941 10643 2975
rect 12909 2941 12943 2975
rect 2605 2873 2639 2907
rect 10793 2873 10827 2907
rect 10057 2805 10091 2839
rect 5089 2601 5123 2635
rect 7757 2601 7791 2635
rect 10701 2601 10735 2635
rect 4077 2465 4111 2499
rect 4813 2465 4847 2499
rect 5372 2465 5406 2499
rect 5641 2465 5675 2499
rect 7941 2465 7975 2499
rect 8953 2465 8987 2499
rect 12725 2465 12759 2499
rect 3249 2397 3283 2431
rect 3433 2397 3467 2431
rect 3525 2397 3559 2431
rect 5273 2397 5307 2431
rect 7573 2397 7607 2431
rect 7757 2397 7791 2431
rect 8033 2397 8067 2431
rect 8309 2397 8343 2431
rect 8401 2397 8435 2431
rect 8677 2397 8711 2431
rect 12817 2397 12851 2431
rect 13093 2397 13127 2431
rect 3157 2329 3191 2363
rect 7297 2329 7331 2363
rect 9229 2329 9263 2363
rect 12449 2329 12483 2363
rect 1869 2261 1903 2295
rect 7113 2261 7147 2295
rect 8677 2261 8711 2295
rect 10977 2261 11011 2295
rect 12909 2261 12943 2295
rect 1501 2057 1535 2091
rect 3801 2057 3835 2091
rect 4077 2057 4111 2091
rect 10425 2057 10459 2091
rect 11069 2057 11103 2091
rect 13277 2057 13311 2091
rect 5549 1989 5583 2023
rect 6745 1989 6779 2023
rect 1685 1921 1719 1955
rect 1869 1921 1903 1955
rect 2053 1921 2087 1955
rect 5825 1921 5859 1955
rect 6193 1921 6227 1955
rect 8677 1921 8711 1955
rect 10885 1921 10919 1955
rect 10977 1921 11011 1955
rect 11253 1921 11287 1955
rect 11529 1921 11563 1955
rect 2329 1853 2363 1887
rect 6469 1853 6503 1887
rect 8217 1853 8251 1887
rect 8953 1853 8987 1887
rect 11805 1853 11839 1887
rect 1869 1717 1903 1751
rect 6009 1717 6043 1751
rect 10701 1717 10735 1751
rect 3341 1513 3375 1547
rect 9045 1513 9079 1547
rect 2881 1445 2915 1479
rect 6929 1445 6963 1479
rect 7757 1445 7791 1479
rect 4445 1377 4479 1411
rect 6193 1377 6227 1411
rect 7389 1377 7423 1411
rect 9689 1377 9723 1411
rect 12081 1377 12115 1411
rect 1409 1309 1443 1343
rect 3525 1309 3559 1343
rect 3875 1309 3909 1343
rect 4721 1309 4755 1343
rect 4813 1309 4847 1343
rect 4997 1309 5031 1343
rect 5549 1309 5583 1343
rect 5825 1309 5859 1343
rect 6745 1309 6779 1343
rect 7481 1309 7515 1343
rect 7757 1309 7791 1343
rect 7941 1309 7975 1343
rect 8585 1309 8619 1343
rect 9229 1309 9263 1343
rect 9413 1309 9447 1343
rect 9505 1309 9539 1343
rect 10057 1309 10091 1343
rect 11529 1309 11563 1343
rect 11713 1309 11747 1343
rect 11897 1309 11931 1343
rect 12633 1309 12667 1343
rect 12725 1309 12759 1343
rect 4169 1241 4203 1275
rect 4353 1241 4387 1275
rect 7389 1241 7423 1275
rect 6561 1173 6595 1207
rect 8401 1173 8435 1207
rect 9873 1173 9907 1207
rect 11253 1173 11287 1207
<< metal1 >>
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 14366 13920 14372 13932
rect 9364 13892 14372 13920
rect 9364 13880 9370 13892
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 11514 13852 11520 13864
rect 8812 13824 11520 13852
rect 8812 13812 8818 13824
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 7006 13744 7012 13796
rect 7064 13784 7070 13796
rect 13354 13784 13360 13796
rect 7064 13756 13360 13784
rect 7064 13744 7070 13756
rect 13354 13744 13360 13756
rect 13412 13744 13418 13796
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 11606 13716 11612 13728
rect 9088 13688 11612 13716
rect 9088 13676 9094 13688
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 1104 13626 13892 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 13892 13626
rect 1104 13552 13892 13574
rect 3510 13512 3516 13524
rect 3471 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 10778 13512 10784 13524
rect 7239 13484 10784 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 2866 13404 2872 13456
rect 2924 13444 2930 13456
rect 6089 13447 6147 13453
rect 6089 13444 6101 13447
rect 2924 13416 6101 13444
rect 2924 13404 2930 13416
rect 6089 13413 6101 13416
rect 6135 13444 6147 13447
rect 7558 13444 7564 13456
rect 6135 13416 7564 13444
rect 6135 13413 6147 13416
rect 6089 13407 6147 13413
rect 7558 13404 7564 13416
rect 7616 13404 7622 13456
rect 7650 13404 7656 13456
rect 7708 13444 7714 13456
rect 8665 13447 8723 13453
rect 7708 13416 7753 13444
rect 7708 13404 7714 13416
rect 8665 13413 8677 13447
rect 8711 13444 8723 13447
rect 9030 13444 9036 13456
rect 8711 13416 9036 13444
rect 8711 13413 8723 13416
rect 8665 13407 8723 13413
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 9125 13447 9183 13453
rect 9125 13413 9137 13447
rect 9171 13444 9183 13447
rect 9171 13416 11560 13444
rect 9171 13413 9183 13416
rect 9125 13407 9183 13413
rect 6917 13379 6975 13385
rect 3160 13348 6592 13376
rect 1854 13308 1860 13320
rect 1815 13280 1860 13308
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 3160 13317 3188 13348
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13277 3203 13311
rect 3145 13271 3203 13277
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 3510 13308 3516 13320
rect 3467 13280 3516 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 1581 13243 1639 13249
rect 1581 13209 1593 13243
rect 1627 13209 1639 13243
rect 2038 13240 2044 13252
rect 1999 13212 2044 13240
rect 1581 13203 1639 13209
rect 1394 13172 1400 13184
rect 1355 13144 1400 13172
rect 1394 13132 1400 13144
rect 1452 13172 1458 13184
rect 1596 13172 1624 13203
rect 2038 13200 2044 13212
rect 2096 13240 2102 13252
rect 2240 13240 2268 13271
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 4212 13280 4353 13308
rect 4212 13268 4218 13280
rect 4341 13277 4353 13280
rect 4387 13277 4399 13311
rect 4890 13308 4896 13320
rect 4851 13280 4896 13308
rect 4341 13271 4399 13277
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 5074 13308 5080 13320
rect 5035 13280 5080 13308
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13308 5595 13311
rect 6178 13308 6184 13320
rect 5583 13280 6184 13308
rect 5583 13277 5595 13280
rect 5537 13271 5595 13277
rect 6178 13268 6184 13280
rect 6236 13308 6242 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6236 13280 6469 13308
rect 6236 13268 6242 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 2682 13240 2688 13252
rect 2096 13212 2268 13240
rect 2643 13212 2688 13240
rect 2096 13200 2102 13212
rect 2682 13200 2688 13212
rect 2740 13200 2746 13252
rect 2774 13200 2780 13252
rect 2832 13240 2838 13252
rect 2961 13243 3019 13249
rect 2832 13212 2877 13240
rect 2832 13200 2838 13212
rect 2961 13209 2973 13243
rect 3007 13240 3019 13243
rect 3050 13240 3056 13252
rect 3007 13212 3056 13240
rect 3007 13209 3019 13212
rect 2961 13203 3019 13209
rect 3050 13200 3056 13212
rect 3108 13200 3114 13252
rect 3878 13200 3884 13252
rect 3936 13240 3942 13252
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 3936 13212 4077 13240
rect 3936 13200 3942 13212
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 4433 13243 4491 13249
rect 4433 13209 4445 13243
rect 4479 13240 4491 13243
rect 4798 13240 4804 13252
rect 4479 13212 4804 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 4798 13200 4804 13212
rect 4856 13200 4862 13252
rect 5626 13200 5632 13252
rect 5684 13240 5690 13252
rect 5684 13212 5729 13240
rect 5684 13200 5690 13212
rect 1452 13144 1624 13172
rect 1673 13175 1731 13181
rect 1452 13132 1458 13144
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 3142 13172 3148 13184
rect 1719 13144 3148 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 3142 13132 3148 13144
rect 3200 13172 3206 13184
rect 3329 13175 3387 13181
rect 3329 13172 3341 13175
rect 3200 13144 3341 13172
rect 3200 13132 3206 13144
rect 3329 13141 3341 13144
rect 3375 13141 3387 13175
rect 3329 13135 3387 13141
rect 4157 13175 4215 13181
rect 4157 13141 4169 13175
rect 4203 13172 4215 13175
rect 4982 13172 4988 13184
rect 4203 13144 4988 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 4982 13132 4988 13144
rect 5040 13172 5046 13184
rect 5442 13172 5448 13184
rect 5040 13144 5448 13172
rect 5040 13132 5046 13144
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 6564 13172 6592 13348
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 9306 13376 9312 13388
rect 6963 13348 9312 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 11146 13376 11152 13388
rect 9539 13348 11152 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 11532 13385 11560 13416
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13345 11575 13379
rect 11517 13339 11575 13345
rect 11606 13336 11612 13388
rect 11664 13376 11670 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 11664 13348 12725 13376
rect 11664 13336 11670 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 7006 13308 7012 13320
rect 6967 13280 7012 13308
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 7432 13280 7481 13308
rect 7432 13268 7438 13280
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 7785 13311 7843 13317
rect 7785 13308 7797 13311
rect 7616 13280 7797 13308
rect 7616 13268 7622 13280
rect 7785 13277 7797 13280
rect 7831 13277 7843 13311
rect 7785 13271 7843 13277
rect 8110 13268 8116 13320
rect 8168 13308 8174 13320
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 8168 13280 8217 13308
rect 8168 13268 8174 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13277 8355 13311
rect 8754 13308 8760 13320
rect 8715 13280 8760 13308
rect 8297 13271 8355 13277
rect 6641 13243 6699 13249
rect 6641 13209 6653 13243
rect 6687 13240 6699 13243
rect 7282 13240 7288 13252
rect 6687 13212 7144 13240
rect 7243 13212 7288 13240
rect 6687 13209 6699 13212
rect 6641 13203 6699 13209
rect 7006 13172 7012 13184
rect 6564 13144 7012 13172
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 7116 13172 7144 13212
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 7926 13240 7932 13252
rect 7887 13212 7932 13240
rect 7926 13200 7932 13212
rect 7984 13200 7990 13252
rect 8018 13200 8024 13252
rect 8076 13240 8082 13252
rect 8076 13212 8121 13240
rect 8076 13200 8082 13212
rect 7558 13172 7564 13184
rect 7116 13144 7564 13172
rect 7558 13132 7564 13144
rect 7616 13172 7622 13184
rect 8312 13172 8340 13271
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13308 9459 13311
rect 9582 13308 9588 13320
rect 9447 13280 9588 13308
rect 9447 13277 9459 13280
rect 9401 13271 9459 13277
rect 8956 13240 8984 13271
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13308 10103 13311
rect 10226 13308 10232 13320
rect 10091 13280 10232 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 10468 13280 10609 13308
rect 10468 13268 10474 13280
rect 10597 13277 10609 13280
rect 10643 13277 10655 13311
rect 10778 13308 10784 13320
rect 10739 13280 10784 13308
rect 10597 13271 10655 13277
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11112 13280 11345 13308
rect 11112 13268 11118 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 12069 13311 12127 13317
rect 12069 13308 12081 13311
rect 11333 13271 11391 13277
rect 11440 13280 12081 13308
rect 10318 13240 10324 13252
rect 8956 13212 10180 13240
rect 10279 13212 10324 13240
rect 7616 13144 8340 13172
rect 8481 13175 8539 13181
rect 7616 13132 7622 13144
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 8570 13172 8576 13184
rect 8527 13144 8576 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 9306 13172 9312 13184
rect 9267 13144 9312 13172
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 10152 13172 10180 13212
rect 10318 13200 10324 13212
rect 10376 13200 10382 13252
rect 10873 13243 10931 13249
rect 10873 13209 10885 13243
rect 10919 13209 10931 13243
rect 10873 13203 10931 13209
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 10152 13144 10425 13172
rect 10413 13141 10425 13144
rect 10459 13172 10471 13175
rect 10686 13172 10692 13184
rect 10459 13144 10692 13172
rect 10459 13141 10471 13144
rect 10413 13135 10471 13141
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 10888 13172 10916 13203
rect 11238 13200 11244 13252
rect 11296 13240 11302 13252
rect 11440 13240 11468 13280
rect 12069 13277 12081 13280
rect 12115 13277 12127 13311
rect 12069 13271 12127 13277
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12802 13308 12808 13320
rect 12216 13280 12261 13308
rect 12763 13280 12808 13308
rect 12216 13268 12222 13280
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 12952 13280 13369 13308
rect 12952 13268 12958 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 11296 13212 11468 13240
rect 11296 13200 11302 13212
rect 11514 13200 11520 13252
rect 11572 13240 11578 13252
rect 11609 13243 11667 13249
rect 11609 13240 11621 13243
rect 11572 13212 11621 13240
rect 11572 13200 11578 13212
rect 11609 13209 11621 13212
rect 11655 13209 11667 13243
rect 12618 13240 12624 13252
rect 12579 13212 12624 13240
rect 11609 13203 11667 13209
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 13262 13240 13268 13252
rect 13223 13212 13268 13240
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13170 13172 13176 13184
rect 10836 13144 13176 13172
rect 10836 13132 10842 13144
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 13541 13175 13599 13181
rect 13541 13141 13553 13175
rect 13587 13172 13599 13175
rect 13722 13172 13728 13184
rect 13587 13144 13728 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 1104 13082 13892 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 13892 13082
rect 1104 13008 13892 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 2774 12968 2780 12980
rect 1627 12940 2780 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 2774 12928 2780 12940
rect 2832 12928 2838 12980
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 9490 12968 9496 12980
rect 7708 12940 9496 12968
rect 7708 12928 7714 12940
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9640 12940 10456 12968
rect 9640 12928 9646 12940
rect 1946 12860 1952 12912
rect 2004 12900 2010 12912
rect 4433 12903 4491 12909
rect 4433 12900 4445 12903
rect 2004 12872 4445 12900
rect 2004 12860 2010 12872
rect 4433 12869 4445 12872
rect 4479 12900 4491 12903
rect 5258 12900 5264 12912
rect 4479 12872 5264 12900
rect 4479 12869 4491 12872
rect 4433 12863 4491 12869
rect 5258 12860 5264 12872
rect 5316 12860 5322 12912
rect 6178 12900 6184 12912
rect 6139 12872 6184 12900
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 8018 12900 8024 12912
rect 7064 12872 8024 12900
rect 7064 12860 7070 12872
rect 8018 12860 8024 12872
rect 8076 12860 8082 12912
rect 8389 12903 8447 12909
rect 8389 12869 8401 12903
rect 8435 12900 8447 12903
rect 10042 12900 10048 12912
rect 8435 12872 9444 12900
rect 9955 12872 10048 12900
rect 8435 12869 8447 12872
rect 8389 12863 8447 12869
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 2590 12832 2596 12844
rect 2551 12804 2596 12832
rect 1673 12795 1731 12801
rect 1688 12696 1716 12795
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 3050 12832 3056 12844
rect 2823 12804 3056 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3476 12804 3709 12832
rect 3476 12792 3482 12804
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 4614 12832 4620 12844
rect 4527 12804 4620 12832
rect 3697 12795 3755 12801
rect 4614 12792 4620 12804
rect 4672 12832 4678 12844
rect 5074 12832 5080 12844
rect 4672 12804 5080 12832
rect 4672 12792 4678 12804
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5442 12792 5448 12844
rect 5500 12832 5506 12844
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5500 12804 5549 12832
rect 5500 12792 5506 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 6362 12832 6368 12844
rect 6323 12804 6368 12832
rect 5537 12795 5595 12801
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7558 12832 7564 12844
rect 7248 12804 7564 12832
rect 7248 12792 7254 12804
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 9416 12841 9444 12872
rect 10042 12860 10048 12872
rect 10100 12900 10106 12912
rect 10318 12900 10324 12912
rect 10100 12872 10324 12900
rect 10100 12860 10106 12872
rect 10318 12860 10324 12872
rect 10376 12860 10382 12912
rect 10428 12909 10456 12940
rect 10778 12928 10784 12980
rect 10836 12968 10842 12980
rect 10962 12968 10968 12980
rect 10836 12940 10968 12968
rect 10836 12928 10842 12940
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 13354 12968 13360 12980
rect 13315 12940 13360 12968
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 10413 12903 10471 12909
rect 10413 12869 10425 12903
rect 10459 12869 10471 12903
rect 10413 12863 10471 12869
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 11882 12900 11888 12912
rect 10744 12872 11888 12900
rect 10744 12860 10750 12872
rect 11882 12860 11888 12872
rect 11940 12900 11946 12912
rect 11940 12872 12480 12900
rect 11940 12860 11946 12872
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7668 12804 8217 12832
rect 1762 12724 1768 12776
rect 1820 12764 1826 12776
rect 2317 12767 2375 12773
rect 1820 12736 1865 12764
rect 1820 12724 1826 12736
rect 2317 12733 2329 12767
rect 2363 12733 2375 12767
rect 2317 12727 2375 12733
rect 2222 12696 2228 12708
rect 1688 12668 2228 12696
rect 2222 12656 2228 12668
rect 2280 12656 2286 12708
rect 2332 12696 2360 12727
rect 7668 12708 7696 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 10137 12835 10195 12841
rect 10137 12832 10149 12835
rect 9447 12804 10149 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 10137 12801 10149 12804
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 2409 12699 2467 12705
rect 2409 12696 2421 12699
rect 2332 12668 2421 12696
rect 2409 12665 2421 12668
rect 2455 12665 2467 12699
rect 2409 12659 2467 12665
rect 3510 12656 3516 12708
rect 3568 12696 3574 12708
rect 3878 12696 3884 12708
rect 3568 12668 3884 12696
rect 3568 12656 3574 12668
rect 3878 12656 3884 12668
rect 3936 12696 3942 12708
rect 4249 12699 4307 12705
rect 4249 12696 4261 12699
rect 3936 12668 4261 12696
rect 3936 12656 3942 12668
rect 4249 12665 4261 12668
rect 4295 12665 4307 12699
rect 7650 12696 7656 12708
rect 7611 12668 7656 12696
rect 4249 12659 4307 12665
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 8496 12628 8524 12795
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 10152 12764 10180 12795
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10778 12832 10784 12844
rect 10284 12804 10784 12832
rect 10284 12792 10290 12804
rect 10778 12792 10784 12804
rect 10836 12832 10842 12844
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 10836 12804 11069 12832
rect 10836 12792 10842 12804
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 12158 12832 12164 12844
rect 11563 12804 12164 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 11348 12764 11376 12795
rect 9548 12736 10088 12764
rect 10152 12736 11376 12764
rect 9548 12724 9554 12736
rect 9306 12656 9312 12708
rect 9364 12696 9370 12708
rect 10060 12696 10088 12736
rect 11532 12696 11560 12795
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 12452 12841 12480 12872
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12676 12872 13093 12900
rect 12676 12860 12682 12872
rect 13081 12869 13093 12872
rect 13127 12900 13139 12903
rect 13265 12903 13323 12909
rect 13265 12900 13277 12903
rect 13127 12872 13277 12900
rect 13127 12869 13139 12872
rect 13081 12863 13139 12869
rect 13265 12869 13277 12872
rect 13311 12869 13323 12903
rect 13265 12863 13323 12869
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 9364 12668 9812 12696
rect 10060 12668 11560 12696
rect 9364 12656 9370 12668
rect 9674 12628 9680 12640
rect 5408 12600 9680 12628
rect 5408 12588 5414 12600
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 9784 12628 9812 12668
rect 9950 12628 9956 12640
rect 9784 12600 9956 12628
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10134 12588 10140 12640
rect 10192 12628 10198 12640
rect 12894 12628 12900 12640
rect 10192 12600 12900 12628
rect 10192 12588 10198 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 1104 12538 13892 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 13892 12538
rect 1104 12464 13892 12486
rect 4062 12424 4068 12436
rect 4023 12396 4068 12424
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4982 12424 4988 12436
rect 4212 12396 4988 12424
rect 4212 12384 4218 12396
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 5261 12427 5319 12433
rect 5261 12393 5273 12427
rect 5307 12424 5319 12427
rect 5626 12424 5632 12436
rect 5307 12396 5632 12424
rect 5307 12393 5319 12396
rect 5261 12387 5319 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 8757 12427 8815 12433
rect 5736 12396 7788 12424
rect 2682 12316 2688 12368
rect 2740 12356 2746 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2740 12328 2789 12356
rect 2740 12316 2746 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 3418 12356 3424 12368
rect 3379 12328 3424 12356
rect 2777 12319 2835 12325
rect 1489 12223 1547 12229
rect 1489 12189 1501 12223
rect 1535 12220 1547 12223
rect 2038 12220 2044 12232
rect 1535 12192 2044 12220
rect 1535 12189 1547 12192
rect 1489 12183 1547 12189
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 2792 12220 2820 12319
rect 3418 12316 3424 12328
rect 3476 12316 3482 12368
rect 4890 12316 4896 12368
rect 4948 12356 4954 12368
rect 5736 12356 5764 12396
rect 4948 12328 5764 12356
rect 6825 12359 6883 12365
rect 4948 12316 4954 12328
rect 6825 12325 6837 12359
rect 6871 12356 6883 12359
rect 7650 12356 7656 12368
rect 6871 12328 7656 12356
rect 6871 12325 6883 12328
rect 6825 12319 6883 12325
rect 7650 12316 7656 12328
rect 7708 12316 7714 12368
rect 7760 12356 7788 12396
rect 8757 12393 8769 12427
rect 8803 12424 8815 12427
rect 8846 12424 8852 12436
rect 8803 12396 8852 12424
rect 8803 12393 8815 12396
rect 8757 12387 8815 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 10505 12427 10563 12433
rect 10505 12393 10517 12427
rect 10551 12424 10563 12427
rect 10686 12424 10692 12436
rect 10551 12396 10692 12424
rect 10551 12393 10563 12396
rect 10505 12387 10563 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 9033 12359 9091 12365
rect 9033 12356 9045 12359
rect 7760 12328 9045 12356
rect 9033 12325 9045 12328
rect 9079 12325 9091 12359
rect 9766 12356 9772 12368
rect 9033 12319 9091 12325
rect 9692 12328 9772 12356
rect 4908 12288 4936 12316
rect 4172 12260 4936 12288
rect 4172 12229 4200 12260
rect 4982 12248 4988 12300
rect 5040 12288 5046 12300
rect 6546 12288 6552 12300
rect 5040 12260 6552 12288
rect 5040 12248 5046 12260
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 7282 12288 7288 12300
rect 6963 12260 7288 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 7834 12248 7840 12300
rect 7892 12288 7898 12300
rect 8570 12288 8576 12300
rect 7892 12260 8156 12288
rect 8531 12260 8576 12288
rect 7892 12248 7898 12260
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 2792 12192 3249 12220
rect 3237 12189 3249 12192
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4798 12220 4804 12232
rect 4759 12192 4804 12220
rect 4157 12183 4215 12189
rect 3896 12152 3924 12183
rect 4798 12180 4804 12192
rect 4856 12220 4862 12232
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 4856 12192 5181 12220
rect 4856 12180 4862 12192
rect 5169 12189 5181 12192
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 6362 12220 6368 12232
rect 5592 12192 6368 12220
rect 5592 12180 5598 12192
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12220 7067 12223
rect 7190 12220 7196 12232
rect 7055 12192 7196 12220
rect 7055 12189 7067 12192
rect 7009 12183 7067 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7616 12192 7941 12220
rect 7616 12180 7622 12192
rect 7929 12189 7941 12192
rect 7975 12220 7987 12223
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7975 12192 8033 12220
rect 7975 12189 7987 12192
rect 7929 12183 7987 12189
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8128 12220 8156 12260
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 8938 12248 8944 12300
rect 8996 12288 9002 12300
rect 9692 12297 9720 12328
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 10042 12316 10048 12368
rect 10100 12356 10106 12368
rect 10137 12359 10195 12365
rect 10137 12356 10149 12359
rect 10100 12328 10149 12356
rect 10100 12316 10106 12328
rect 10137 12325 10149 12328
rect 10183 12325 10195 12359
rect 10137 12319 10195 12325
rect 10318 12316 10324 12368
rect 10376 12316 10382 12368
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 11388 12328 11928 12356
rect 11388 12316 11394 12328
rect 9677 12291 9735 12297
rect 8996 12260 9347 12288
rect 8996 12248 9002 12260
rect 9214 12229 9220 12232
rect 9212 12220 9220 12229
rect 8128 12192 9076 12220
rect 9175 12192 9220 12220
rect 8021 12183 8079 12189
rect 5074 12152 5080 12164
rect 3896 12124 5080 12152
rect 5074 12112 5080 12124
rect 5132 12112 5138 12164
rect 5445 12155 5503 12161
rect 5445 12121 5457 12155
rect 5491 12121 5503 12155
rect 5445 12115 5503 12121
rect 5629 12155 5687 12161
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 5718 12152 5724 12164
rect 5675 12124 5724 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 3602 12084 3608 12096
rect 3384 12056 3608 12084
rect 3384 12044 3390 12056
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 4982 12044 4988 12096
rect 5040 12084 5046 12096
rect 5460 12084 5488 12115
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 5813 12155 5871 12161
rect 5813 12121 5825 12155
rect 5859 12152 5871 12155
rect 5902 12152 5908 12164
rect 5859 12124 5908 12152
rect 5859 12121 5871 12124
rect 5813 12115 5871 12121
rect 5902 12112 5908 12124
rect 5960 12112 5966 12164
rect 6086 12152 6092 12164
rect 6047 12124 6092 12152
rect 6086 12112 6092 12124
rect 6144 12112 6150 12164
rect 6273 12155 6331 12161
rect 6273 12121 6285 12155
rect 6319 12152 6331 12155
rect 6638 12152 6644 12164
rect 6319 12124 6644 12152
rect 6319 12121 6331 12124
rect 6273 12115 6331 12121
rect 6638 12112 6644 12124
rect 6696 12112 6702 12164
rect 7285 12155 7343 12161
rect 7285 12121 7297 12155
rect 7331 12152 7343 12155
rect 7374 12152 7380 12164
rect 7331 12124 7380 12152
rect 7331 12121 7343 12124
rect 7285 12115 7343 12121
rect 7374 12112 7380 12124
rect 7432 12152 7438 12164
rect 8481 12155 8539 12161
rect 8481 12152 8493 12155
rect 7432 12124 8493 12152
rect 7432 12112 7438 12124
rect 8481 12121 8493 12124
rect 8527 12121 8539 12155
rect 9048 12152 9076 12192
rect 9212 12183 9220 12192
rect 9214 12180 9220 12183
rect 9272 12180 9278 12232
rect 9319 12220 9347 12260
rect 9677 12257 9689 12291
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10229 12291 10287 12297
rect 10229 12288 10241 12291
rect 10008 12260 10241 12288
rect 10008 12248 10014 12260
rect 10229 12257 10241 12260
rect 10275 12257 10287 12291
rect 10336 12288 10364 12316
rect 11698 12288 11704 12300
rect 10336 12260 11704 12288
rect 10229 12251 10287 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11900 12288 11928 12328
rect 11900 12260 12020 12288
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 9319 12192 9413 12220
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 9585 12223 9643 12229
rect 9585 12220 9597 12223
rect 9548 12192 9597 12220
rect 9548 12180 9554 12192
rect 9585 12189 9597 12192
rect 9631 12189 9643 12223
rect 9585 12183 9643 12189
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 9824 12192 10333 12220
rect 9824 12180 9830 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 10686 12220 10692 12232
rect 10551 12192 10692 12220
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10962 12220 10968 12232
rect 10875 12192 10968 12220
rect 10962 12180 10968 12192
rect 11020 12220 11026 12232
rect 11238 12220 11244 12232
rect 11020 12192 11244 12220
rect 11020 12180 11026 12192
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11572 12192 11621 12220
rect 11572 12180 11578 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 11609 12183 11667 12189
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 11992 12229 12020 12260
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 11977 12183 12035 12189
rect 12084 12192 12541 12220
rect 9309 12155 9367 12161
rect 9309 12152 9321 12155
rect 9048 12124 9321 12152
rect 8481 12115 8539 12121
rect 9309 12121 9321 12124
rect 9355 12152 9367 12155
rect 9355 12124 11008 12152
rect 9355 12121 9367 12124
rect 9309 12115 9367 12121
rect 5040 12056 5488 12084
rect 5040 12044 5046 12056
rect 6178 12044 6184 12096
rect 6236 12084 6242 12096
rect 7650 12084 7656 12096
rect 6236 12056 7656 12084
rect 6236 12044 6242 12056
rect 7650 12044 7656 12056
rect 7708 12084 7714 12096
rect 8018 12084 8024 12096
rect 7708 12056 8024 12084
rect 7708 12044 7714 12056
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 10980 12084 11008 12124
rect 11054 12112 11060 12164
rect 11112 12152 11118 12164
rect 12084 12152 12112 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 13170 12220 13176 12232
rect 13131 12192 13176 12220
rect 12529 12183 12587 12189
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 12342 12152 12348 12164
rect 11112 12124 12112 12152
rect 12303 12124 12348 12152
rect 11112 12112 11118 12124
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 13446 12152 13452 12164
rect 13407 12124 13452 12152
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 12066 12084 12072 12096
rect 10980 12056 12072 12084
rect 12066 12044 12072 12056
rect 12124 12084 12130 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 12124 12056 12173 12084
rect 12124 12044 12130 12056
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 12161 12047 12219 12053
rect 1104 11994 13892 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 13892 11994
rect 1104 11920 13892 11942
rect 6178 11880 6184 11892
rect 4908 11852 6184 11880
rect 2222 11812 2228 11824
rect 2183 11784 2228 11812
rect 2222 11772 2228 11784
rect 2280 11772 2286 11824
rect 2501 11815 2559 11821
rect 2501 11781 2513 11815
rect 2547 11812 2559 11815
rect 2590 11812 2596 11824
rect 2547 11784 2596 11812
rect 2547 11781 2559 11784
rect 2501 11775 2559 11781
rect 2590 11772 2596 11784
rect 2648 11772 2654 11824
rect 3602 11772 3608 11824
rect 3660 11812 3666 11824
rect 4617 11815 4675 11821
rect 3660 11784 4200 11812
rect 3660 11772 3666 11784
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 1762 11744 1768 11756
rect 1627 11716 1768 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 1762 11704 1768 11716
rect 1820 11704 1826 11756
rect 2682 11704 2688 11756
rect 2740 11744 2746 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2740 11716 2789 11744
rect 2740 11704 2746 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 3050 11744 3056 11756
rect 3011 11716 3056 11744
rect 2777 11707 2835 11713
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 3786 11744 3792 11756
rect 3476 11716 3792 11744
rect 3476 11704 3482 11716
rect 3786 11704 3792 11716
rect 3844 11744 3850 11756
rect 3881 11747 3939 11753
rect 3881 11744 3893 11747
rect 3844 11716 3893 11744
rect 3844 11704 3850 11716
rect 3881 11713 3893 11716
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 3970 11704 3976 11756
rect 4028 11744 4034 11756
rect 4172 11744 4200 11784
rect 4617 11781 4629 11815
rect 4663 11812 4675 11815
rect 4798 11812 4804 11824
rect 4663 11784 4804 11812
rect 4663 11781 4675 11784
rect 4617 11775 4675 11781
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 4473 11747 4531 11753
rect 4473 11744 4485 11747
rect 4028 11716 4073 11744
rect 4172 11716 4485 11744
rect 4028 11704 4034 11716
rect 4473 11713 4485 11716
rect 4519 11713 4531 11747
rect 4706 11744 4712 11756
rect 4667 11716 4712 11744
rect 4473 11707 4531 11713
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 4908 11753 4936 11852
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 6328 11852 6469 11880
rect 6328 11840 6334 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 7377 11883 7435 11889
rect 7377 11880 7389 11883
rect 6604 11852 7389 11880
rect 6604 11840 6610 11852
rect 7377 11849 7389 11852
rect 7423 11880 7435 11883
rect 7834 11880 7840 11892
rect 7423 11852 7840 11880
rect 7423 11849 7435 11852
rect 7377 11843 7435 11849
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 7926 11840 7932 11892
rect 7984 11840 7990 11892
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 8113 11883 8171 11889
rect 8113 11880 8125 11883
rect 8076 11852 8125 11880
rect 8076 11840 8082 11852
rect 8113 11849 8125 11852
rect 8159 11849 8171 11883
rect 8113 11843 8171 11849
rect 8404 11852 8616 11880
rect 5997 11815 6055 11821
rect 5997 11781 6009 11815
rect 6043 11812 6055 11815
rect 6086 11812 6092 11824
rect 6043 11784 6092 11812
rect 6043 11781 6055 11784
rect 5997 11775 6055 11781
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 7944 11812 7972 11840
rect 8202 11812 8208 11824
rect 6420 11784 6868 11812
rect 6420 11772 6426 11784
rect 5258 11753 5264 11756
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11713 4951 11747
rect 5256 11744 5264 11753
rect 5219 11716 5264 11744
rect 4893 11707 4951 11713
rect 5256 11707 5264 11716
rect 5258 11704 5264 11707
rect 5316 11704 5322 11756
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11713 5411 11747
rect 5353 11707 5411 11713
rect 1394 11608 1400 11620
rect 1355 11580 1400 11608
rect 1394 11568 1400 11580
rect 1452 11568 1458 11620
rect 1780 11608 1808 11704
rect 2866 11636 2872 11688
rect 2924 11676 2930 11688
rect 3510 11676 3516 11688
rect 2924 11648 3516 11676
rect 2924 11636 2930 11648
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 4065 11679 4123 11685
rect 4065 11676 4077 11679
rect 3651 11648 4077 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 4065 11645 4077 11648
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 4264 11648 4752 11676
rect 4264 11608 4292 11648
rect 1780 11580 4292 11608
rect 4341 11611 4399 11617
rect 4341 11577 4353 11611
rect 4387 11608 4399 11611
rect 4614 11608 4620 11620
rect 4387 11580 4620 11608
rect 4387 11577 4399 11580
rect 4341 11571 4399 11577
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 4724 11608 4752 11648
rect 4798 11636 4804 11688
rect 4856 11676 4862 11688
rect 5373 11676 5401 11707
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 5629 11747 5687 11753
rect 5500 11716 5545 11744
rect 5500 11704 5506 11716
rect 5629 11713 5641 11747
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6454 11744 6460 11756
rect 6227 11716 6460 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 5644 11676 5672 11707
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 6840 11753 6868 11784
rect 6932 11784 8208 11812
rect 6932 11753 6960 11784
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 6825 11747 6883 11753
rect 6696 11716 6741 11744
rect 6696 11704 6702 11716
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 7061 11747 7119 11753
rect 7061 11713 7073 11747
rect 7107 11744 7119 11747
rect 7466 11744 7472 11756
rect 7107 11716 7472 11744
rect 7107 11713 7119 11716
rect 7061 11707 7119 11713
rect 5718 11676 5724 11688
rect 4856 11648 5401 11676
rect 5631 11648 5724 11676
rect 4856 11636 4862 11648
rect 5718 11636 5724 11648
rect 5776 11676 5782 11688
rect 6546 11676 6552 11688
rect 5776 11648 6552 11676
rect 5776 11636 5782 11648
rect 6546 11636 6552 11648
rect 6604 11636 6610 11688
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 6932 11676 6960 11707
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 7742 11744 7748 11756
rect 7703 11716 7748 11744
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 8001 11747 8059 11753
rect 8001 11713 8013 11747
rect 8047 11744 8059 11747
rect 8404 11744 8432 11852
rect 8588 11812 8616 11852
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 10502 11880 10508 11892
rect 8812 11852 10508 11880
rect 8812 11840 8818 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10873 11883 10931 11889
rect 10873 11849 10885 11883
rect 10919 11880 10931 11883
rect 11422 11880 11428 11892
rect 10919 11852 11428 11880
rect 10919 11849 10931 11852
rect 10873 11843 10931 11849
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11572 11852 11652 11880
rect 11572 11840 11578 11852
rect 8846 11812 8852 11824
rect 8588 11784 8852 11812
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 9122 11772 9128 11824
rect 9180 11812 9186 11824
rect 9180 11784 10180 11812
rect 9180 11772 9186 11784
rect 8047 11716 8432 11744
rect 8047 11713 8059 11716
rect 8001 11707 8059 11713
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 9217 11747 9275 11753
rect 8536 11716 8581 11744
rect 8536 11704 8542 11716
rect 9217 11713 9229 11747
rect 9263 11713 9275 11747
rect 9398 11744 9404 11756
rect 9359 11716 9404 11744
rect 9217 11707 9275 11713
rect 6788 11648 6960 11676
rect 6788 11636 6794 11648
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 7892 11648 8217 11676
rect 7892 11636 7898 11648
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8846 11676 8852 11688
rect 8343 11648 8852 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 8941 11679 8999 11685
rect 8941 11645 8953 11679
rect 8987 11676 8999 11679
rect 9232 11676 9260 11707
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 9508 11753 9536 11784
rect 10152 11756 10180 11784
rect 10226 11772 10232 11824
rect 10284 11812 10290 11824
rect 10284 11784 10329 11812
rect 10284 11772 10290 11784
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11713 9551 11747
rect 9766 11744 9772 11756
rect 9727 11716 9772 11744
rect 9493 11707 9551 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 8987 11648 9260 11676
rect 8987 11645 8999 11648
rect 8941 11639 8999 11645
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 10060 11676 10088 11707
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10192 11716 10517 11744
rect 10192 11704 10198 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 10761 11747 10819 11753
rect 10761 11713 10773 11747
rect 10807 11744 10819 11747
rect 11238 11744 11244 11756
rect 10807 11716 11244 11744
rect 10807 11713 10819 11716
rect 10761 11707 10819 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 11514 11744 11520 11756
rect 11379 11716 11520 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 11624 11744 11652 11852
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11624 11716 11713 11744
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11848 11716 11897 11744
rect 11848 11704 11854 11716
rect 11885 11713 11897 11716
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12802 11744 12808 11756
rect 12032 11716 12808 11744
rect 12032 11704 12038 11716
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13446 11744 13452 11756
rect 13407 11716 13452 11744
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 9364 11648 10456 11676
rect 9364 11636 9370 11648
rect 10321 11611 10379 11617
rect 10321 11608 10333 11611
rect 4724 11580 10333 11608
rect 10321 11577 10333 11580
rect 10367 11577 10379 11611
rect 10321 11571 10379 11577
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 3697 11543 3755 11549
rect 3697 11540 3709 11543
rect 3660 11512 3709 11540
rect 3660 11500 3666 11512
rect 3697 11509 3709 11512
rect 3743 11509 3755 11543
rect 3697 11503 3755 11509
rect 5077 11543 5135 11549
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 5350 11540 5356 11552
rect 5123 11512 5356 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 5994 11500 6000 11552
rect 6052 11540 6058 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 6052 11512 7205 11540
rect 6052 11500 6058 11512
rect 7193 11509 7205 11512
rect 7239 11509 7251 11543
rect 7558 11540 7564 11552
rect 7519 11512 7564 11540
rect 7193 11503 7251 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 7926 11500 7932 11552
rect 7984 11540 7990 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 7984 11512 8585 11540
rect 7984 11500 7990 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 8573 11503 8631 11509
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9490 11540 9496 11552
rect 9088 11512 9496 11540
rect 9088 11500 9094 11512
rect 9490 11500 9496 11512
rect 9548 11540 9554 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9548 11512 9965 11540
rect 9548 11500 9554 11512
rect 9953 11509 9965 11512
rect 9999 11509 10011 11543
rect 10428 11540 10456 11648
rect 10594 11636 10600 11688
rect 10652 11676 10658 11688
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10652 11648 10977 11676
rect 10652 11636 10658 11648
rect 10965 11645 10977 11648
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11146 11676 11152 11688
rect 11103 11648 11152 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11256 11676 11284 11704
rect 12158 11676 12164 11688
rect 11256 11648 12164 11676
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 10502 11568 10508 11620
rect 10560 11608 10566 11620
rect 12342 11608 12348 11620
rect 10560 11580 12348 11608
rect 10560 11568 10566 11580
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 13262 11608 13268 11620
rect 13223 11580 13268 11608
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 10870 11540 10876 11552
rect 10428 11512 10876 11540
rect 9953 11503 10011 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 11238 11540 11244 11552
rect 11199 11512 11244 11540
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11609 11543 11667 11549
rect 11609 11509 11621 11543
rect 11655 11540 11667 11543
rect 11974 11540 11980 11552
rect 11655 11512 11980 11540
rect 11655 11509 11667 11512
rect 11609 11503 11667 11509
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 1104 11450 13892 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 13892 11450
rect 1104 11376 13892 11398
rect 4893 11339 4951 11345
rect 4893 11305 4905 11339
rect 4939 11336 4951 11339
rect 5258 11336 5264 11348
rect 4939 11308 5264 11336
rect 4939 11305 4951 11308
rect 4893 11299 4951 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 5534 11336 5540 11348
rect 5495 11308 5540 11336
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6914 11336 6920 11348
rect 6503 11308 6920 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7469 11339 7527 11345
rect 7469 11305 7481 11339
rect 7515 11336 7527 11339
rect 7558 11336 7564 11348
rect 7515 11308 7564 11336
rect 7515 11305 7527 11308
rect 7469 11299 7527 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 7926 11336 7932 11348
rect 7699 11308 7932 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 7926 11296 7932 11308
rect 7984 11336 7990 11348
rect 8662 11336 8668 11348
rect 7984 11308 8668 11336
rect 7984 11296 7990 11308
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 9088 11308 9137 11336
rect 9088 11296 9094 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9125 11299 9183 11305
rect 10781 11339 10839 11345
rect 10781 11305 10793 11339
rect 10827 11336 10839 11339
rect 10962 11336 10968 11348
rect 10827 11308 10968 11336
rect 10827 11305 10839 11308
rect 10781 11299 10839 11305
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 11514 11296 11520 11348
rect 11572 11336 11578 11348
rect 11572 11308 11617 11336
rect 11572 11296 11578 11308
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 11940 11308 12480 11336
rect 11940 11296 11946 11308
rect 1857 11271 1915 11277
rect 1857 11237 1869 11271
rect 1903 11268 1915 11271
rect 2682 11268 2688 11280
rect 1903 11240 2688 11268
rect 1903 11237 1915 11240
rect 1857 11231 1915 11237
rect 2682 11228 2688 11240
rect 2740 11228 2746 11280
rect 3068 11240 4752 11268
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 3068 11209 3096 11240
rect 3053 11203 3111 11209
rect 1452 11172 2452 11200
rect 1452 11160 1458 11172
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2424 11141 2452 11172
rect 3053 11169 3065 11203
rect 3099 11169 3111 11203
rect 3602 11200 3608 11212
rect 3563 11172 3608 11200
rect 3053 11163 3111 11169
rect 3602 11160 3608 11172
rect 3660 11160 3666 11212
rect 4724 11200 4752 11240
rect 5166 11228 5172 11280
rect 5224 11268 5230 11280
rect 5721 11271 5779 11277
rect 5721 11268 5733 11271
rect 5224 11240 5733 11268
rect 5224 11228 5230 11240
rect 5721 11237 5733 11240
rect 5767 11268 5779 11271
rect 6178 11268 6184 11280
rect 5767 11240 6184 11268
rect 5767 11237 5779 11240
rect 5721 11231 5779 11237
rect 6178 11228 6184 11240
rect 6236 11228 6242 11280
rect 6270 11228 6276 11280
rect 6328 11228 6334 11280
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 7282 11268 7288 11280
rect 7064 11240 7288 11268
rect 7064 11228 7070 11240
rect 7282 11228 7288 11240
rect 7340 11228 7346 11280
rect 9674 11268 9680 11280
rect 7835 11240 9680 11268
rect 4890 11200 4896 11212
rect 4724 11172 4896 11200
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 3513 11135 3571 11141
rect 2731 11104 3464 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 1765 11067 1823 11073
rect 1765 11064 1777 11067
rect 1627 11036 1777 11064
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 1765 11033 1777 11036
rect 1811 11033 1823 11067
rect 2332 11064 2360 11092
rect 2869 11067 2927 11073
rect 2869 11064 2881 11067
rect 2332 11036 2881 11064
rect 1765 11027 1823 11033
rect 2869 11033 2881 11036
rect 2915 11033 2927 11067
rect 3436 11064 3464 11104
rect 3513 11101 3525 11135
rect 3559 11132 3571 11135
rect 3970 11132 3976 11144
rect 3559 11104 3976 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 4724 11141 4752 11172
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4982 11132 4988 11144
rect 4943 11104 4988 11132
rect 4709 11095 4767 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5350 11092 5356 11144
rect 5408 11141 5414 11144
rect 5408 11132 5416 11141
rect 5902 11132 5908 11144
rect 5408 11104 5453 11132
rect 5863 11104 5908 11132
rect 5408 11095 5416 11104
rect 5408 11092 5414 11095
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6293 11141 6321 11228
rect 6454 11160 6460 11212
rect 6512 11200 6518 11212
rect 6512 11172 6994 11200
rect 6512 11160 6518 11172
rect 6278 11135 6336 11141
rect 6278 11101 6290 11135
rect 6324 11101 6336 11135
rect 6278 11095 6336 11101
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 6822 11132 6828 11144
rect 6696 11104 6741 11132
rect 6783 11104 6828 11132
rect 6696 11092 6702 11104
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 6966 11119 6994 11172
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 7835 11200 7863 11240
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 10134 11228 10140 11280
rect 10192 11228 10198 11280
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 11974 11268 11980 11280
rect 10928 11240 11192 11268
rect 10928 11228 10934 11240
rect 7616 11172 7863 11200
rect 7616 11160 7622 11172
rect 8202 11160 8208 11212
rect 8260 11160 8266 11212
rect 8665 11203 8723 11209
rect 8665 11169 8677 11203
rect 8711 11200 8723 11203
rect 9950 11200 9956 11212
rect 8711 11172 9956 11200
rect 8711 11169 8723 11172
rect 8665 11163 8723 11169
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 10152 11200 10180 11228
rect 10152 11172 10640 11200
rect 6942 11113 7000 11119
rect 6942 11079 6954 11113
rect 6988 11079 7000 11113
rect 3602 11064 3608 11076
rect 3436 11036 3608 11064
rect 2869 11027 2927 11033
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 3786 11064 3792 11076
rect 3747 11036 3792 11064
rect 3786 11024 3792 11036
rect 3844 11024 3850 11076
rect 5166 11064 5172 11076
rect 5127 11036 5172 11064
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 6089 11067 6147 11073
rect 6089 11064 6101 11067
rect 5316 11036 5361 11064
rect 5460 11036 6101 11064
rect 5316 11024 5322 11036
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 1946 10996 1952 11008
rect 1719 10968 1952 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 1946 10956 1952 10968
rect 2004 10956 2010 11008
rect 2501 10999 2559 11005
rect 2501 10965 2513 10999
rect 2547 10996 2559 10999
rect 3142 10996 3148 11008
rect 2547 10968 3148 10996
rect 2547 10965 2559 10968
rect 2501 10959 2559 10965
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 3620 10996 3648 11024
rect 5460 11008 5488 11036
rect 5442 10996 5448 11008
rect 3620 10968 5448 10996
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 6012 10996 6040 11036
rect 6089 11033 6101 11036
rect 6135 11033 6147 11067
rect 6089 11027 6147 11033
rect 6181 11067 6239 11073
rect 6181 11033 6193 11067
rect 6227 11064 6239 11067
rect 6730 11064 6736 11076
rect 6227 11036 6736 11064
rect 6227 11033 6239 11036
rect 6181 11027 6239 11033
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 6942 11073 7000 11079
rect 7043 11113 7101 11119
rect 7043 11079 7055 11113
rect 7089 11110 7101 11113
rect 7089 11079 7104 11110
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 7820 11135 7878 11141
rect 7820 11132 7832 11135
rect 7524 11104 7832 11132
rect 7524 11092 7530 11104
rect 7820 11101 7832 11104
rect 7866 11101 7878 11135
rect 7820 11095 7878 11101
rect 7926 11092 7932 11144
rect 7984 11141 7990 11144
rect 7984 11135 8027 11141
rect 8015 11101 8027 11135
rect 7984 11095 8027 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8220 11132 8248 11160
rect 8159 11104 8248 11132
rect 8389 11135 8447 11141
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 9214 11132 9220 11144
rect 8435 11104 9220 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 7984 11092 7990 11095
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 10134 11132 10140 11144
rect 9447 11104 10140 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10502 11132 10508 11144
rect 10284 11104 10329 11132
rect 10463 11104 10508 11132
rect 10284 11092 10290 11104
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 7043 11073 7104 11079
rect 6546 10996 6552 11008
rect 6012 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10996 6610 11008
rect 6822 10996 6828 11008
rect 6604 10968 6828 10996
rect 6604 10956 6610 10968
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 7076 10996 7104 11073
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 8205 11067 8263 11073
rect 7340 11036 8064 11064
rect 7340 11024 7346 11036
rect 7926 10996 7932 11008
rect 7076 10968 7932 10996
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8036 10996 8064 11036
rect 8205 11033 8217 11067
rect 8251 11033 8263 11067
rect 8754 11064 8760 11076
rect 8715 11036 8760 11064
rect 8205 11027 8263 11033
rect 8220 10996 8248 11027
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 8938 11064 8944 11076
rect 8899 11036 8944 11064
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9493 11067 9551 11073
rect 9493 11033 9505 11067
rect 9539 11033 9551 11067
rect 9674 11064 9680 11076
rect 9635 11036 9680 11064
rect 9493 11027 9551 11033
rect 9122 10996 9128 11008
rect 8036 10968 8248 10996
rect 9083 10968 9128 10996
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 9508 10996 9536 11027
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 9858 11064 9864 11076
rect 9819 11036 9864 11064
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 10042 11064 10048 11076
rect 10003 11036 10048 11064
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 10612 11064 10640 11172
rect 11054 11141 11060 11144
rect 11037 11135 11060 11141
rect 11037 11101 11049 11135
rect 11037 11095 11060 11101
rect 11054 11092 11060 11095
rect 11112 11092 11118 11144
rect 11164 11132 11192 11240
rect 11348 11240 11980 11268
rect 11348 11209 11376 11240
rect 11974 11228 11980 11240
rect 12032 11228 12038 11280
rect 12452 11277 12480 11308
rect 12437 11271 12495 11277
rect 12437 11237 12449 11271
rect 12483 11237 12495 11271
rect 12437 11231 12495 11237
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12986 11200 12992 11212
rect 12124 11172 12204 11200
rect 12124 11160 12130 11172
rect 11882 11132 11888 11144
rect 11164 11104 11652 11132
rect 11843 11104 11888 11132
rect 11624 11073 11652 11104
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12176 11141 12204 11172
rect 12406 11172 12992 11200
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11101 12219 11135
rect 12161 11095 12219 11101
rect 12305 11135 12363 11141
rect 12305 11101 12317 11135
rect 12351 11132 12363 11135
rect 12406 11132 12434 11172
rect 12986 11160 12992 11172
rect 13044 11160 13050 11212
rect 12618 11132 12624 11144
rect 12351 11104 12434 11132
rect 12579 11104 12624 11132
rect 12351 11101 12363 11104
rect 12305 11095 12363 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 13320 11104 13369 11132
rect 13320 11092 13326 11104
rect 13357 11101 13369 11104
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 10612 11036 10793 11064
rect 10781 11033 10793 11036
rect 10827 11033 10839 11067
rect 10781 11027 10839 11033
rect 11609 11067 11667 11073
rect 11609 11033 11621 11067
rect 11655 11033 11667 11067
rect 11790 11064 11796 11076
rect 11751 11036 11796 11064
rect 11609 11027 11667 11033
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 12066 11064 12072 11076
rect 12027 11036 12072 11064
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 13078 11064 13084 11076
rect 13039 11036 13084 11064
rect 13078 11024 13084 11036
rect 13136 11024 13142 11076
rect 13173 11067 13231 11073
rect 13173 11033 13185 11067
rect 13219 11064 13231 11067
rect 13630 11064 13636 11076
rect 13219 11036 13636 11064
rect 13219 11033 13231 11036
rect 13173 11027 13231 11033
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 9582 10996 9588 11008
rect 9508 10968 9588 10996
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 10376 10968 10425 10996
rect 10376 10956 10382 10968
rect 10413 10965 10425 10968
rect 10459 10965 10471 10999
rect 10413 10959 10471 10965
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 11149 10999 11207 11005
rect 11149 10996 11161 10999
rect 10652 10968 11161 10996
rect 10652 10956 10658 10968
rect 11149 10965 11161 10968
rect 11195 10965 11207 10999
rect 11149 10959 11207 10965
rect 11241 10999 11299 11005
rect 11241 10965 11253 10999
rect 11287 10996 11299 10999
rect 11330 10996 11336 11008
rect 11287 10968 11336 10996
rect 11287 10965 11299 10968
rect 11241 10959 11299 10965
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13449 10999 13507 11005
rect 13449 10996 13461 10999
rect 13412 10968 13461 10996
rect 13412 10956 13418 10968
rect 13449 10965 13461 10968
rect 13495 10965 13507 10999
rect 13449 10959 13507 10965
rect 1104 10906 13892 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 13892 10906
rect 1104 10832 13892 10854
rect 3694 10752 3700 10804
rect 3752 10752 3758 10804
rect 5350 10792 5356 10804
rect 3804 10764 5356 10792
rect 3421 10727 3479 10733
rect 3421 10693 3433 10727
rect 3467 10724 3479 10727
rect 3712 10724 3740 10752
rect 3467 10696 3740 10724
rect 3467 10693 3479 10696
rect 3421 10687 3479 10693
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 2314 10656 2320 10668
rect 1443 10628 2320 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2866 10656 2872 10668
rect 2731 10628 2872 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 3326 10665 3332 10668
rect 3324 10656 3332 10665
rect 3287 10628 3332 10656
rect 3324 10619 3332 10628
rect 3326 10616 3332 10619
rect 3384 10616 3390 10668
rect 3510 10656 3516 10668
rect 3471 10628 3516 10656
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3602 10616 3608 10668
rect 3660 10656 3666 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3660 10628 3709 10656
rect 3660 10616 3666 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 566 10548 572 10600
rect 624 10588 630 10600
rect 624 10560 3280 10588
rect 624 10548 630 10560
rect 2682 10520 2688 10532
rect 2643 10492 2688 10520
rect 2682 10480 2688 10492
rect 2740 10480 2746 10532
rect 3252 10520 3280 10560
rect 3804 10529 3832 10764
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6512 10764 6561 10792
rect 6512 10752 6518 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 6549 10755 6607 10761
rect 7300 10764 7972 10792
rect 4249 10727 4307 10733
rect 4249 10693 4261 10727
rect 4295 10724 4307 10727
rect 4890 10724 4896 10736
rect 4295 10696 4896 10724
rect 4295 10693 4307 10696
rect 4249 10687 4307 10693
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 4264 10656 4292 10687
rect 4890 10684 4896 10696
rect 4948 10684 4954 10736
rect 5258 10724 5264 10736
rect 5219 10696 5264 10724
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 7193 10727 7251 10733
rect 7193 10724 7205 10727
rect 6012 10696 7205 10724
rect 4019 10628 4292 10656
rect 4525 10659 4583 10665
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5810 10656 5816 10668
rect 5215 10628 5816 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 4540 10588 4568 10619
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 5353 10591 5411 10597
rect 5353 10588 5365 10591
rect 4540 10560 5365 10588
rect 5353 10557 5365 10560
rect 5399 10588 5411 10591
rect 6012 10588 6040 10696
rect 7193 10693 7205 10696
rect 7239 10693 7251 10727
rect 7193 10687 7251 10693
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 6144 10628 6193 10656
rect 6144 10616 6150 10628
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6270 10616 6276 10668
rect 6328 10656 6334 10668
rect 6661 10659 6719 10665
rect 6661 10656 6673 10659
rect 6328 10628 6673 10656
rect 6328 10616 6334 10628
rect 6661 10625 6673 10628
rect 6707 10625 6719 10659
rect 6661 10619 6719 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7300 10656 7328 10764
rect 7944 10724 7972 10764
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 8168 10764 8401 10792
rect 8168 10752 8174 10764
rect 8389 10761 8401 10764
rect 8435 10761 8447 10795
rect 8389 10755 8447 10761
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8536 10764 9720 10792
rect 8536 10752 8542 10764
rect 9490 10724 9496 10736
rect 7944 10696 9496 10724
rect 9490 10684 9496 10696
rect 9548 10684 9554 10736
rect 7147 10628 7328 10656
rect 7837 10659 7895 10665
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 5399 10560 6040 10588
rect 6365 10591 6423 10597
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 6365 10557 6377 10591
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 6457 10591 6515 10597
rect 6457 10557 6469 10591
rect 6503 10588 6515 10591
rect 6546 10588 6552 10600
rect 6503 10560 6552 10588
rect 6503 10557 6515 10560
rect 6457 10551 6515 10557
rect 3789 10523 3847 10529
rect 3789 10520 3801 10523
rect 3252 10492 3801 10520
rect 3789 10489 3801 10492
rect 3835 10489 3847 10523
rect 3789 10483 3847 10489
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 5258 10520 5264 10532
rect 4203 10492 5264 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 6380 10520 6408 10551
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 6932 10588 6960 10619
rect 7374 10588 7380 10600
rect 6932 10560 7380 10588
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 7852 10588 7880 10619
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8555 10659 8613 10665
rect 8555 10656 8567 10659
rect 7984 10628 8029 10656
rect 8312 10628 8567 10656
rect 7984 10616 7990 10628
rect 7800 10560 7880 10588
rect 6914 10520 6920 10532
rect 6380 10492 6920 10520
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 7800 10520 7828 10560
rect 8018 10548 8024 10600
rect 8076 10588 8082 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 8076 10560 8217 10588
rect 8076 10548 8082 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8110 10520 8116 10532
rect 7156 10492 7828 10520
rect 8071 10492 8116 10520
rect 7156 10480 7162 10492
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 3108 10424 3157 10452
rect 3108 10412 3114 10424
rect 3145 10421 3157 10424
rect 3191 10421 3203 10455
rect 3145 10415 3203 10421
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 5997 10455 6055 10461
rect 5997 10452 6009 10455
rect 3568 10424 6009 10452
rect 3568 10412 3574 10424
rect 5997 10421 6009 10424
rect 6043 10452 6055 10455
rect 6454 10452 6460 10464
rect 6043 10424 6460 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 6788 10424 7297 10452
rect 6788 10412 6794 10424
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 7285 10415 7343 10421
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 7653 10455 7711 10461
rect 7653 10452 7665 10455
rect 7524 10424 7665 10452
rect 7524 10412 7530 10424
rect 7653 10421 7665 10424
rect 7699 10421 7711 10455
rect 7800 10452 7828 10492
rect 8110 10480 8116 10492
rect 8168 10520 8174 10532
rect 8312 10520 8340 10628
rect 8555 10625 8567 10628
rect 8601 10625 8613 10659
rect 8555 10619 8613 10625
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 8680 10588 8708 10619
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 9088 10628 9137 10656
rect 9088 10616 9094 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9308 10659 9366 10665
rect 9308 10625 9320 10659
rect 9354 10656 9366 10659
rect 9582 10656 9588 10668
rect 9354 10628 9588 10656
rect 9354 10625 9366 10628
rect 9308 10619 9366 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 9692 10665 9720 10764
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10100 10764 10149 10792
rect 10100 10752 10106 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10137 10755 10195 10761
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 10744 10764 11100 10792
rect 10744 10752 10750 10764
rect 9941 10727 9999 10733
rect 9941 10693 9953 10727
rect 9987 10693 9999 10727
rect 10962 10724 10968 10736
rect 10923 10696 10968 10724
rect 9941 10687 9999 10693
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 9944 10600 9972 10687
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 11072 10724 11100 10764
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11330 10792 11336 10804
rect 11204 10764 11336 10792
rect 11204 10752 11210 10764
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11480 10764 11744 10792
rect 11480 10752 11486 10764
rect 11072 10696 11192 10724
rect 10594 10656 10600 10668
rect 10432 10628 10600 10656
rect 8938 10588 8944 10600
rect 8444 10560 8708 10588
rect 8899 10560 8944 10588
rect 8444 10548 8450 10560
rect 8168 10492 8340 10520
rect 8680 10520 8708 10560
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10557 9551 10591
rect 9944 10560 9956 10600
rect 9493 10551 9551 10557
rect 9416 10520 9444 10551
rect 8680 10492 9444 10520
rect 8168 10480 8174 10492
rect 8294 10452 8300 10464
rect 7800 10424 8300 10452
rect 7653 10415 7711 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 8849 10455 8907 10461
rect 8849 10452 8861 10455
rect 8444 10424 8861 10452
rect 8444 10412 8450 10424
rect 8849 10421 8861 10424
rect 8895 10452 8907 10455
rect 9122 10452 9128 10464
rect 8895 10424 9128 10452
rect 8895 10421 8907 10424
rect 8849 10415 8907 10421
rect 9122 10412 9128 10424
rect 9180 10452 9186 10464
rect 9508 10452 9536 10551
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 9861 10523 9919 10529
rect 9861 10489 9873 10523
rect 9907 10520 9919 10523
rect 10432 10520 10460 10628
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 10686 10616 10692 10668
rect 10744 10665 10750 10668
rect 11164 10665 11192 10696
rect 11716 10665 11744 10764
rect 12158 10724 12164 10736
rect 11808 10696 12164 10724
rect 10744 10659 10787 10665
rect 10775 10625 10787 10659
rect 10744 10619 10787 10625
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10656 10931 10659
rect 11149 10659 11207 10665
rect 10919 10646 11008 10656
rect 10919 10628 11083 10646
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 10744 10616 10750 10619
rect 10980 10618 11083 10628
rect 11149 10625 11161 10659
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11055 10588 11083 10618
rect 11808 10588 11836 10696
rect 12158 10684 12164 10696
rect 12216 10684 12222 10736
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 11055 10560 11836 10588
rect 11900 10588 11928 10619
rect 11974 10616 11980 10668
rect 12032 10656 12038 10668
rect 12618 10656 12624 10668
rect 12032 10628 12624 10656
rect 12032 10616 12038 10628
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 13354 10656 13360 10668
rect 13315 10628 13360 10656
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 12066 10588 12072 10600
rect 11900 10560 12072 10588
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 10594 10520 10600 10532
rect 9907 10492 10460 10520
rect 10555 10492 10600 10520
rect 9907 10489 9919 10492
rect 9861 10483 9919 10489
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 11054 10480 11060 10532
rect 11112 10520 11118 10532
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 11112 10492 11253 10520
rect 11112 10480 11118 10492
rect 11241 10489 11253 10492
rect 11287 10489 11299 10523
rect 11241 10483 11299 10489
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 13078 10520 13084 10532
rect 11388 10492 13084 10520
rect 11388 10480 11394 10492
rect 13078 10480 13084 10492
rect 13136 10520 13142 10532
rect 13265 10523 13323 10529
rect 13265 10520 13277 10523
rect 13136 10492 13277 10520
rect 13136 10480 13142 10492
rect 13265 10489 13277 10492
rect 13311 10489 13323 10523
rect 13265 10483 13323 10489
rect 9180 10424 9536 10452
rect 9180 10412 9186 10424
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 9732 10424 10149 10452
rect 9732 10412 9738 10424
rect 10137 10421 10149 10424
rect 10183 10421 10195 10455
rect 10137 10415 10195 10421
rect 10321 10455 10379 10461
rect 10321 10421 10333 10455
rect 10367 10452 10379 10455
rect 11146 10452 11152 10464
rect 10367 10424 11152 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11422 10412 11428 10464
rect 11480 10452 11486 10464
rect 11609 10455 11667 10461
rect 11609 10452 11621 10455
rect 11480 10424 11621 10452
rect 11480 10412 11486 10424
rect 11609 10421 11621 10424
rect 11655 10421 11667 10455
rect 11609 10415 11667 10421
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 13170 10452 13176 10464
rect 11848 10424 13176 10452
rect 11848 10412 11854 10424
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 1104 10362 13892 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 13892 10362
rect 1104 10288 13892 10310
rect 6270 10248 6276 10260
rect 2700 10220 6276 10248
rect 2700 10056 2728 10220
rect 6270 10208 6276 10220
rect 6328 10208 6334 10260
rect 6454 10248 6460 10260
rect 6415 10220 6460 10248
rect 6454 10208 6460 10220
rect 6512 10248 6518 10260
rect 8110 10248 8116 10260
rect 6512 10220 8116 10248
rect 6512 10208 6518 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8352 10220 8708 10248
rect 8352 10208 8358 10220
rect 5074 10180 5080 10192
rect 5035 10152 5080 10180
rect 5074 10140 5080 10152
rect 5132 10140 5138 10192
rect 5718 10180 5724 10192
rect 5679 10152 5724 10180
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 7558 10180 7564 10192
rect 6236 10152 7564 10180
rect 6236 10140 6242 10152
rect 7558 10140 7564 10152
rect 7616 10180 7622 10192
rect 8478 10180 8484 10192
rect 7616 10152 8484 10180
rect 7616 10140 7622 10152
rect 8478 10140 8484 10152
rect 8536 10140 8542 10192
rect 8570 10140 8576 10192
rect 8628 10140 8634 10192
rect 8680 10180 8708 10220
rect 9122 10208 9128 10260
rect 9180 10248 9186 10260
rect 9493 10251 9551 10257
rect 9180 10220 9444 10248
rect 9180 10208 9186 10220
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 8680 10152 9045 10180
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 9416 10180 9444 10220
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 9674 10248 9680 10260
rect 9539 10220 9680 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 9861 10251 9919 10257
rect 9861 10217 9873 10251
rect 9907 10248 9919 10251
rect 10042 10248 10048 10260
rect 9907 10220 10048 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 11164 10220 12388 10248
rect 11164 10180 11192 10220
rect 9416 10152 11192 10180
rect 11241 10183 11299 10189
rect 9033 10143 9091 10149
rect 11241 10149 11253 10183
rect 11287 10180 11299 10183
rect 11287 10152 12296 10180
rect 11287 10149 11299 10152
rect 11241 10143 11299 10149
rect 5166 10112 5172 10124
rect 3344 10084 5172 10112
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10044 1547 10047
rect 1765 10047 1823 10053
rect 1765 10044 1777 10047
rect 1535 10016 1777 10044
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 1765 10013 1777 10016
rect 1811 10044 1823 10047
rect 2682 10044 2688 10056
rect 1811 10016 2176 10044
rect 2595 10016 2688 10044
rect 1811 10013 1823 10016
rect 1765 10007 1823 10013
rect 1946 9976 1952 9988
rect 1907 9948 1952 9976
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 2148 9976 2176 10016
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3234 10044 3240 10056
rect 2823 10016 3240 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3344 10053 3372 10084
rect 5166 10072 5172 10084
rect 5224 10112 5230 10124
rect 6362 10112 6368 10124
rect 5224 10084 6368 10112
rect 5224 10072 5230 10084
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10044 3571 10047
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3559 10016 3801 10044
rect 3559 10013 3571 10016
rect 3513 10007 3571 10013
rect 3789 10013 3801 10016
rect 3835 10044 3847 10047
rect 3970 10044 3976 10056
rect 3835 10016 3976 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4890 10044 4896 10056
rect 4851 10016 4896 10044
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 5902 10044 5908 10056
rect 5863 10016 5908 10044
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 6196 10053 6224 10084
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 7282 10112 7288 10124
rect 6472 10084 7288 10112
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6472 10044 6500 10084
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 6328 10016 6500 10044
rect 6733 10047 6791 10053
rect 6328 10004 6334 10016
rect 6733 10013 6745 10047
rect 6779 10044 6791 10047
rect 6822 10044 6828 10056
rect 6779 10016 6828 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 7135 10047 7193 10053
rect 6917 10007 6975 10013
rect 7010 10025 7068 10031
rect 2866 9976 2872 9988
rect 2148 9948 2872 9976
rect 2866 9936 2872 9948
rect 2924 9936 2930 9988
rect 3053 9979 3111 9985
rect 3053 9945 3065 9979
rect 3099 9976 3111 9979
rect 6086 9976 6092 9988
rect 3099 9948 3280 9976
rect 6047 9948 6092 9976
rect 3099 9945 3111 9948
rect 3053 9939 3111 9945
rect 3252 9920 3280 9948
rect 6086 9936 6092 9948
rect 6144 9936 6150 9988
rect 6457 9979 6515 9985
rect 6457 9945 6469 9979
rect 6503 9976 6515 9979
rect 6546 9976 6552 9988
rect 6503 9948 6552 9976
rect 6503 9945 6515 9948
rect 6457 9939 6515 9945
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 6638 9936 6644 9988
rect 6696 9976 6702 9988
rect 6696 9948 6741 9976
rect 6696 9936 6702 9948
rect 1670 9908 1676 9920
rect 1631 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 2958 9908 2964 9920
rect 2919 9880 2964 9908
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 3142 9908 3148 9920
rect 3103 9880 3148 9908
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 3234 9868 3240 9920
rect 3292 9868 3298 9920
rect 5442 9908 5448 9920
rect 5403 9880 5448 9908
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6932 9908 6960 10007
rect 7010 9991 7022 10025
rect 7056 9991 7068 10025
rect 7135 10013 7147 10047
rect 7181 10044 7193 10047
rect 7558 10044 7564 10056
rect 7181 10016 7564 10044
rect 7181 10013 7193 10016
rect 7135 10007 7193 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8202 10044 8208 10056
rect 7984 10016 8208 10044
rect 7984 10004 7990 10016
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8386 10044 8392 10056
rect 8347 10016 8392 10044
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8478 10038 8484 10090
rect 8536 10038 8542 10090
rect 8588 10053 8616 10140
rect 9858 10072 9864 10124
rect 9916 10112 9922 10124
rect 10042 10112 10048 10124
rect 9916 10084 10048 10112
rect 9916 10072 9922 10084
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10134 10072 10140 10124
rect 10192 10112 10198 10124
rect 10962 10112 10968 10124
rect 10192 10084 10968 10112
rect 10192 10072 10198 10084
rect 8573 10047 8631 10053
rect 8481 10013 8493 10038
rect 8527 10013 8539 10038
rect 8481 10007 8539 10013
rect 8573 10013 8585 10047
rect 8619 10013 8631 10047
rect 8941 10047 8999 10053
rect 8941 10046 8953 10047
rect 8573 10007 8631 10013
rect 8752 10018 8953 10046
rect 7010 9988 7068 9991
rect 7006 9936 7012 9988
rect 7064 9936 7070 9988
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 7377 9979 7435 9985
rect 7377 9976 7389 9979
rect 7340 9948 7389 9976
rect 7340 9936 7346 9948
rect 7377 9945 7389 9948
rect 7423 9945 7435 9979
rect 7377 9939 7435 9945
rect 8021 9979 8079 9985
rect 8021 9945 8033 9979
rect 8067 9976 8079 9979
rect 8110 9976 8116 9988
rect 8067 9948 8116 9976
rect 8067 9945 8079 9948
rect 8021 9939 8079 9945
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 8220 9976 8248 10004
rect 8752 9976 8780 10018
rect 8941 10013 8953 10018
rect 8987 10013 8999 10047
rect 9217 10047 9275 10053
rect 9217 10022 9229 10047
rect 8941 10007 8999 10013
rect 9140 10013 9229 10022
rect 9263 10013 9275 10047
rect 9140 10007 9275 10013
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 9582 10044 9588 10056
rect 9355 10016 9588 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 9140 9994 9260 10007
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 10336 10053 10364 10084
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10044 10011 10047
rect 10321 10047 10379 10053
rect 9999 10016 10272 10044
rect 9999 10013 10011 10016
rect 9953 10007 10011 10013
rect 8220 9948 8780 9976
rect 9030 9936 9036 9988
rect 9088 9976 9094 9988
rect 9140 9976 9168 9994
rect 10137 9979 10195 9985
rect 10137 9976 10149 9979
rect 9088 9948 9168 9976
rect 9324 9948 10149 9976
rect 9088 9936 9094 9948
rect 9324 9920 9352 9948
rect 10137 9945 10149 9948
rect 10183 9945 10195 9979
rect 10137 9939 10195 9945
rect 5776 9880 6960 9908
rect 5776 9868 5782 9880
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 7558 9908 7564 9920
rect 7248 9880 7564 9908
rect 7248 9868 7254 9880
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 8757 9911 8815 9917
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 9122 9908 9128 9920
rect 8803 9880 9128 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9306 9868 9312 9920
rect 9364 9868 9370 9920
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 10244 9908 10272 10016
rect 10321 10013 10333 10047
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10686 10044 10692 10056
rect 10647 10016 10692 10044
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 10888 10053 10916 10084
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 11974 10112 11980 10124
rect 11532 10084 11980 10112
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 11109 10047 11167 10053
rect 11109 10013 11121 10047
rect 11155 10044 11167 10047
rect 11532 10044 11560 10084
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 11155 10016 11560 10044
rect 11155 10013 11167 10016
rect 11109 10007 11167 10013
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11664 10016 11713 10044
rect 11664 10004 11670 10016
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 12268 10044 12296 10152
rect 12360 10112 12388 10220
rect 13170 10208 13176 10260
rect 13228 10248 13234 10260
rect 13265 10251 13323 10257
rect 13265 10248 13277 10251
rect 13228 10220 13277 10248
rect 13228 10208 13234 10220
rect 13265 10217 13277 10220
rect 13311 10217 13323 10251
rect 13265 10211 13323 10217
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 12360 10084 12541 10112
rect 12529 10081 12541 10084
rect 12575 10081 12587 10115
rect 13081 10115 13139 10121
rect 13081 10112 13093 10115
rect 12529 10075 12587 10081
rect 12636 10084 13093 10112
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 12268 10016 12449 10044
rect 11701 10007 11759 10013
rect 12437 10013 12449 10016
rect 12483 10044 12495 10047
rect 12636 10044 12664 10084
rect 13081 10081 13093 10084
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 12483 10016 12664 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 10428 9976 10456 10004
rect 10594 9976 10600 9988
rect 10428 9948 10600 9976
rect 10594 9936 10600 9948
rect 10652 9936 10658 9988
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 10965 9979 11023 9985
rect 10965 9976 10977 9979
rect 10836 9948 10977 9976
rect 10836 9936 10842 9948
rect 10965 9945 10977 9948
rect 11011 9945 11023 9979
rect 10965 9939 11023 9945
rect 11422 9936 11428 9988
rect 11480 9976 11486 9988
rect 11517 9979 11575 9985
rect 11517 9976 11529 9979
rect 11480 9948 11529 9976
rect 11480 9936 11486 9948
rect 11517 9945 11529 9948
rect 11563 9945 11575 9979
rect 11716 9976 11744 10007
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12768 10016 13185 10044
rect 12768 10004 12774 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 12621 9979 12679 9985
rect 12621 9976 12633 9979
rect 11716 9948 12633 9976
rect 11517 9939 11575 9945
rect 12621 9945 12633 9948
rect 12667 9945 12679 9979
rect 12621 9939 12679 9945
rect 12894 9936 12900 9988
rect 12952 9976 12958 9988
rect 13372 9976 13400 10007
rect 12952 9948 13400 9976
rect 12952 9936 12958 9948
rect 10100 9880 10272 9908
rect 10100 9868 10106 9880
rect 10410 9868 10416 9920
rect 10468 9908 10474 9920
rect 10505 9911 10563 9917
rect 10505 9908 10517 9911
rect 10468 9880 10517 9908
rect 10468 9868 10474 9880
rect 10505 9877 10517 9880
rect 10551 9877 10563 9911
rect 10505 9871 10563 9877
rect 10686 9868 10692 9920
rect 10744 9908 10750 9920
rect 12434 9908 12440 9920
rect 10744 9880 12440 9908
rect 10744 9868 10750 9880
rect 12434 9868 12440 9880
rect 12492 9868 12498 9920
rect 1104 9818 13892 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 13892 9818
rect 1104 9744 13892 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 3476 9676 4629 9704
rect 3476 9664 3482 9676
rect 4617 9673 4629 9676
rect 4663 9673 4675 9707
rect 4890 9704 4896 9716
rect 4851 9676 4896 9704
rect 4617 9667 4675 9673
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 5997 9707 6055 9713
rect 5997 9673 6009 9707
rect 6043 9704 6055 9707
rect 6546 9704 6552 9716
rect 6043 9676 6552 9704
rect 6043 9673 6055 9676
rect 5997 9667 6055 9673
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 7653 9707 7711 9713
rect 7653 9673 7665 9707
rect 7699 9704 7711 9707
rect 7834 9704 7840 9716
rect 7699 9676 7840 9704
rect 7699 9673 7711 9676
rect 7653 9667 7711 9673
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 8110 9704 8116 9716
rect 8071 9676 8116 9704
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8573 9707 8631 9713
rect 8220 9676 8524 9704
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 1857 9639 1915 9645
rect 1857 9636 1869 9639
rect 1728 9608 1869 9636
rect 1728 9596 1734 9608
rect 1857 9605 1869 9608
rect 1903 9605 1915 9639
rect 1857 9599 1915 9605
rect 1946 9596 1952 9648
rect 2004 9636 2010 9648
rect 2004 9608 2049 9636
rect 2004 9596 2010 9608
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 3145 9639 3203 9645
rect 3145 9636 3157 9639
rect 2924 9608 3157 9636
rect 2924 9596 2930 9608
rect 3145 9605 3157 9608
rect 3191 9605 3203 9639
rect 3145 9599 3203 9605
rect 3789 9639 3847 9645
rect 3789 9605 3801 9639
rect 3835 9636 3847 9639
rect 4433 9639 4491 9645
rect 4433 9636 4445 9639
rect 3835 9608 4445 9636
rect 3835 9605 3847 9608
rect 3789 9599 3847 9605
rect 4433 9605 4445 9608
rect 4479 9636 4491 9639
rect 5074 9636 5080 9648
rect 4479 9608 5080 9636
rect 4479 9605 4491 9608
rect 4433 9599 4491 9605
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5169 9639 5227 9645
rect 5169 9605 5181 9639
rect 5215 9636 5227 9639
rect 5442 9636 5448 9648
rect 5215 9608 5448 9636
rect 5215 9605 5227 9608
rect 5169 9599 5227 9605
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 6362 9636 6368 9648
rect 6323 9608 6368 9636
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 6638 9596 6644 9648
rect 6696 9636 6702 9648
rect 7282 9636 7288 9648
rect 6696 9608 6868 9636
rect 7243 9608 7288 9636
rect 6696 9596 6702 9608
rect 1762 9568 1768 9580
rect 1723 9540 1768 9568
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2148 9540 2513 9568
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 2148 9500 2176 9540
rect 2501 9537 2513 9540
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 2639 9540 3341 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 3329 9537 3341 9540
rect 3375 9568 3387 9571
rect 3418 9568 3424 9580
rect 3375 9540 3424 9568
rect 3375 9537 3387 9540
rect 3329 9531 3387 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 3970 9568 3976 9580
rect 3931 9540 3976 9568
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 4890 9528 4896 9580
rect 4948 9568 4954 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4948 9540 4997 9568
rect 4948 9528 4954 9540
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9568 5779 9571
rect 5994 9568 6000 9580
rect 5767 9540 6000 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 6454 9568 6460 9580
rect 6227 9540 6460 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6454 9528 6460 9540
rect 6512 9568 6518 9580
rect 6840 9577 6868 9608
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 7469 9639 7527 9645
rect 7469 9605 7481 9639
rect 7515 9636 7527 9639
rect 8220 9636 8248 9676
rect 7515 9608 7880 9636
rect 7515 9605 7527 9608
rect 7469 9599 7527 9605
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6512 9540 6561 9568
rect 6512 9528 6518 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 6951 9571 7009 9577
rect 6951 9537 6963 9571
rect 6997 9568 7009 9571
rect 7098 9568 7104 9580
rect 6997 9540 7104 9568
rect 6997 9537 7009 9540
rect 6951 9531 7009 9537
rect 1719 9472 2176 9500
rect 2409 9503 2467 9509
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2409 9469 2421 9503
rect 2455 9500 2467 9503
rect 2682 9500 2688 9512
rect 2455 9472 2688 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 3050 9500 3056 9512
rect 3011 9472 3056 9500
rect 3050 9460 3056 9472
rect 3108 9460 3114 9512
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 4571 9472 5948 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 3605 9435 3663 9441
rect 3605 9432 3617 9435
rect 3384 9404 3617 9432
rect 3384 9392 3390 9404
rect 3605 9401 3617 9404
rect 3651 9401 3663 9435
rect 5258 9432 5264 9444
rect 5219 9404 5264 9432
rect 3605 9395 3663 9401
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 5920 9432 5948 9472
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 6748 9500 6776 9531
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7852 9577 7880 9608
rect 8036 9608 8248 9636
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9537 7895 9571
rect 7837 9531 7895 9537
rect 6144 9472 6868 9500
rect 6144 9460 6150 9472
rect 6840 9444 6868 9472
rect 6730 9432 6736 9444
rect 5920 9404 6736 9432
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 6822 9392 6828 9444
rect 6880 9392 6886 9444
rect 7193 9435 7251 9441
rect 7193 9401 7205 9435
rect 7239 9432 7251 9435
rect 8036 9432 8064 9608
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 8496 9636 8524 9676
rect 8573 9673 8585 9707
rect 8619 9704 8631 9707
rect 8938 9704 8944 9716
rect 8619 9676 8944 9704
rect 8619 9673 8631 9676
rect 8573 9667 8631 9673
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 9950 9704 9956 9716
rect 9048 9676 9956 9704
rect 9048 9636 9076 9676
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10045 9707 10103 9713
rect 10045 9673 10057 9707
rect 10091 9704 10103 9707
rect 10226 9704 10232 9716
rect 10091 9676 10232 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 11624 9676 11836 9704
rect 11624 9648 11652 9676
rect 8352 9608 8397 9636
rect 8496 9608 9076 9636
rect 9217 9639 9275 9645
rect 8352 9596 8358 9608
rect 9217 9605 9229 9639
rect 9263 9636 9275 9639
rect 9263 9608 10272 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 8386 9568 8392 9580
rect 8347 9540 8392 9568
rect 8386 9528 8392 9540
rect 8444 9568 8450 9580
rect 8754 9568 8760 9580
rect 8444 9540 8760 9568
rect 8444 9528 8450 9540
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 8941 9571 8999 9577
rect 8941 9537 8953 9571
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 8294 9460 8300 9512
rect 8352 9500 8358 9512
rect 8956 9500 8984 9531
rect 9122 9528 9128 9580
rect 9180 9568 9186 9580
rect 9309 9571 9367 9577
rect 9309 9568 9321 9571
rect 9180 9540 9321 9568
rect 9180 9528 9186 9540
rect 9309 9537 9321 9540
rect 9355 9537 9367 9571
rect 9582 9568 9588 9580
rect 9543 9540 9588 9568
rect 9309 9531 9367 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 9766 9528 9772 9580
rect 9824 9577 9830 9580
rect 9950 9577 9956 9580
rect 9824 9571 9873 9577
rect 9824 9537 9827 9571
rect 9861 9537 9873 9571
rect 9824 9531 9873 9537
rect 9929 9571 9956 9577
rect 9929 9537 9941 9571
rect 9929 9531 9956 9537
rect 9824 9528 9830 9531
rect 9950 9528 9956 9531
rect 10008 9528 10014 9580
rect 10244 9577 10272 9608
rect 10318 9596 10324 9648
rect 10376 9636 10382 9648
rect 10873 9639 10931 9645
rect 10376 9608 10456 9636
rect 10376 9596 10382 9608
rect 10428 9577 10456 9608
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 11054 9636 11060 9648
rect 10919 9608 11060 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 11296 9608 11529 9636
rect 11296 9596 11302 9608
rect 11517 9605 11529 9608
rect 11563 9605 11575 9639
rect 11517 9599 11575 9605
rect 11606 9596 11612 9648
rect 11664 9596 11670 9648
rect 11808 9636 11836 9676
rect 12345 9639 12403 9645
rect 12345 9636 12357 9639
rect 11808 9608 12357 9636
rect 12345 9605 12357 9608
rect 12391 9605 12403 9639
rect 12345 9599 12403 9605
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 10560 9540 10701 9568
rect 10560 9528 10566 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 11072 9568 11100 9596
rect 11333 9571 11391 9577
rect 11072 9540 11284 9568
rect 10689 9531 10747 9537
rect 8352 9472 8984 9500
rect 9033 9503 9091 9509
rect 8352 9460 8358 9472
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9674 9500 9680 9512
rect 9079 9472 9680 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9500 10195 9503
rect 11256 9500 11284 9540
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11422 9568 11428 9580
rect 11379 9540 11428 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 11698 9528 11704 9580
rect 11756 9568 11762 9580
rect 12069 9571 12127 9577
rect 12069 9568 12081 9571
rect 11756 9540 12081 9568
rect 11756 9528 11762 9540
rect 12069 9537 12081 9540
rect 12115 9568 12127 9571
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 12115 9540 12173 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 12161 9531 12219 9537
rect 12268 9540 13369 9568
rect 12268 9500 12296 9540
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 10183 9472 10460 9500
rect 11256 9472 12296 9500
rect 12713 9503 12771 9509
rect 10183 9469 10195 9472
rect 10137 9463 10195 9469
rect 8662 9432 8668 9444
rect 7239 9404 8064 9432
rect 8128 9404 8668 9432
rect 7239 9401 7251 9404
rect 7193 9395 7251 9401
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 7208 9364 7236 9395
rect 7466 9364 7472 9376
rect 1912 9336 7236 9364
rect 7427 9336 7472 9364
rect 1912 9324 1918 9336
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 8128 9373 8156 9404
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 10321 9435 10379 9441
rect 10321 9432 10333 9435
rect 8904 9404 10333 9432
rect 8904 9392 8910 9404
rect 10321 9401 10333 9404
rect 10367 9401 10379 9435
rect 10321 9395 10379 9401
rect 8116 9367 8174 9373
rect 8116 9333 8128 9367
rect 8162 9333 8174 9367
rect 8116 9327 8174 9333
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 8996 9336 9413 9364
rect 8996 9324 9002 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 10432 9364 10460 9472
rect 12713 9469 12725 9503
rect 12759 9500 12771 9503
rect 12802 9500 12808 9512
rect 12759 9472 12808 9500
rect 12759 9469 12771 9472
rect 12713 9463 12771 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 13262 9500 13268 9512
rect 13223 9472 13268 9500
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 11057 9435 11115 9441
rect 11057 9432 11069 9435
rect 10704 9404 11069 9432
rect 10704 9364 10732 9404
rect 11057 9401 11069 9404
rect 11103 9401 11115 9435
rect 11057 9395 11115 9401
rect 11146 9392 11152 9444
rect 11204 9432 11210 9444
rect 11609 9435 11667 9441
rect 11609 9432 11621 9435
rect 11204 9404 11621 9432
rect 11204 9392 11210 9404
rect 11609 9401 11621 9404
rect 11655 9401 11667 9435
rect 13170 9432 13176 9444
rect 13131 9404 13176 9432
rect 11609 9395 11667 9401
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 10432 9336 10732 9364
rect 9401 9327 9459 9333
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 10836 9336 11253 9364
rect 10836 9324 10842 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11241 9327 11299 9333
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12618 9364 12624 9376
rect 12483 9336 12624 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 1104 9274 13892 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 13892 9274
rect 1104 9200 13892 9222
rect 1762 9120 1768 9172
rect 1820 9160 1826 9172
rect 2682 9160 2688 9172
rect 1820 9132 2688 9160
rect 1820 9120 1826 9132
rect 2682 9120 2688 9132
rect 2740 9160 2746 9172
rect 3602 9160 3608 9172
rect 2740 9120 2774 9160
rect 3563 9132 3608 9160
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 6178 9160 6184 9172
rect 6139 9132 6184 9160
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6454 9160 6460 9172
rect 6415 9132 6460 9160
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 7098 9160 7104 9172
rect 6656 9132 7104 9160
rect 2746 9092 2774 9120
rect 6656 9101 6684 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 7708 9132 7757 9160
rect 7708 9120 7714 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 7745 9123 7803 9129
rect 7834 9120 7840 9172
rect 7892 9160 7898 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 7892 9132 7941 9160
rect 7892 9120 7898 9132
rect 7929 9129 7941 9132
rect 7975 9160 7987 9163
rect 8662 9160 8668 9172
rect 7975 9132 8668 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 8754 9120 8760 9172
rect 8812 9160 8818 9172
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 8812 9132 9965 9160
rect 8812 9120 8818 9132
rect 9953 9129 9965 9132
rect 9999 9129 10011 9163
rect 9953 9123 10011 9129
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 10100 9132 10241 9160
rect 10100 9120 10106 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 12802 9160 12808 9172
rect 10229 9123 10287 9129
rect 10520 9132 11192 9160
rect 12763 9132 12808 9160
rect 3881 9095 3939 9101
rect 3881 9092 3893 9095
rect 2746 9064 3893 9092
rect 3881 9061 3893 9064
rect 3927 9061 3939 9095
rect 3881 9055 3939 9061
rect 6641 9095 6699 9101
rect 6641 9061 6653 9095
rect 6687 9061 6699 9095
rect 6641 9055 6699 9061
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 7009 9095 7067 9101
rect 7009 9092 7021 9095
rect 6972 9064 7021 9092
rect 6972 9052 6978 9064
rect 7009 9061 7021 9064
rect 7055 9061 7067 9095
rect 7009 9055 7067 9061
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 7558 9092 7564 9104
rect 7248 9064 7564 9092
rect 7248 9052 7254 9064
rect 7558 9052 7564 9064
rect 7616 9092 7622 9104
rect 7616 9064 8432 9092
rect 7616 9052 7622 9064
rect 2774 9024 2780 9036
rect 1780 8996 2780 9024
rect 1780 8965 1808 8996
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3789 9027 3847 9033
rect 3789 9024 3801 9027
rect 3016 8996 3801 9024
rect 3016 8984 3022 8996
rect 3789 8993 3801 8996
rect 3835 8993 3847 9027
rect 3789 8987 3847 8993
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 4028 8996 4353 9024
rect 4028 8984 4034 8996
rect 4341 8993 4353 8996
rect 4387 9024 4399 9027
rect 4387 8996 8340 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8956 1915 8959
rect 3326 8956 3332 8968
rect 1903 8928 2774 8956
rect 3287 8928 3332 8956
rect 1903 8925 1915 8928
rect 1857 8919 1915 8925
rect 2746 8888 2774 8928
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 5077 8959 5135 8965
rect 4488 8928 4533 8956
rect 4488 8916 4494 8928
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5626 8956 5632 8968
rect 5123 8928 5632 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 5994 8956 6000 8968
rect 5955 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8956 6331 8959
rect 6822 8956 6828 8968
rect 6319 8928 6828 8956
rect 6319 8925 6331 8928
rect 6273 8919 6331 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7466 8956 7472 8968
rect 6932 8928 7472 8956
rect 3050 8888 3056 8900
rect 2746 8860 3056 8888
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 3418 8888 3424 8900
rect 3379 8860 3424 8888
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 4890 8888 4896 8900
rect 4851 8860 4896 8888
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 5258 8888 5264 8900
rect 5040 8860 5085 8888
rect 5171 8860 5264 8888
rect 5040 8848 5046 8860
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 6362 8848 6368 8900
rect 6420 8888 6426 8900
rect 6932 8897 6960 8928
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 7892 8928 7941 8956
rect 7892 8916 7898 8928
rect 7929 8925 7941 8928
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8168 8928 8213 8956
rect 8168 8916 8174 8928
rect 6917 8891 6975 8897
rect 6917 8888 6929 8891
rect 6420 8860 6929 8888
rect 6420 8848 6426 8860
rect 6917 8857 6929 8860
rect 6963 8857 6975 8891
rect 7190 8888 7196 8900
rect 7151 8860 7196 8888
rect 6917 8851 6975 8857
rect 7190 8848 7196 8860
rect 7248 8848 7254 8900
rect 7377 8891 7435 8897
rect 7377 8857 7389 8891
rect 7423 8857 7435 8891
rect 8312 8888 8340 8996
rect 8404 8965 8432 9064
rect 8496 9064 9260 9092
rect 8496 9033 8524 9064
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 8754 9024 8760 9036
rect 8481 8987 8539 8993
rect 8588 8996 8760 9024
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8588 8888 8616 8996
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9232 9024 9260 9064
rect 9490 9052 9496 9104
rect 9548 9092 9554 9104
rect 9585 9095 9643 9101
rect 9585 9092 9597 9095
rect 9548 9064 9597 9092
rect 9548 9052 9554 9064
rect 9585 9061 9597 9064
rect 9631 9061 9643 9095
rect 9585 9055 9643 9061
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 10520 9092 10548 9132
rect 11164 9104 11192 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 10686 9092 10692 9104
rect 9824 9064 10548 9092
rect 10647 9064 10692 9092
rect 9824 9052 9830 9064
rect 10686 9052 10692 9064
rect 10744 9052 10750 9104
rect 11146 9092 11152 9104
rect 11059 9064 11152 9092
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 9674 9024 9680 9036
rect 9232 8996 9680 9024
rect 8665 8959 8723 8965
rect 8665 8925 8677 8959
rect 8711 8956 8723 8959
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8711 8928 8953 8956
rect 8711 8925 8723 8928
rect 8665 8919 8723 8925
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9324 8965 9352 8996
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10704 9024 10732 9052
rect 10060 8996 10732 9024
rect 10060 8968 10088 8996
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 11296 8996 13369 9024
rect 11296 8984 11302 8996
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 9088 8928 9137 8956
rect 9088 8916 9094 8928
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9218 8959 9276 8965
rect 9218 8946 9230 8959
rect 9264 8946 9276 8959
rect 9324 8959 9384 8965
rect 9125 8919 9183 8925
rect 8312 8860 8616 8888
rect 8757 8891 8815 8897
rect 9214 8894 9220 8946
rect 9272 8894 9278 8946
rect 9324 8928 9338 8959
rect 9326 8925 9338 8928
rect 9372 8925 9384 8959
rect 9858 8956 9864 8968
rect 9819 8928 9864 8956
rect 9326 8919 9384 8925
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 10042 8956 10048 8968
rect 9955 8928 10048 8956
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 10192 8928 10333 8956
rect 10192 8916 10198 8928
rect 10321 8925 10333 8928
rect 10367 8925 10379 8959
rect 10778 8956 10784 8968
rect 10739 8928 10784 8956
rect 10321 8919 10379 8925
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11054 8956 11060 8968
rect 11011 8928 11060 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11330 8956 11336 8968
rect 11291 8928 11336 8956
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 12618 8956 12624 8968
rect 12579 8928 12624 8956
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 7377 8851 7435 8857
rect 8757 8857 8769 8891
rect 8803 8888 8815 8891
rect 8803 8860 9168 8888
rect 8803 8857 8815 8860
rect 8757 8851 8815 8857
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 5276 8820 5304 8848
rect 2832 8792 5304 8820
rect 2832 8780 2838 8792
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 7392 8820 7420 8851
rect 8846 8820 8852 8832
rect 6696 8792 8852 8820
rect 6696 8780 6702 8792
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 9140 8820 9168 8860
rect 9322 8860 9812 8888
rect 9322 8820 9350 8860
rect 9140 8792 9350 8820
rect 9784 8820 9812 8860
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10505 8891 10563 8897
rect 10505 8888 10517 8891
rect 10008 8860 10517 8888
rect 10008 8848 10014 8860
rect 10505 8857 10517 8860
rect 10551 8888 10563 8891
rect 12066 8888 12072 8900
rect 10551 8860 12072 8888
rect 10551 8857 10563 8860
rect 10505 8851 10563 8857
rect 12066 8848 12072 8860
rect 12124 8848 12130 8900
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 13004 8888 13032 8919
rect 12584 8860 13032 8888
rect 13265 8891 13323 8897
rect 12584 8848 12590 8860
rect 13265 8857 13277 8891
rect 13311 8888 13323 8891
rect 13538 8888 13544 8900
rect 13311 8860 13544 8888
rect 13311 8857 13323 8860
rect 13265 8851 13323 8857
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 10042 8820 10048 8832
rect 9784 8792 10048 8820
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 13173 8823 13231 8829
rect 13173 8820 13185 8823
rect 10468 8792 13185 8820
rect 10468 8780 10474 8792
rect 13173 8789 13185 8792
rect 13219 8789 13231 8823
rect 13173 8783 13231 8789
rect 1104 8730 13892 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 13892 8730
rect 1104 8656 13892 8678
rect 2685 8619 2743 8625
rect 2685 8585 2697 8619
rect 2731 8616 2743 8619
rect 4982 8616 4988 8628
rect 2731 8588 4988 8616
rect 2731 8585 2743 8588
rect 2685 8579 2743 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 6549 8619 6607 8625
rect 6549 8585 6561 8619
rect 6595 8616 6607 8619
rect 7193 8619 7251 8625
rect 6595 8588 7052 8616
rect 6595 8585 6607 8588
rect 6549 8579 6607 8585
rect 2869 8551 2927 8557
rect 2869 8517 2881 8551
rect 2915 8548 2927 8551
rect 3326 8548 3332 8560
rect 2915 8520 3332 8548
rect 2915 8517 2927 8520
rect 2869 8511 2927 8517
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 7024 8548 7052 8588
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 7834 8616 7840 8628
rect 7239 8588 7840 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8481 8619 8539 8625
rect 8481 8585 8493 8619
rect 8527 8616 8539 8619
rect 8570 8616 8576 8628
rect 8527 8588 8576 8616
rect 8527 8585 8539 8588
rect 8481 8579 8539 8585
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 9030 8616 9036 8628
rect 8991 8588 9036 8616
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 9769 8619 9827 8625
rect 9769 8616 9781 8619
rect 9548 8588 9781 8616
rect 9548 8576 9554 8588
rect 9769 8585 9781 8588
rect 9815 8585 9827 8619
rect 9769 8579 9827 8585
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10284 8588 10885 8616
rect 10284 8576 10290 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 11020 8588 11253 8616
rect 11020 8576 11026 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 12710 8616 12716 8628
rect 11241 8579 11299 8585
rect 11624 8588 12716 8616
rect 7282 8548 7288 8560
rect 7024 8520 7288 8548
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 7668 8520 7972 8548
rect 7668 8492 7696 8520
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 3053 8483 3111 8489
rect 2832 8452 2877 8480
rect 2832 8440 2838 8452
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8480 3847 8483
rect 3970 8480 3976 8492
rect 3835 8452 3976 8480
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 3068 8412 3096 8443
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4430 8480 4436 8492
rect 4111 8452 4436 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5626 8480 5632 8492
rect 5583 8452 5632 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5626 8440 5632 8452
rect 5684 8480 5690 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5684 8452 5825 8480
rect 5684 8440 5690 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 6362 8480 6368 8492
rect 6323 8452 6368 8480
rect 5997 8443 6055 8449
rect 6012 8412 6040 8443
rect 6362 8440 6368 8452
rect 6420 8480 6426 8492
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 6420 8452 6745 8480
rect 6420 8440 6426 8452
rect 6733 8449 6745 8452
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6880 8452 7389 8480
rect 6880 8440 6886 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7650 8480 7656 8492
rect 7611 8452 7656 8480
rect 7377 8443 7435 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 7834 8480 7840 8492
rect 7795 8452 7840 8480
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 7944 8489 7972 8520
rect 8110 8508 8116 8560
rect 8168 8548 8174 8560
rect 9398 8548 9404 8560
rect 8168 8520 9404 8548
rect 8168 8508 8174 8520
rect 8220 8489 8248 8520
rect 9398 8508 9404 8520
rect 9456 8508 9462 8560
rect 9858 8548 9864 8560
rect 9600 8520 9864 8548
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8570 8480 8576 8492
rect 8343 8452 8576 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 8754 8480 8760 8492
rect 8715 8452 8760 8480
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 9180 8452 9229 8480
rect 9180 8440 9186 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9490 8480 9496 8492
rect 9364 8452 9409 8480
rect 9451 8452 9496 8480
rect 9364 8440 9370 8452
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9600 8489 9628 8520
rect 9858 8508 9864 8520
rect 9916 8548 9922 8560
rect 9916 8520 11100 8548
rect 9916 8508 9922 8520
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 10686 8489 10692 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9732 8452 10149 8480
rect 9732 8440 9738 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10683 8443 10692 8489
rect 10744 8480 10750 8492
rect 10962 8480 10968 8492
rect 10744 8452 10783 8480
rect 10923 8452 10968 8480
rect 10686 8440 10692 8443
rect 10744 8440 10750 8452
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11072 8489 11100 8520
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 6086 8412 6092 8424
rect 2740 8384 3096 8412
rect 5999 8384 6092 8412
rect 2740 8372 2746 8384
rect 6086 8372 6092 8384
rect 6144 8412 6150 8424
rect 9766 8412 9772 8424
rect 6144 8384 9772 8412
rect 6144 8372 6150 8384
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 10042 8412 10048 8424
rect 10003 8384 10048 8412
rect 10042 8372 10048 8384
rect 10100 8412 10106 8424
rect 10318 8412 10324 8424
rect 10100 8384 10324 8412
rect 10100 8372 10106 8384
rect 10318 8372 10324 8384
rect 10376 8412 10382 8424
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 10376 8384 10609 8412
rect 10376 8372 10382 8384
rect 10597 8381 10609 8384
rect 10643 8412 10655 8415
rect 11532 8412 11560 8443
rect 10643 8384 11560 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 4890 8304 4896 8356
rect 4948 8344 4954 8356
rect 5353 8347 5411 8353
rect 5353 8344 5365 8347
rect 4948 8316 5365 8344
rect 4948 8304 4954 8316
rect 5353 8313 5365 8316
rect 5399 8313 5411 8347
rect 6914 8344 6920 8356
rect 6875 8316 6920 8344
rect 5353 8307 5411 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7745 8347 7803 8353
rect 7745 8313 7757 8347
rect 7791 8344 7803 8347
rect 8018 8344 8024 8356
rect 7791 8316 8024 8344
rect 7791 8313 7803 8316
rect 7745 8307 7803 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 9214 8304 9220 8356
rect 9272 8344 9278 8356
rect 11624 8344 11652 8588
rect 12710 8576 12716 8588
rect 12768 8616 12774 8628
rect 13446 8616 13452 8628
rect 12768 8588 13452 8616
rect 12768 8576 12774 8588
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 12299 8551 12357 8557
rect 12299 8548 12311 8551
rect 11992 8520 12311 8548
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 9272 8316 11652 8344
rect 9272 8304 9278 8316
rect 3234 8236 3240 8288
rect 3292 8276 3298 8288
rect 3881 8279 3939 8285
rect 3881 8276 3893 8279
rect 3292 8248 3893 8276
rect 3292 8236 3298 8248
rect 3881 8245 3893 8248
rect 3927 8276 3939 8279
rect 6362 8276 6368 8288
rect 3927 8248 6368 8276
rect 3927 8245 3939 8248
rect 3881 8239 3939 8245
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 8754 8276 8760 8288
rect 7524 8248 8760 8276
rect 7524 8236 7530 8248
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 9306 8276 9312 8288
rect 8996 8248 9312 8276
rect 8996 8236 9002 8248
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 10152 8285 10180 8316
rect 10520 8288 10548 8316
rect 11698 8304 11704 8356
rect 11756 8344 11762 8356
rect 11992 8344 12020 8520
rect 12299 8517 12311 8520
rect 12345 8548 12357 8551
rect 12894 8548 12900 8560
rect 12345 8520 12900 8548
rect 12345 8517 12357 8520
rect 12299 8511 12357 8517
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8480 12679 8483
rect 12802 8480 12808 8492
rect 12667 8452 12808 8480
rect 12667 8449 12679 8452
rect 12621 8443 12679 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 13170 8412 13176 8424
rect 12952 8384 13176 8412
rect 12952 8372 12958 8384
rect 13170 8372 13176 8384
rect 13228 8412 13234 8424
rect 13280 8412 13308 8443
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 13504 8452 13553 8480
rect 13504 8440 13510 8452
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 13228 8384 13308 8412
rect 13228 8372 13234 8384
rect 12066 8344 12072 8356
rect 11756 8316 12072 8344
rect 11756 8304 11762 8316
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 12158 8304 12164 8356
rect 12216 8344 12222 8356
rect 12802 8344 12808 8356
rect 12216 8316 12808 8344
rect 12216 8304 12222 8316
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 10137 8279 10195 8285
rect 10137 8245 10149 8279
rect 10183 8245 10195 8279
rect 10137 8239 10195 8245
rect 10226 8236 10232 8288
rect 10284 8276 10290 8288
rect 10321 8279 10379 8285
rect 10321 8276 10333 8279
rect 10284 8248 10333 8276
rect 10284 8236 10290 8248
rect 10321 8245 10333 8248
rect 10367 8245 10379 8279
rect 10321 8239 10379 8245
rect 10502 8236 10508 8288
rect 10560 8276 10566 8288
rect 10560 8248 10653 8276
rect 10560 8236 10566 8248
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 12253 8279 12311 8285
rect 12253 8276 12265 8279
rect 11112 8248 12265 8276
rect 11112 8236 11118 8248
rect 12253 8245 12265 8248
rect 12299 8276 12311 8279
rect 13722 8276 13728 8288
rect 12299 8248 13728 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 1104 8186 13892 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 13892 8186
rect 1104 8112 13892 8134
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3694 8072 3700 8084
rect 3467 8044 3700 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3694 8032 3700 8044
rect 3752 8032 3758 8084
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 4614 8072 4620 8084
rect 4387 8044 4620 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 9398 8072 9404 8084
rect 8720 8044 9404 8072
rect 8720 8032 8726 8044
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 10778 8072 10784 8084
rect 9907 8044 10784 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 10888 8044 12434 8072
rect 1670 8004 1676 8016
rect 1631 7976 1676 8004
rect 1670 7964 1676 7976
rect 1728 7964 1734 8016
rect 3712 7936 3740 8032
rect 3878 7964 3884 8016
rect 3936 8004 3942 8016
rect 3936 7976 5028 8004
rect 3936 7964 3942 7976
rect 3970 7936 3976 7948
rect 1596 7908 2360 7936
rect 1596 7880 1624 7908
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1688 7732 1716 7831
rect 1762 7828 1768 7880
rect 1820 7868 1826 7880
rect 1949 7871 2007 7877
rect 1949 7868 1961 7871
rect 1820 7840 1961 7868
rect 1820 7828 1826 7840
rect 1949 7837 1961 7840
rect 1995 7837 2007 7871
rect 2130 7868 2136 7880
rect 2091 7840 2136 7868
rect 1949 7831 2007 7837
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 2332 7877 2360 7908
rect 3160 7908 3976 7936
rect 3160 7877 3188 7908
rect 3970 7896 3976 7908
rect 4028 7936 4034 7948
rect 4028 7908 4108 7936
rect 4028 7896 4034 7908
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7837 2375 7871
rect 2501 7871 2559 7877
rect 2501 7868 2513 7871
rect 2317 7831 2375 7837
rect 2424 7840 2513 7868
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 1946 7732 1952 7744
rect 1688 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7732 2010 7744
rect 2424 7732 2452 7840
rect 2501 7837 2513 7840
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 2774 7760 2780 7812
rect 2832 7800 2838 7812
rect 2976 7800 3004 7831
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 3878 7868 3884 7880
rect 3292 7840 3337 7868
rect 3436 7840 3884 7868
rect 3292 7828 3298 7840
rect 3050 7800 3056 7812
rect 2832 7772 2877 7800
rect 2963 7772 3056 7800
rect 2832 7760 2838 7772
rect 3050 7760 3056 7772
rect 3108 7800 3114 7812
rect 3436 7800 3464 7840
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4080 7877 4108 7908
rect 4706 7896 4712 7948
rect 4764 7896 4770 7948
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4724 7868 4752 7896
rect 4571 7840 4752 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 5000 7877 5028 7976
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 8297 8007 8355 8013
rect 8297 8004 8309 8007
rect 7892 7976 8309 8004
rect 7892 7964 7898 7976
rect 8297 7973 8309 7976
rect 8343 8004 8355 8007
rect 9030 8004 9036 8016
rect 8343 7976 8598 8004
rect 8991 7976 9036 8004
rect 8343 7973 8355 7976
rect 8297 7967 8355 7973
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7936 7619 7939
rect 7650 7936 7656 7948
rect 7607 7908 7656 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 7650 7896 7656 7908
rect 7708 7936 7714 7948
rect 8570 7936 8598 7976
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9214 7964 9220 8016
rect 9272 8004 9278 8016
rect 10888 8004 10916 8044
rect 11238 8004 11244 8016
rect 9272 7976 10916 8004
rect 11199 7976 11244 8004
rect 9272 7964 9278 7976
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 12161 8007 12219 8013
rect 12161 8004 12173 8007
rect 12032 7976 12173 8004
rect 12032 7964 12038 7976
rect 12161 7973 12173 7976
rect 12207 7973 12219 8007
rect 12406 8004 12434 8044
rect 13078 8004 13084 8016
rect 12406 7976 13084 8004
rect 12161 7967 12219 7973
rect 13078 7964 13084 7976
rect 13136 7964 13142 8016
rect 7708 7908 8524 7936
rect 8570 7908 9628 7936
rect 7708 7896 7714 7908
rect 4985 7871 5043 7877
rect 4856 7840 4901 7868
rect 4856 7828 4862 7840
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 5442 7868 5448 7880
rect 5403 7840 5448 7868
rect 4985 7831 5043 7837
rect 3108 7772 3464 7800
rect 3108 7760 3114 7772
rect 3786 7760 3792 7812
rect 3844 7800 3850 7812
rect 4709 7803 4767 7809
rect 4709 7800 4721 7803
rect 3844 7772 4721 7800
rect 3844 7760 3850 7772
rect 4709 7769 4721 7772
rect 4755 7769 4767 7803
rect 5000 7800 5028 7831
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 5626 7868 5632 7880
rect 5587 7840 5632 7868
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 6086 7868 6092 7880
rect 6047 7840 6092 7868
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6236 7840 6469 7868
rect 6236 7828 6242 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7466 7868 7472 7880
rect 6963 7840 7472 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 8496 7877 8524 7908
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7760 7840 8125 7868
rect 5350 7800 5356 7812
rect 5000 7772 5356 7800
rect 4709 7763 4767 7769
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5721 7803 5779 7809
rect 5721 7769 5733 7803
rect 5767 7800 5779 7803
rect 5810 7800 5816 7812
rect 5767 7772 5816 7800
rect 5767 7769 5779 7772
rect 5721 7763 5779 7769
rect 5810 7760 5816 7772
rect 5868 7760 5874 7812
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 7760 7809 7788 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9306 7868 9312 7880
rect 9263 7840 9312 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 7745 7803 7803 7809
rect 7745 7800 7757 7803
rect 6880 7772 7757 7800
rect 6880 7760 6886 7772
rect 7745 7769 7757 7772
rect 7791 7769 7803 7803
rect 7926 7800 7932 7812
rect 7887 7772 7932 7800
rect 7745 7763 7803 7769
rect 7926 7760 7932 7772
rect 7984 7800 7990 7812
rect 8404 7800 8432 7831
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9600 7877 9628 7908
rect 10042 7896 10048 7948
rect 10100 7936 10106 7948
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10100 7908 10241 7936
rect 10100 7896 10106 7908
rect 10229 7905 10241 7908
rect 10275 7905 10287 7939
rect 10962 7936 10968 7948
rect 10229 7899 10287 7905
rect 10428 7908 10968 7936
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9508 7800 9536 7831
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9732 7840 9781 7868
rect 9732 7828 9738 7840
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 10428 7877 10456 7908
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11388 7908 11897 7936
rect 11388 7896 11394 7908
rect 11885 7905 11897 7908
rect 11931 7936 11943 7939
rect 11931 7908 12434 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 10413 7871 10471 7877
rect 9916 7840 9961 7868
rect 9916 7828 9922 7840
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10778 7868 10784 7880
rect 10739 7840 10784 7868
rect 10413 7831 10471 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10873 7871 10931 7877
rect 10873 7837 10885 7871
rect 10919 7868 10931 7871
rect 11054 7868 11060 7880
rect 10919 7840 11060 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 11054 7828 11060 7840
rect 11112 7868 11118 7880
rect 11514 7868 11520 7880
rect 11112 7840 11520 7868
rect 11112 7828 11118 7840
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 11698 7868 11704 7880
rect 11659 7840 11704 7868
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 7984 7772 9536 7800
rect 7984 7760 7990 7772
rect 10594 7760 10600 7812
rect 10652 7800 10658 7812
rect 11333 7803 11391 7809
rect 11333 7800 11345 7803
rect 10652 7772 11345 7800
rect 10652 7760 10658 7772
rect 11333 7769 11345 7772
rect 11379 7769 11391 7803
rect 11333 7763 11391 7769
rect 11882 7760 11888 7812
rect 11940 7800 11946 7812
rect 11977 7803 12035 7809
rect 11977 7800 11989 7803
rect 11940 7772 11989 7800
rect 11940 7760 11946 7772
rect 11977 7769 11989 7772
rect 12023 7769 12035 7803
rect 11977 7763 12035 7769
rect 12066 7760 12072 7812
rect 12124 7800 12130 7812
rect 12124 7772 12169 7800
rect 12124 7760 12130 7772
rect 2590 7732 2596 7744
rect 2004 7704 2452 7732
rect 2551 7704 2596 7732
rect 2004 7692 2010 7704
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 4062 7732 4068 7744
rect 4023 7704 4068 7732
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7732 5227 7735
rect 5534 7732 5540 7744
rect 5215 7704 5540 7732
rect 5215 7701 5227 7704
rect 5169 7695 5227 7701
rect 5534 7692 5540 7704
rect 5592 7692 5598 7744
rect 5902 7732 5908 7744
rect 5863 7704 5908 7732
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 7282 7732 7288 7744
rect 7243 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 8110 7732 8116 7744
rect 7524 7704 8116 7732
rect 7524 7692 7530 7704
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8665 7735 8723 7741
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 8754 7732 8760 7744
rect 8711 7704 8760 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 8754 7692 8760 7704
rect 8812 7732 8818 7744
rect 9122 7732 9128 7744
rect 8812 7704 9128 7732
rect 8812 7692 8818 7704
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 10045 7735 10103 7741
rect 10045 7701 10057 7735
rect 10091 7732 10103 7735
rect 10226 7732 10232 7744
rect 10091 7704 10232 7732
rect 10091 7701 10103 7704
rect 10045 7695 10103 7701
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 10410 7732 10416 7744
rect 10371 7704 10416 7732
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 11241 7735 11299 7741
rect 11241 7732 11253 7735
rect 11204 7704 11253 7732
rect 11204 7692 11210 7704
rect 11241 7701 11253 7704
rect 11287 7701 11299 7735
rect 12406 7732 12434 7908
rect 12710 7868 12716 7880
rect 12671 7840 12716 7868
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 12986 7868 12992 7880
rect 12947 7840 12992 7868
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 12618 7732 12624 7744
rect 12406 7704 12624 7732
rect 11241 7695 11299 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 13449 7735 13507 7741
rect 13449 7732 13461 7735
rect 13412 7704 13461 7732
rect 13412 7692 13418 7704
rect 13449 7701 13461 7704
rect 13495 7701 13507 7735
rect 13449 7695 13507 7701
rect 1104 7642 13892 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 13892 7642
rect 1104 7568 13892 7590
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 1765 7531 1823 7537
rect 1765 7528 1777 7531
rect 1544 7500 1777 7528
rect 1544 7488 1550 7500
rect 1765 7497 1777 7500
rect 1811 7528 1823 7531
rect 2130 7528 2136 7540
rect 1811 7500 2136 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2498 7528 2504 7540
rect 2459 7500 2504 7528
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 3878 7528 3884 7540
rect 3344 7500 3884 7528
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 3344 7460 3372 7500
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7340 7500 7972 7528
rect 7340 7488 7346 7500
rect 1719 7432 3372 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 6914 7420 6920 7472
rect 6972 7420 6978 7472
rect 7944 7469 7972 7500
rect 8110 7488 8116 7540
rect 8168 7488 8174 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8260 7500 8861 7528
rect 8260 7488 8266 7500
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 9214 7528 9220 7540
rect 9175 7500 9220 7528
rect 8849 7491 8907 7497
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 10410 7528 10416 7540
rect 9784 7500 10416 7528
rect 7929 7463 7987 7469
rect 7929 7429 7941 7463
rect 7975 7429 7987 7463
rect 8128 7460 8156 7488
rect 9309 7463 9367 7469
rect 9309 7460 9321 7463
rect 8128 7432 9321 7460
rect 7929 7423 7987 7429
rect 9309 7429 9321 7432
rect 9355 7429 9367 7463
rect 9309 7423 9367 7429
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4264 7364 4629 7392
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 2961 7327 3019 7333
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 3510 7324 3516 7336
rect 3007 7296 3516 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 2222 7188 2228 7200
rect 2183 7160 2228 7188
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 2700 7188 2728 7287
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 3970 7284 3976 7336
rect 4028 7324 4034 7336
rect 4264 7324 4292 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 5350 7392 5356 7404
rect 4939 7364 5356 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5902 7392 5908 7404
rect 5863 7364 5908 7392
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 8754 7401 8760 7404
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 8737 7395 8760 7401
rect 8737 7361 8749 7395
rect 8737 7355 8760 7361
rect 4028 7296 4292 7324
rect 5169 7327 5227 7333
rect 4028 7284 4034 7296
rect 5169 7293 5181 7327
rect 5215 7324 5227 7327
rect 5258 7324 5264 7336
rect 5215 7296 5264 7324
rect 5215 7293 5227 7296
rect 5169 7287 5227 7293
rect 5258 7284 5264 7296
rect 5316 7324 5322 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 5316 7296 8217 7324
rect 5316 7284 5322 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8496 7324 8524 7355
rect 8754 7352 8760 7355
rect 8812 7352 8818 7404
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 9122 7392 9128 7404
rect 8987 7364 9128 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 9784 7401 9812 7500
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 10560 7500 10824 7528
rect 10560 7488 10566 7500
rect 10226 7420 10232 7472
rect 10284 7460 10290 7472
rect 10284 7432 10548 7460
rect 10284 7420 10290 7432
rect 9551 7395 9609 7401
rect 9551 7392 9563 7395
rect 9456 7364 9563 7392
rect 9456 7352 9462 7364
rect 9551 7361 9563 7364
rect 9597 7361 9609 7395
rect 9551 7355 9609 7361
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7392 10011 7395
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9999 7364 10057 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 10045 7361 10057 7364
rect 10091 7392 10103 7395
rect 10134 7392 10140 7404
rect 10091 7364 10140 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 8352 7296 8524 7324
rect 9033 7327 9091 7333
rect 8352 7284 8358 7296
rect 9033 7293 9045 7327
rect 9079 7324 9091 7327
rect 9692 7324 9720 7355
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 10520 7401 10548 7432
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 9858 7324 9864 7336
rect 9079 7296 9864 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 10336 7324 10364 7355
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10652 7364 10697 7392
rect 10652 7352 10658 7364
rect 10796 7324 10824 7500
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 12253 7531 12311 7537
rect 12253 7528 12265 7531
rect 11756 7500 12265 7528
rect 11756 7488 11762 7500
rect 12253 7497 12265 7500
rect 12299 7497 12311 7531
rect 12253 7491 12311 7497
rect 10965 7463 11023 7469
rect 10965 7429 10977 7463
rect 11011 7460 11023 7463
rect 11011 7432 11836 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7361 11207 7395
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 11149 7355 11207 7361
rect 10336 7296 10824 7324
rect 11164 7324 11192 7355
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11808 7401 11836 7432
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 12158 7392 12164 7404
rect 11940 7364 11985 7392
rect 12119 7364 12164 7392
rect 11940 7352 11946 7364
rect 12158 7352 12164 7364
rect 12216 7392 12222 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12216 7364 12909 7392
rect 12216 7352 12222 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 11698 7324 11704 7336
rect 11164 7296 11704 7324
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 12066 7324 12072 7336
rect 12027 7296 12072 7324
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 12526 7284 12532 7336
rect 12584 7324 12590 7336
rect 12986 7324 12992 7336
rect 12584 7296 12992 7324
rect 12584 7284 12590 7296
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 4798 7216 4804 7268
rect 4856 7256 4862 7268
rect 4893 7259 4951 7265
rect 4893 7256 4905 7259
rect 4856 7228 4905 7256
rect 4856 7216 4862 7228
rect 4893 7225 4905 7228
rect 4939 7225 4951 7259
rect 4893 7219 4951 7225
rect 6457 7259 6515 7265
rect 6457 7225 6469 7259
rect 6503 7256 6515 7259
rect 6822 7256 6828 7268
rect 6503 7228 6828 7256
rect 6503 7225 6515 7228
rect 6457 7219 6515 7225
rect 6822 7216 6828 7228
rect 6880 7216 6886 7268
rect 10410 7256 10416 7268
rect 10468 7265 10474 7268
rect 10375 7228 10416 7256
rect 10410 7216 10416 7228
rect 10468 7219 10475 7265
rect 12802 7256 12808 7268
rect 10520 7228 12808 7256
rect 10468 7216 10474 7219
rect 2958 7188 2964 7200
rect 2700 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4614 7188 4620 7200
rect 4479 7160 4620 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 10520 7188 10548 7228
rect 12802 7216 12808 7228
rect 12860 7256 12866 7268
rect 13170 7256 13176 7268
rect 12860 7228 13176 7256
rect 12860 7216 12866 7228
rect 13170 7216 13176 7228
rect 13228 7216 13234 7268
rect 11606 7188 11612 7200
rect 8343 7160 10548 7188
rect 11567 7160 11612 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 13538 7188 13544 7200
rect 13499 7160 13544 7188
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 1104 7098 13892 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 13892 7098
rect 1104 7024 13892 7046
rect 1486 6984 1492 6996
rect 1447 6956 1492 6984
rect 1486 6944 1492 6956
rect 1544 6944 1550 6996
rect 3510 6984 3516 6996
rect 3471 6956 3516 6984
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6822 6984 6828 6996
rect 5592 6956 6828 6984
rect 5592 6944 5598 6956
rect 6822 6944 6828 6956
rect 6880 6984 6886 6996
rect 6880 6956 7788 6984
rect 6880 6944 6886 6956
rect 7760 6916 7788 6956
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10410 6984 10416 6996
rect 10008 6956 10416 6984
rect 10008 6944 10014 6956
rect 10410 6944 10416 6956
rect 10468 6984 10474 6996
rect 10962 6984 10968 6996
rect 10468 6956 10968 6984
rect 10468 6944 10474 6956
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11606 6944 11612 6996
rect 11664 6984 11670 6996
rect 12081 6987 12139 6993
rect 12081 6984 12093 6987
rect 11664 6956 12093 6984
rect 11664 6944 11670 6956
rect 12081 6953 12093 6956
rect 12127 6953 12139 6987
rect 12618 6984 12624 6996
rect 12579 6956 12624 6984
rect 12081 6947 12139 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 11054 6916 11060 6928
rect 7760 6888 11060 6916
rect 11054 6876 11060 6888
rect 11112 6876 11118 6928
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3237 6851 3295 6857
rect 3237 6848 3249 6851
rect 3016 6820 3249 6848
rect 3016 6808 3022 6820
rect 3237 6817 3249 6820
rect 3283 6848 3295 6851
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3283 6820 3985 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3973 6817 3985 6820
rect 4019 6848 4031 6851
rect 5258 6848 5264 6860
rect 4019 6820 5264 6848
rect 4019 6817 4031 6820
rect 3973 6811 4031 6817
rect 5258 6808 5264 6820
rect 5316 6848 5322 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 5316 6820 6469 6848
rect 5316 6808 5322 6820
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 7926 6808 7932 6860
rect 7984 6848 7990 6860
rect 7984 6820 8156 6848
rect 7984 6808 7990 6820
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6780 3387 6783
rect 3418 6780 3424 6792
rect 3375 6752 3424 6780
rect 3375 6749 3387 6752
rect 3329 6743 3387 6749
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 3786 6780 3792 6792
rect 3747 6752 3792 6780
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6749 6239 6783
rect 6362 6780 6368 6792
rect 6323 6752 6368 6780
rect 6181 6743 6239 6749
rect 2682 6712 2688 6724
rect 2530 6684 2688 6712
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 2958 6712 2964 6724
rect 2919 6684 2964 6712
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 4246 6712 4252 6724
rect 4207 6684 4252 6712
rect 4246 6672 4252 6684
rect 4304 6672 4310 6724
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 5474 6684 6009 6712
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 5721 6647 5779 6653
rect 5721 6644 5733 6647
rect 5684 6616 5733 6644
rect 5684 6604 5690 6616
rect 5721 6613 5733 6616
rect 5767 6613 5779 6647
rect 6196 6644 6224 6743
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6733 6715 6791 6721
rect 6733 6681 6745 6715
rect 6779 6712 6791 6715
rect 7006 6712 7012 6724
rect 6779 6684 7012 6712
rect 6779 6681 6791 6684
rect 6733 6675 6791 6681
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7282 6672 7288 6724
rect 7340 6672 7346 6724
rect 8128 6656 8156 6820
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10376 6820 10609 6848
rect 10376 6808 10382 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12345 6851 12403 6857
rect 12345 6848 12357 6851
rect 12124 6820 12357 6848
rect 12124 6808 12130 6820
rect 12345 6817 12357 6820
rect 12391 6817 12403 6851
rect 12986 6848 12992 6860
rect 12345 6811 12403 6817
rect 12636 6820 12992 6848
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 9180 6752 9229 6780
rect 9180 6740 9186 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 9858 6780 9864 6792
rect 9723 6752 9864 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 12636 6789 12664 6820
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 13170 6848 13176 6860
rect 13131 6820 13176 6848
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 12851 6783 12909 6789
rect 12851 6780 12863 6783
rect 12768 6752 12863 6780
rect 12768 6740 12774 6752
rect 12851 6749 12863 6752
rect 12897 6749 12909 6783
rect 13446 6780 13452 6792
rect 13407 6752 13452 6780
rect 12851 6743 12909 6749
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 8294 6672 8300 6724
rect 8352 6712 8358 6724
rect 10410 6712 10416 6724
rect 8352 6684 10416 6712
rect 8352 6672 8358 6684
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 11054 6672 11060 6724
rect 11112 6672 11118 6724
rect 13354 6712 13360 6724
rect 13004 6684 13360 6712
rect 7098 6644 7104 6656
rect 6196 6616 7104 6644
rect 5721 6607 5779 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 8168 6616 8217 6644
rect 8168 6604 8174 6616
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 10045 6647 10103 6653
rect 10045 6644 10057 6647
rect 9364 6616 10057 6644
rect 9364 6604 9370 6616
rect 10045 6613 10057 6616
rect 10091 6613 10103 6647
rect 10318 6644 10324 6656
rect 10231 6616 10324 6644
rect 10045 6607 10103 6613
rect 10318 6604 10324 6616
rect 10376 6644 10382 6656
rect 11790 6644 11796 6656
rect 10376 6616 11796 6644
rect 10376 6604 10382 6616
rect 11790 6604 11796 6616
rect 11848 6644 11854 6656
rect 12158 6644 12164 6656
rect 11848 6616 12164 6644
rect 11848 6604 11854 6616
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 13004 6653 13032 6684
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 12989 6647 13047 6653
rect 12989 6613 13001 6647
rect 13035 6613 13047 6647
rect 12989 6607 13047 6613
rect 13078 6604 13084 6656
rect 13136 6644 13142 6656
rect 13262 6644 13268 6656
rect 13136 6616 13181 6644
rect 13223 6616 13268 6644
rect 13136 6604 13142 6616
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 1104 6554 13892 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 13892 6554
rect 1104 6480 13892 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 2685 6443 2743 6449
rect 1820 6412 1992 6440
rect 1820 6400 1826 6412
rect 1486 6332 1492 6384
rect 1544 6372 1550 6384
rect 1857 6375 1915 6381
rect 1857 6372 1869 6375
rect 1544 6344 1869 6372
rect 1544 6332 1550 6344
rect 1857 6341 1869 6344
rect 1903 6341 1915 6375
rect 1964 6372 1992 6412
rect 2685 6409 2697 6443
rect 2731 6440 2743 6443
rect 2958 6440 2964 6452
rect 2731 6412 2964 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 4304 6412 4445 6440
rect 4304 6400 4310 6412
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 4433 6403 4491 6409
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6972 6412 7021 6440
rect 6972 6400 6978 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 7282 6440 7288 6452
rect 7243 6412 7288 6440
rect 7009 6403 7067 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 8757 6443 8815 6449
rect 8757 6409 8769 6443
rect 8803 6440 8815 6443
rect 9122 6440 9128 6452
rect 8803 6412 9128 6440
rect 8803 6409 8815 6412
rect 8757 6403 8815 6409
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 9306 6440 9312 6452
rect 9267 6412 9312 6440
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 10318 6440 10324 6452
rect 9600 6412 10324 6440
rect 3881 6375 3939 6381
rect 1964 6344 3832 6372
rect 1857 6335 1915 6341
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 1762 6304 1768 6316
rect 1719 6276 1768 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1872 6276 2145 6304
rect 1489 6239 1547 6245
rect 1489 6205 1501 6239
rect 1535 6236 1547 6239
rect 1872 6236 1900 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2222 6264 2228 6316
rect 2280 6304 2286 6316
rect 2501 6307 2559 6313
rect 2501 6304 2513 6307
rect 2280 6276 2513 6304
rect 2280 6264 2286 6276
rect 2501 6273 2513 6276
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2924 6276 2973 6304
rect 2924 6264 2930 6276
rect 2961 6273 2973 6276
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 3694 6304 3700 6316
rect 3283 6276 3700 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 3804 6304 3832 6344
rect 3881 6341 3893 6375
rect 3927 6372 3939 6375
rect 4614 6372 4620 6384
rect 3927 6344 4620 6372
rect 3927 6341 3939 6344
rect 3881 6335 3939 6341
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 7116 6344 7420 6372
rect 7116 6316 7144 6344
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 3804 6276 4905 6304
rect 1535 6208 1900 6236
rect 1949 6239 2007 6245
rect 1535 6205 1547 6208
rect 1489 6199 1547 6205
rect 1949 6205 1961 6239
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6205 3939 6239
rect 3881 6199 3939 6205
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 1964 6168 1992 6199
rect 1912 6140 1992 6168
rect 1912 6128 1918 6140
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 3145 6171 3203 6177
rect 3145 6168 3157 6171
rect 3108 6140 3157 6168
rect 3108 6128 3114 6140
rect 3145 6137 3157 6140
rect 3191 6137 3203 6171
rect 3418 6168 3424 6180
rect 3379 6140 3424 6168
rect 3145 6131 3203 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 3896 6168 3924 6199
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 4617 6239 4675 6245
rect 4617 6236 4629 6239
rect 4028 6208 4629 6236
rect 4028 6196 4034 6208
rect 4617 6205 4629 6208
rect 4663 6205 4675 6239
rect 4617 6199 4675 6205
rect 4062 6168 4068 6180
rect 3896 6140 4068 6168
rect 4062 6128 4068 6140
rect 4120 6128 4126 6180
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 1544 6072 2329 6100
rect 1544 6060 1550 6072
rect 2317 6069 2329 6072
rect 2363 6069 2375 6103
rect 2317 6063 2375 6069
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 3752 6072 4169 6100
rect 3752 6060 3758 6072
rect 4157 6069 4169 6072
rect 4203 6069 4215 6103
rect 4632 6100 4660 6199
rect 4724 6168 4752 6276
rect 4893 6273 4905 6276
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5500 6276 5549 6304
rect 5500 6264 5506 6276
rect 5537 6273 5549 6276
rect 5583 6304 5595 6307
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5583 6276 5733 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5721 6273 5733 6276
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6178 6304 6184 6316
rect 5951 6276 6184 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6420 6276 6745 6304
rect 6420 6264 6426 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7098 6304 7104 6316
rect 7055 6276 7104 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6236 4859 6239
rect 5460 6236 5488 6264
rect 6086 6236 6092 6248
rect 4847 6208 5488 6236
rect 6047 6208 6092 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 6086 6196 6092 6208
rect 6144 6196 6150 6248
rect 6748 6236 6776 6267
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7392 6313 7420 6344
rect 7193 6307 7251 6313
rect 7193 6273 7205 6307
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7208 6236 7236 6267
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7800 6276 7941 6304
rect 7800 6264 7806 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 9307 6307 9365 6313
rect 9307 6304 9319 6307
rect 9180 6276 9319 6304
rect 9180 6264 9186 6276
rect 9307 6273 9319 6276
rect 9353 6304 9365 6307
rect 9600 6304 9628 6412
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10836 6412 10885 6440
rect 10836 6400 10842 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 11241 6443 11299 6449
rect 11241 6409 11253 6443
rect 11287 6440 11299 6443
rect 11882 6440 11888 6452
rect 11287 6412 11888 6440
rect 11287 6409 11299 6412
rect 11241 6403 11299 6409
rect 9858 6372 9864 6384
rect 9819 6344 9864 6372
rect 9858 6332 9864 6344
rect 9916 6332 9922 6384
rect 10410 6332 10416 6384
rect 10468 6372 10474 6384
rect 10962 6372 10968 6384
rect 10468 6344 10824 6372
rect 10875 6344 10968 6372
rect 10468 6332 10474 6344
rect 9353 6276 9628 6304
rect 9353 6273 9365 6276
rect 9307 6267 9365 6273
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 10134 6313 10140 6316
rect 10103 6307 10140 6313
rect 10103 6304 10115 6307
rect 9732 6276 10115 6304
rect 9732 6264 9738 6276
rect 10103 6273 10115 6276
rect 10103 6267 10140 6273
rect 10134 6264 10140 6267
rect 10192 6264 10198 6316
rect 10597 6307 10655 6313
rect 10597 6304 10609 6307
rect 10244 6276 10609 6304
rect 6748 6208 7236 6236
rect 6932 6180 6960 6208
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 7340 6208 7849 6236
rect 7340 6196 7346 6208
rect 7837 6205 7849 6208
rect 7883 6236 7895 6239
rect 8018 6236 8024 6248
rect 7883 6208 8024 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 8168 6208 9781 6236
rect 8168 6196 8174 6208
rect 9769 6205 9781 6208
rect 9815 6236 9827 6239
rect 10244 6236 10272 6276
rect 10597 6273 10609 6276
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 10410 6236 10416 6248
rect 9815 6208 10272 6236
rect 10371 6208 10416 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 10796 6236 10824 6344
rect 10888 6313 10916 6344
rect 10962 6332 10968 6344
rect 11020 6372 11026 6384
rect 11256 6372 11284 6403
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12161 6443 12219 6449
rect 12161 6409 12173 6443
rect 12207 6440 12219 6443
rect 12894 6440 12900 6452
rect 12207 6412 12900 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 12894 6400 12900 6412
rect 12952 6400 12958 6452
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 13722 6440 13728 6452
rect 13495 6412 13728 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 11020 6344 11284 6372
rect 11020 6332 11026 6344
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 12069 6375 12127 6381
rect 11480 6344 11836 6372
rect 11480 6332 11486 6344
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6273 11115 6307
rect 11514 6304 11520 6316
rect 11475 6276 11520 6304
rect 11057 6267 11115 6273
rect 11072 6236 11100 6267
rect 11514 6264 11520 6276
rect 11572 6264 11578 6316
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11808 6304 11836 6344
rect 12069 6341 12081 6375
rect 12115 6372 12127 6375
rect 13630 6372 13636 6384
rect 12115 6344 13636 6372
rect 12115 6341 12127 6344
rect 12069 6335 12127 6341
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 11882 6304 11888 6316
rect 11808 6276 11888 6304
rect 11882 6264 11888 6276
rect 11940 6304 11946 6316
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 11940 6276 12265 6304
rect 11940 6264 11946 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 12434 6304 12440 6316
rect 12395 6276 12440 6304
rect 12253 6267 12311 6273
rect 10560 6208 10605 6236
rect 10796 6208 11100 6236
rect 12268 6236 12296 6267
rect 12434 6264 12440 6276
rect 12492 6304 12498 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12492 6276 12909 6304
rect 12492 6264 12498 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13096 6236 13124 6267
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13265 6307 13323 6313
rect 13265 6304 13277 6307
rect 13228 6276 13277 6304
rect 13228 6264 13234 6276
rect 13265 6273 13277 6276
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 12268 6208 13124 6236
rect 10560 6196 10566 6208
rect 5626 6168 5632 6180
rect 4724 6140 5632 6168
rect 4706 6100 4712 6112
rect 4632 6072 4712 6100
rect 4157 6063 4215 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5276 6109 5304 6140
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 6914 6128 6920 6180
rect 6972 6128 6978 6180
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 9125 6171 9183 6177
rect 9125 6168 9137 6171
rect 7064 6140 9137 6168
rect 7064 6128 7070 6140
rect 9125 6137 9137 6140
rect 9171 6137 9183 6171
rect 9125 6131 9183 6137
rect 9677 6171 9735 6177
rect 9677 6137 9689 6171
rect 9723 6168 9735 6171
rect 9858 6168 9864 6180
rect 9723 6140 9864 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 9858 6128 9864 6140
rect 9916 6168 9922 6180
rect 10594 6168 10600 6180
rect 9916 6140 10600 6168
rect 9916 6128 9922 6140
rect 10594 6128 10600 6140
rect 10652 6128 10658 6180
rect 12894 6168 12900 6180
rect 12855 6140 12900 6168
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 5077 6103 5135 6109
rect 5077 6100 5089 6103
rect 4948 6072 5089 6100
rect 4948 6060 4954 6072
rect 5077 6069 5089 6072
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 5261 6103 5319 6109
rect 5261 6069 5273 6103
rect 5307 6069 5319 6103
rect 5261 6063 5319 6069
rect 5350 6060 5356 6112
rect 5408 6100 5414 6112
rect 7190 6100 7196 6112
rect 5408 6072 7196 6100
rect 5408 6060 5414 6072
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10042 6100 10048 6112
rect 9824 6072 10048 6100
rect 9824 6060 9830 6072
rect 10042 6060 10048 6072
rect 10100 6100 10106 6112
rect 10502 6100 10508 6112
rect 10100 6072 10508 6100
rect 10100 6060 10106 6072
rect 10502 6060 10508 6072
rect 10560 6100 10566 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 10560 6072 11805 6100
rect 10560 6060 10566 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 12618 6100 12624 6112
rect 12579 6072 12624 6100
rect 11793 6063 11851 6069
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 1104 6010 13892 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 13892 6010
rect 1104 5936 13892 5958
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3329 5899 3387 5905
rect 3329 5896 3341 5899
rect 2924 5868 3341 5896
rect 2924 5856 2930 5868
rect 3329 5865 3341 5868
rect 3375 5865 3387 5899
rect 3329 5859 3387 5865
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4982 5896 4988 5908
rect 4212 5868 4988 5896
rect 4212 5856 4218 5868
rect 1578 5788 1584 5840
rect 1636 5828 1642 5840
rect 2314 5828 2320 5840
rect 1636 5800 2320 5828
rect 1636 5788 1642 5800
rect 2314 5788 2320 5800
rect 2372 5828 2378 5840
rect 2372 5800 3004 5828
rect 2372 5788 2378 5800
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 2777 5763 2835 5769
rect 2777 5760 2789 5763
rect 1811 5732 2789 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 2777 5729 2789 5732
rect 2823 5729 2835 5763
rect 2777 5723 2835 5729
rect 1486 5692 1492 5704
rect 1447 5664 1492 5692
rect 1486 5652 1492 5664
rect 1544 5652 1550 5704
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 1596 5556 1624 5655
rect 1854 5652 1860 5704
rect 1912 5692 1918 5704
rect 1949 5695 2007 5701
rect 1949 5692 1961 5695
rect 1912 5664 1961 5692
rect 1912 5652 1918 5664
rect 1949 5661 1961 5664
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 1670 5584 1676 5636
rect 1728 5624 1734 5636
rect 2148 5624 2176 5655
rect 1728 5596 2176 5624
rect 2240 5624 2268 5655
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 2682 5692 2688 5704
rect 2372 5664 2417 5692
rect 2516 5664 2688 5692
rect 2372 5652 2378 5664
rect 2516 5624 2544 5664
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2976 5701 3004 5800
rect 4264 5769 4292 5868
rect 4982 5856 4988 5868
rect 5040 5896 5046 5908
rect 6086 5896 6092 5908
rect 5040 5868 6092 5896
rect 5040 5856 5046 5868
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5729 4307 5763
rect 4614 5760 4620 5772
rect 4249 5723 4307 5729
rect 4356 5732 4620 5760
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3513 5695 3571 5701
rect 3513 5692 3525 5695
rect 3007 5664 3525 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3513 5661 3525 5664
rect 3559 5661 3571 5695
rect 3513 5655 3571 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4356 5692 4384 5732
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 5092 5711 5120 5868
rect 6086 5856 6092 5868
rect 6144 5896 6150 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6144 5868 7205 5896
rect 6144 5856 6150 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 9674 5896 9680 5908
rect 7193 5859 7251 5865
rect 8588 5868 9680 5896
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 6972 5732 7788 5760
rect 6972 5720 6978 5732
rect 5078 5705 5136 5711
rect 4111 5664 4384 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 4706 5692 4712 5704
rect 4580 5664 4625 5692
rect 4667 5664 4712 5692
rect 4580 5652 4586 5664
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 4890 5692 4896 5704
rect 4851 5664 4896 5692
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 5078 5671 5090 5705
rect 5124 5671 5136 5705
rect 5442 5692 5448 5704
rect 5078 5665 5136 5671
rect 5403 5664 5448 5692
rect 4985 5655 5043 5661
rect 2240 5596 2544 5624
rect 2593 5627 2651 5633
rect 1728 5584 1734 5596
rect 2593 5593 2605 5627
rect 2639 5624 2651 5627
rect 2866 5624 2872 5636
rect 2639 5596 2872 5624
rect 2639 5593 2651 5596
rect 2593 5587 2651 5593
rect 2866 5584 2872 5596
rect 2924 5584 2930 5636
rect 5000 5624 5028 5655
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 7190 5652 7196 5704
rect 7248 5692 7254 5704
rect 7760 5701 7788 5732
rect 8588 5701 8616 5868
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 10762 5899 10820 5905
rect 10762 5896 10774 5899
rect 10060 5868 10774 5896
rect 8665 5831 8723 5837
rect 8665 5797 8677 5831
rect 8711 5797 8723 5831
rect 8665 5791 8723 5797
rect 9033 5831 9091 5837
rect 9033 5797 9045 5831
rect 9079 5828 9091 5831
rect 10060 5828 10088 5868
rect 10762 5865 10774 5868
rect 10808 5865 10820 5899
rect 10762 5859 10820 5865
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 12710 5896 12716 5908
rect 12584 5868 12716 5896
rect 12584 5856 12590 5868
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 9079 5800 10088 5828
rect 9079 5797 9091 5800
rect 9033 5791 9091 5797
rect 8680 5760 8708 5791
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 8680 5732 9505 5760
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 10318 5760 10324 5772
rect 9493 5723 9551 5729
rect 9600 5732 10324 5760
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 7248 5664 7389 5692
rect 7248 5652 7254 5664
rect 7377 5661 7389 5664
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 8573 5655 8631 5661
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 8846 5692 8852 5704
rect 8803 5664 8852 5692
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 5353 5627 5411 5633
rect 5000 5596 5120 5624
rect 1946 5556 1952 5568
rect 1596 5528 1952 5556
rect 1946 5516 1952 5528
rect 2004 5556 2010 5568
rect 2222 5556 2228 5568
rect 2004 5528 2228 5556
rect 2004 5516 2010 5528
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 3145 5559 3203 5565
rect 3145 5556 3157 5559
rect 3108 5528 3157 5556
rect 3108 5516 3114 5528
rect 3145 5525 3157 5528
rect 3191 5525 3203 5559
rect 3878 5556 3884 5568
rect 3839 5528 3884 5556
rect 3145 5519 3203 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 4433 5559 4491 5565
rect 4433 5556 4445 5559
rect 4212 5528 4445 5556
rect 4212 5516 4218 5528
rect 4433 5525 4445 5528
rect 4479 5525 4491 5559
rect 5092 5556 5120 5596
rect 5353 5593 5365 5627
rect 5399 5624 5411 5627
rect 5721 5627 5779 5633
rect 5721 5624 5733 5627
rect 5399 5596 5733 5624
rect 5399 5593 5411 5596
rect 5353 5587 5411 5593
rect 5721 5593 5733 5596
rect 5767 5593 5779 5627
rect 5721 5587 5779 5593
rect 6454 5584 6460 5636
rect 6512 5584 6518 5636
rect 7098 5584 7104 5636
rect 7156 5624 7162 5636
rect 7944 5624 7972 5655
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9600 5692 9628 5732
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 12066 5760 12072 5772
rect 10520 5732 12072 5760
rect 9263 5664 9628 5692
rect 9769 5695 9827 5701
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9769 5661 9781 5695
rect 9815 5692 9827 5695
rect 9950 5692 9956 5704
rect 9815 5664 9956 5692
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10042 5652 10048 5704
rect 10100 5692 10106 5704
rect 10520 5701 10548 5732
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 12986 5720 12992 5772
rect 13044 5760 13050 5772
rect 13265 5763 13323 5769
rect 13265 5760 13277 5763
rect 13044 5732 13277 5760
rect 13044 5720 13050 5732
rect 13265 5729 13277 5732
rect 13311 5729 13323 5763
rect 13265 5723 13323 5729
rect 12808 5704 12860 5710
rect 10505 5695 10563 5701
rect 10505 5692 10517 5695
rect 10100 5664 10517 5692
rect 10100 5652 10106 5664
rect 10505 5661 10517 5664
rect 10551 5661 10563 5695
rect 10505 5655 10563 5661
rect 12808 5646 12860 5652
rect 7156 5596 7972 5624
rect 8113 5627 8171 5633
rect 7156 5584 7162 5596
rect 8113 5593 8125 5627
rect 8159 5624 8171 5627
rect 8159 5596 11270 5624
rect 8159 5593 8171 5596
rect 8113 5587 8171 5593
rect 12066 5584 12072 5636
rect 12124 5624 12130 5636
rect 12437 5627 12495 5633
rect 12437 5624 12449 5627
rect 12124 5596 12449 5624
rect 12124 5584 12130 5596
rect 12437 5593 12449 5596
rect 12483 5593 12495 5627
rect 12437 5587 12495 5593
rect 6086 5556 6092 5568
rect 5092 5528 6092 5556
rect 4433 5519 4491 5525
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 7561 5559 7619 5565
rect 7561 5525 7573 5559
rect 7607 5556 7619 5559
rect 7742 5556 7748 5568
rect 7607 5528 7748 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 8846 5516 8852 5568
rect 8904 5556 8910 5568
rect 10226 5556 10232 5568
rect 8904 5528 10232 5556
rect 8904 5516 8910 5528
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10410 5556 10416 5568
rect 10371 5528 10416 5556
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 12253 5559 12311 5565
rect 12253 5525 12265 5559
rect 12299 5556 12311 5559
rect 12802 5556 12808 5568
rect 12299 5528 12808 5556
rect 12299 5525 12311 5528
rect 12253 5519 12311 5525
rect 12802 5516 12808 5528
rect 12860 5556 12866 5568
rect 13262 5556 13268 5568
rect 12860 5528 13268 5556
rect 12860 5516 12866 5528
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 1104 5466 13892 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 13892 5466
rect 1104 5392 13892 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3602 5352 3608 5364
rect 3191 5324 3608 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5352 3755 5355
rect 4154 5352 4160 5364
rect 3743 5324 4160 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 8110 5352 8116 5364
rect 5500 5324 8116 5352
rect 5500 5312 5506 5324
rect 1581 5287 1639 5293
rect 1581 5253 1593 5287
rect 1627 5284 1639 5287
rect 1949 5287 2007 5293
rect 1627 5256 1900 5284
rect 1627 5253 1639 5256
rect 1581 5247 1639 5253
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5185 1823 5219
rect 1872 5216 1900 5256
rect 1949 5253 1961 5287
rect 1995 5284 2007 5287
rect 3878 5284 3884 5296
rect 1995 5256 3884 5284
rect 1995 5253 2007 5256
rect 1949 5247 2007 5253
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 4798 5244 4804 5296
rect 4856 5244 4862 5296
rect 2406 5216 2412 5228
rect 1872 5188 2268 5216
rect 2367 5188 2412 5216
rect 1765 5179 1823 5185
rect 1780 5012 1808 5179
rect 2038 5148 2044 5160
rect 1999 5120 2044 5148
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 2240 5148 2268 5188
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2516 5188 2973 5216
rect 2516 5148 2544 5188
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5216 3295 5219
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 3283 5188 3525 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 3513 5185 3525 5188
rect 3559 5216 3571 5219
rect 3970 5216 3976 5228
rect 3559 5188 3976 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 2240 5120 2544 5148
rect 2593 5151 2651 5157
rect 2593 5117 2605 5151
rect 2639 5148 2651 5151
rect 2774 5148 2780 5160
rect 2639 5120 2780 5148
rect 2639 5117 2651 5120
rect 2593 5111 2651 5117
rect 2774 5108 2780 5120
rect 2832 5148 2838 5160
rect 2976 5148 3004 5179
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 5828 5225 5856 5324
rect 8110 5312 8116 5324
rect 8168 5352 8174 5364
rect 9858 5352 9864 5364
rect 8168 5324 9168 5352
rect 9819 5324 9864 5352
rect 8168 5312 8174 5324
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 6512 5256 6561 5284
rect 6512 5244 6518 5256
rect 6549 5253 6561 5256
rect 6595 5253 6607 5287
rect 7098 5284 7104 5296
rect 6549 5247 6607 5253
rect 6748 5256 7104 5284
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5902 5176 5908 5228
rect 5960 5216 5966 5228
rect 6748 5225 6776 5256
rect 7098 5244 7104 5256
rect 7156 5244 7162 5296
rect 7834 5244 7840 5296
rect 7892 5244 7898 5296
rect 6733 5219 6791 5225
rect 5960 5188 6005 5216
rect 5960 5176 5966 5188
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6914 5216 6920 5228
rect 6875 5188 6920 5216
rect 6733 5179 6791 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 9140 5225 9168 5324
rect 9858 5312 9864 5324
rect 9916 5352 9922 5364
rect 9916 5324 10180 5352
rect 9916 5312 9922 5324
rect 9585 5287 9643 5293
rect 9585 5253 9597 5287
rect 9631 5284 9643 5287
rect 9950 5284 9956 5296
rect 9631 5256 9956 5284
rect 9631 5253 9643 5256
rect 9585 5247 9643 5253
rect 9950 5244 9956 5256
rect 10008 5244 10014 5296
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9490 5216 9496 5228
rect 9451 5188 9496 5216
rect 9125 5179 9183 5185
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 9858 5216 9864 5228
rect 9723 5188 9864 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 10152 5216 10180 5324
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 11591 5355 11649 5361
rect 11591 5352 11603 5355
rect 10376 5324 11603 5352
rect 10376 5312 10382 5324
rect 11591 5321 11603 5324
rect 11637 5321 11649 5355
rect 12066 5352 12072 5364
rect 12027 5324 12072 5352
rect 11591 5315 11649 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 12406 5324 13461 5352
rect 10226 5244 10232 5296
rect 10284 5284 10290 5296
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 10284 5256 10701 5284
rect 10284 5244 10290 5256
rect 10689 5253 10701 5256
rect 10735 5253 10747 5287
rect 11238 5284 11244 5296
rect 10689 5247 10747 5253
rect 10888 5256 11244 5284
rect 10888 5225 10916 5256
rect 11238 5244 11244 5256
rect 11296 5284 11302 5296
rect 11698 5284 11704 5296
rect 11296 5256 11704 5284
rect 11296 5244 11302 5256
rect 11698 5244 11704 5256
rect 11756 5244 11762 5296
rect 11790 5244 11796 5296
rect 11848 5284 11854 5296
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 11848 5256 12173 5284
rect 11848 5244 11854 5256
rect 12161 5253 12173 5256
rect 12207 5253 12219 5287
rect 12161 5247 12219 5253
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10152 5188 10517 5216
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 11057 5219 11115 5225
rect 11057 5185 11069 5219
rect 11103 5216 11115 5219
rect 11514 5216 11520 5228
rect 11103 5188 11520 5216
rect 11103 5185 11115 5188
rect 11057 5179 11115 5185
rect 3786 5148 3792 5160
rect 2832 5120 2877 5148
rect 2976 5120 3792 5148
rect 2832 5108 2838 5120
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 8849 5151 8907 5157
rect 5583 5120 6132 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 1946 5040 1952 5092
rect 2004 5080 2010 5092
rect 2133 5083 2191 5089
rect 2133 5080 2145 5083
rect 2004 5052 2145 5080
rect 2004 5040 2010 5052
rect 2133 5049 2145 5052
rect 2179 5049 2191 5083
rect 2133 5043 2191 5049
rect 2222 5040 2228 5092
rect 2280 5080 2286 5092
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 2280 5052 3341 5080
rect 2280 5040 2286 5052
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 4522 5080 4528 5092
rect 3329 5043 3387 5049
rect 3988 5052 4528 5080
rect 3878 5012 3884 5024
rect 1780 4984 3884 5012
rect 3878 4972 3884 4984
rect 3936 5012 3942 5024
rect 3988 5012 4016 5052
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 6104 5089 6132 5120
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 8895 5120 10149 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10318 5148 10324 5160
rect 10279 5120 10324 5148
rect 10137 5111 10195 5117
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 10612 5148 10640 5179
rect 11072 5148 11100 5179
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 11882 5216 11888 5228
rect 11795 5188 11888 5216
rect 11882 5176 11888 5188
rect 11940 5216 11946 5228
rect 12406 5216 12434 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 11940 5188 12434 5216
rect 11940 5176 11946 5188
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 12851 5219 12909 5225
rect 12851 5216 12863 5219
rect 12768 5188 12863 5216
rect 12768 5176 12774 5188
rect 12851 5185 12863 5188
rect 12897 5185 12909 5219
rect 12986 5216 12992 5228
rect 12947 5188 12992 5216
rect 12851 5179 12909 5185
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 13262 5216 13268 5228
rect 13223 5188 13268 5216
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 12618 5148 12624 5160
rect 10612 5120 11100 5148
rect 12531 5120 12624 5148
rect 6089 5083 6147 5089
rect 6089 5049 6101 5083
rect 6135 5049 6147 5083
rect 9306 5080 9312 5092
rect 9267 5052 9312 5080
rect 6089 5043 6147 5049
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 10042 5080 10048 5092
rect 9456 5052 10048 5080
rect 9456 5040 9462 5052
rect 10042 5040 10048 5052
rect 10100 5040 10106 5092
rect 3936 4984 4016 5012
rect 4065 5015 4123 5021
rect 3936 4972 3942 4984
rect 4065 4981 4077 5015
rect 4111 5012 4123 5015
rect 4890 5012 4896 5024
rect 4111 4984 4896 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 7377 5015 7435 5021
rect 7377 4981 7389 5015
rect 7423 5012 7435 5015
rect 9214 5012 9220 5024
rect 7423 4984 9220 5012
rect 7423 4981 7435 4984
rect 7377 4975 7435 4981
rect 9214 4972 9220 4984
rect 9272 5012 9278 5024
rect 10612 5012 10640 5120
rect 12618 5108 12624 5120
rect 12676 5148 12682 5160
rect 13078 5148 13084 5160
rect 12676 5120 13084 5148
rect 12676 5108 12682 5120
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 12710 5080 12716 5092
rect 12671 5052 12716 5080
rect 12710 5040 12716 5052
rect 12768 5040 12774 5092
rect 9272 4984 10640 5012
rect 9272 4972 9278 4984
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12618 5012 12624 5024
rect 12584 4984 12624 5012
rect 12584 4972 12590 4984
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 1104 4922 13892 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 13892 4922
rect 1104 4848 13892 4870
rect 1489 4811 1547 4817
rect 1489 4777 1501 4811
rect 1535 4808 1547 4811
rect 3329 4811 3387 4817
rect 1535 4780 3004 4808
rect 1535 4777 1547 4780
rect 1489 4771 1547 4777
rect 2130 4740 2136 4752
rect 1872 4712 2136 4740
rect 1872 4681 1900 4712
rect 2130 4700 2136 4712
rect 2188 4700 2194 4752
rect 2976 4749 3004 4780
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 5371 4811 5429 4817
rect 3375 4780 5316 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 2961 4743 3019 4749
rect 2961 4709 2973 4743
rect 3007 4709 3019 4743
rect 5288 4740 5316 4780
rect 5371 4777 5383 4811
rect 5417 4808 5429 4811
rect 5902 4808 5908 4820
rect 5417 4780 5908 4808
rect 5417 4777 5429 4780
rect 5371 4771 5429 4777
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7561 4811 7619 4817
rect 7561 4808 7573 4811
rect 6972 4780 7573 4808
rect 6972 4768 6978 4780
rect 7561 4777 7573 4780
rect 7607 4777 7619 4811
rect 7561 4771 7619 4777
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 10318 4808 10324 4820
rect 9355 4780 10324 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 7009 4743 7067 4749
rect 5288 4712 6960 4740
rect 2961 4703 3019 4709
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4641 1915 4675
rect 3326 4672 3332 4684
rect 1857 4635 1915 4641
rect 2148 4644 3332 4672
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 2148 4613 2176 4644
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 3602 4632 3608 4684
rect 3660 4672 3666 4684
rect 3660 4644 4476 4672
rect 3660 4632 3666 4644
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4573 2191 4607
rect 2363 4607 2421 4613
rect 2363 4604 2375 4607
rect 2133 4567 2191 4573
rect 2240 4576 2375 4604
rect 1486 4496 1492 4548
rect 1544 4536 1550 4548
rect 2240 4536 2268 4576
rect 2363 4573 2375 4576
rect 2409 4573 2421 4607
rect 2363 4567 2421 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 2774 4604 2780 4616
rect 2731 4576 2780 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 3050 4604 3056 4616
rect 2924 4576 2969 4604
rect 3011 4576 3056 4604
rect 2924 4564 2930 4576
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3786 4604 3792 4616
rect 3200 4576 3245 4604
rect 3747 4576 3792 4604
rect 3200 4564 3206 4576
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4448 4613 4476 4644
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4764 4644 4813 4672
rect 4764 4632 4770 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 4890 4632 4896 4684
rect 4948 4672 4954 4684
rect 6932 4672 6960 4712
rect 7009 4709 7021 4743
rect 7055 4740 7067 4743
rect 7098 4740 7104 4752
rect 7055 4712 7104 4740
rect 7055 4709 7067 4712
rect 7009 4703 7067 4709
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 7282 4672 7288 4684
rect 4948 4644 5948 4672
rect 6932 4644 7288 4672
rect 4948 4632 4954 4644
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 4028 4576 4077 4604
rect 4028 4564 4034 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 4479 4576 5549 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 4341 4539 4399 4545
rect 4341 4536 4353 4539
rect 1544 4508 2268 4536
rect 2746 4508 4353 4536
rect 1544 4496 1550 4508
rect 2746 4480 2774 4508
rect 4341 4505 4353 4508
rect 4387 4505 4399 4539
rect 4341 4499 4399 4505
rect 4890 4496 4896 4548
rect 4948 4536 4954 4548
rect 5077 4539 5135 4545
rect 4948 4508 4993 4536
rect 4948 4496 4954 4508
rect 5077 4505 5089 4539
rect 5123 4536 5135 4539
rect 5718 4536 5724 4548
rect 5123 4508 5724 4536
rect 5123 4505 5135 4508
rect 5077 4499 5135 4505
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 5920 4545 5948 4644
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 7576 4672 7604 4771
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 11238 4808 11244 4820
rect 11199 4780 11244 4808
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 7834 4700 7840 4752
rect 7892 4740 7898 4752
rect 8021 4743 8079 4749
rect 8021 4740 8033 4743
rect 7892 4712 8033 4740
rect 7892 4700 7898 4712
rect 8021 4709 8033 4712
rect 8067 4709 8079 4743
rect 8021 4703 8079 4709
rect 12161 4743 12219 4749
rect 12161 4709 12173 4743
rect 12207 4740 12219 4743
rect 13262 4740 13268 4752
rect 12207 4712 13268 4740
rect 12207 4709 12219 4712
rect 12161 4703 12219 4709
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 7576 4644 8248 4672
rect 6362 4604 6368 4616
rect 6323 4576 6368 4604
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6454 4564 6460 4616
rect 6512 4604 6518 4616
rect 6512 4576 6557 4604
rect 6512 4564 6518 4576
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 7190 4604 7196 4616
rect 6696 4576 6741 4604
rect 7151 4576 7196 4604
rect 6696 4564 6702 4576
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 7374 4604 7380 4616
rect 7335 4576 7380 4604
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 7576 4604 7604 4644
rect 8220 4613 8248 4644
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9180 4644 9352 4672
rect 9180 4632 9186 4644
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7576 4576 7757 4604
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 9214 4604 9220 4616
rect 9175 4576 9220 4604
rect 8389 4567 8447 4573
rect 5905 4539 5963 4545
rect 5905 4505 5917 4539
rect 5951 4505 5963 4539
rect 5905 4499 5963 4505
rect 5994 4496 6000 4548
rect 6052 4536 6058 4548
rect 6052 4508 6097 4536
rect 6052 4496 6058 4508
rect 6178 4496 6184 4548
rect 6236 4536 6242 4548
rect 6236 4508 6281 4536
rect 6236 4496 6242 4508
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 7944 4536 7972 4567
rect 8404 4536 8432 4567
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9324 4613 9352 4644
rect 10778 4632 10784 4684
rect 10836 4672 10842 4684
rect 11609 4675 11667 4681
rect 11609 4672 11621 4675
rect 10836 4644 11621 4672
rect 10836 4632 10842 4644
rect 11609 4641 11621 4644
rect 11655 4672 11667 4675
rect 11790 4672 11796 4684
rect 11655 4644 11796 4672
rect 11655 4641 11667 4644
rect 11609 4635 11667 4641
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9456 4576 9505 4604
rect 9456 4564 9462 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12768 4576 12817 4604
rect 12768 4564 12774 4576
rect 12805 4573 12817 4576
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4604 13323 4607
rect 13354 4604 13360 4616
rect 13311 4576 13360 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 7156 4508 8432 4536
rect 8573 4539 8631 4545
rect 7156 4496 7162 4508
rect 8573 4505 8585 4539
rect 8619 4536 8631 4539
rect 8662 4536 8668 4548
rect 8619 4508 8668 4536
rect 8619 4505 8631 4508
rect 8573 4499 8631 4505
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 9766 4496 9772 4548
rect 9824 4536 9830 4548
rect 9824 4508 9869 4536
rect 9824 4496 9830 4508
rect 10226 4496 10232 4548
rect 10284 4496 10290 4548
rect 11885 4539 11943 4545
rect 11885 4505 11897 4539
rect 11931 4536 11943 4539
rect 13722 4536 13728 4548
rect 11931 4508 13728 4536
rect 11931 4505 11943 4508
rect 11885 4499 11943 4505
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 2501 4471 2559 4477
rect 2501 4468 2513 4471
rect 2096 4440 2513 4468
rect 2096 4428 2102 4440
rect 2501 4437 2513 4440
rect 2547 4437 2559 4471
rect 2501 4431 2559 4437
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4468 2651 4471
rect 2682 4468 2688 4480
rect 2639 4440 2688 4468
rect 2639 4437 2651 4440
rect 2593 4431 2651 4437
rect 2682 4428 2688 4440
rect 2740 4440 2774 4480
rect 3602 4468 3608 4480
rect 3563 4440 3608 4468
rect 2740 4428 2746 4440
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 4430 4428 4436 4480
rect 4488 4468 4494 4480
rect 4525 4471 4583 4477
rect 4525 4468 4537 4471
rect 4488 4440 4537 4468
rect 4488 4428 4494 4440
rect 4525 4437 4537 4440
rect 4571 4437 4583 4471
rect 4525 4431 4583 4437
rect 4982 4428 4988 4480
rect 5040 4468 5046 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 5040 4440 6561 4468
rect 5040 4428 5046 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 6549 4431 6607 4437
rect 7374 4428 7380 4480
rect 7432 4468 7438 4480
rect 9582 4468 9588 4480
rect 7432 4440 9588 4468
rect 7432 4428 7438 4440
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 11701 4471 11759 4477
rect 11701 4437 11713 4471
rect 11747 4468 11759 4471
rect 12437 4471 12495 4477
rect 12437 4468 12449 4471
rect 11747 4440 12449 4468
rect 11747 4437 11759 4440
rect 11701 4431 11759 4437
rect 12437 4437 12449 4440
rect 12483 4437 12495 4471
rect 12437 4431 12495 4437
rect 1104 4378 13892 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 13892 4378
rect 1104 4304 13892 4326
rect 2685 4267 2743 4273
rect 2685 4233 2697 4267
rect 2731 4264 2743 4267
rect 3142 4264 3148 4276
rect 2731 4236 3148 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 3878 4224 3884 4276
rect 3936 4264 3942 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 3936 4236 4629 4264
rect 3936 4224 3942 4236
rect 4617 4233 4629 4236
rect 4663 4233 4675 4267
rect 4617 4227 4675 4233
rect 6089 4267 6147 4273
rect 6089 4233 6101 4267
rect 6135 4264 6147 4267
rect 9309 4267 9367 4273
rect 6135 4236 7972 4264
rect 6135 4233 6147 4236
rect 6089 4227 6147 4233
rect 1486 4196 1492 4208
rect 1447 4168 1492 4196
rect 1486 4156 1492 4168
rect 1544 4156 1550 4208
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 2924 4168 3188 4196
rect 2924 4156 2930 4168
rect 3160 4140 3188 4168
rect 3602 4156 3608 4208
rect 3660 4196 3666 4208
rect 4982 4196 4988 4208
rect 3660 4168 3740 4196
rect 3660 4156 3666 4168
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 1857 4131 1915 4137
rect 1857 4128 1869 4131
rect 1820 4100 1869 4128
rect 1820 4088 1826 4100
rect 1857 4097 1869 4100
rect 1903 4097 1915 4131
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 1857 4091 1915 4097
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2498 4128 2504 4140
rect 2459 4100 2504 4128
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4128 2835 4131
rect 3050 4128 3056 4140
rect 2823 4100 3056 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3142 4088 3148 4140
rect 3200 4088 3206 4140
rect 3326 4128 3332 4140
rect 3287 4100 3332 4128
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 1946 4060 1952 4072
rect 1907 4032 1952 4060
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2590 4060 2596 4072
rect 2551 4032 2596 4060
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 2866 4060 2872 4072
rect 2827 4032 2872 4060
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 3145 3995 3203 4001
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 3602 3992 3608 4004
rect 3191 3964 3608 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 3602 3952 3608 3964
rect 3660 3952 3666 4004
rect 3712 3992 3740 4168
rect 4356 4168 4988 4196
rect 4356 4137 4384 4168
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 6362 4196 6368 4208
rect 5644 4168 6368 4196
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4614 4128 4620 4140
rect 4575 4100 4620 4128
rect 4341 4091 4399 4097
rect 4172 4060 4200 4091
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 4798 4128 4804 4140
rect 4759 4100 4804 4128
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5166 4128 5172 4140
rect 4948 4100 5172 4128
rect 4948 4088 4954 4100
rect 5166 4088 5172 4100
rect 5224 4128 5230 4140
rect 5644 4137 5672 4168
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 6914 4156 6920 4208
rect 6972 4156 6978 4208
rect 7944 4205 7972 4236
rect 9309 4233 9321 4267
rect 9355 4264 9367 4267
rect 9490 4264 9496 4276
rect 9355 4236 9496 4264
rect 9355 4233 9367 4236
rect 9309 4227 9367 4233
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 9677 4267 9735 4273
rect 9677 4233 9689 4267
rect 9723 4264 9735 4267
rect 9766 4264 9772 4276
rect 9723 4236 9772 4264
rect 9723 4233 9735 4236
rect 9677 4227 9735 4233
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 10468 4236 10517 4264
rect 10468 4224 10474 4236
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 11054 4264 11060 4276
rect 11015 4236 11060 4264
rect 10505 4227 10563 4233
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 11238 4224 11244 4276
rect 11296 4224 11302 4276
rect 7929 4199 7987 4205
rect 7929 4165 7941 4199
rect 7975 4165 7987 4199
rect 9398 4196 9404 4208
rect 7929 4159 7987 4165
rect 8220 4168 9404 4196
rect 8220 4140 8248 4168
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 10321 4199 10379 4205
rect 10321 4196 10333 4199
rect 9784 4168 10333 4196
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 5224 4100 5273 4128
rect 5224 4088 5230 4100
rect 5261 4097 5273 4100
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 5902 4128 5908 4140
rect 5859 4100 5908 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8260 4100 8305 4128
rect 8260 4088 8266 4100
rect 8570 4088 8576 4140
rect 8628 4128 8634 4140
rect 8757 4131 8815 4137
rect 8757 4128 8769 4131
rect 8628 4100 8769 4128
rect 8628 4088 8634 4100
rect 8757 4097 8769 4100
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9784 4128 9812 4168
rect 10321 4165 10333 4168
rect 10367 4196 10379 4199
rect 11256 4196 11284 4224
rect 10367 4168 11284 4196
rect 10367 4165 10379 4168
rect 10321 4159 10379 4165
rect 11882 4156 11888 4208
rect 11940 4196 11946 4208
rect 11940 4168 12282 4196
rect 11940 4156 11946 4168
rect 9171 4100 9812 4128
rect 9861 4131 9919 4137
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 10597 4131 10655 4137
rect 9907 4100 10088 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 5074 4060 5080 4072
rect 4172 4032 5080 4060
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 5718 4060 5724 4072
rect 5491 4032 5724 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4060 6239 4063
rect 6730 4060 6736 4072
rect 6227 4032 6736 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6730 4020 6736 4032
rect 6788 4020 6794 4072
rect 7282 4020 7288 4072
rect 7340 4060 7346 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 7340 4032 8677 4060
rect 7340 4020 7346 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 9766 4060 9772 4072
rect 8665 4023 8723 4029
rect 9646 4032 9772 4060
rect 5258 3992 5264 4004
rect 3712 3964 5264 3992
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 5736 3992 5764 4020
rect 6457 3995 6515 4001
rect 6457 3992 6469 3995
rect 5736 3964 6469 3992
rect 6457 3961 6469 3964
rect 6503 3992 6515 3995
rect 6546 3992 6552 4004
rect 6503 3964 6552 3992
rect 6503 3961 6515 3964
rect 6457 3955 6515 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 9646 3992 9674 4032
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 10060 4001 10088 4100
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 10778 4128 10784 4140
rect 10643 4100 10784 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11238 4128 11244 4140
rect 11199 4100 11244 4128
rect 11057 4091 11115 4097
rect 8128 3964 9674 3992
rect 10045 3995 10103 4001
rect 2958 3924 2964 3936
rect 2919 3896 2964 3924
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4672 3896 5089 3924
rect 4672 3884 4678 3896
rect 5077 3893 5089 3896
rect 5123 3924 5135 3927
rect 6638 3924 6644 3936
rect 5123 3896 6644 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 8128 3924 8156 3964
rect 10045 3961 10057 3995
rect 10091 3961 10103 3995
rect 10045 3955 10103 3961
rect 6880 3896 8156 3924
rect 9125 3927 9183 3933
rect 6880 3884 6886 3896
rect 9125 3893 9137 3927
rect 9171 3924 9183 3927
rect 9214 3924 9220 3936
rect 9171 3896 9220 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 11072 3924 11100 4091
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11388 4032 11529 4060
rect 11388 4020 11394 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11517 4023 11575 4029
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 13446 4060 13452 4072
rect 11839 4032 13452 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13170 3952 13176 4004
rect 13228 3992 13234 4004
rect 13265 3995 13323 4001
rect 13265 3992 13277 3995
rect 13228 3964 13277 3992
rect 13228 3952 13234 3964
rect 13265 3961 13277 3964
rect 13311 3961 13323 3995
rect 13265 3955 13323 3961
rect 11514 3924 11520 3936
rect 11072 3896 11520 3924
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 1104 3834 13892 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 13892 3834
rect 1104 3760 13892 3782
rect 1857 3723 1915 3729
rect 1857 3689 1869 3723
rect 1903 3720 1915 3723
rect 1946 3720 1952 3732
rect 1903 3692 1952 3720
rect 1903 3689 1915 3692
rect 1857 3683 1915 3689
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 2041 3723 2099 3729
rect 2041 3689 2053 3723
rect 2087 3720 2099 3723
rect 2866 3720 2872 3732
rect 2087 3692 2872 3720
rect 2087 3689 2099 3692
rect 2041 3683 2099 3689
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3689 3295 3723
rect 3510 3720 3516 3732
rect 3471 3692 3516 3720
rect 3237 3683 3295 3689
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 2317 3655 2375 3661
rect 2317 3652 2329 3655
rect 1728 3624 2329 3652
rect 1728 3612 1734 3624
rect 2317 3621 2329 3624
rect 2363 3621 2375 3655
rect 2317 3615 2375 3621
rect 2498 3612 2504 3664
rect 2556 3652 2562 3664
rect 3252 3652 3280 3683
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 3970 3720 3976 3732
rect 3931 3692 3976 3720
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 5074 3720 5080 3732
rect 5035 3692 5080 3720
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 5684 3692 6377 3720
rect 5684 3680 5690 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 6365 3683 6423 3689
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7926 3720 7932 3732
rect 7064 3692 7932 3720
rect 7064 3680 7070 3692
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 9950 3720 9956 3732
rect 9911 3692 9956 3720
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 10100 3692 10149 3720
rect 10100 3680 10106 3692
rect 10137 3689 10149 3692
rect 10183 3720 10195 3723
rect 10962 3720 10968 3732
rect 10183 3692 10968 3720
rect 10183 3689 10195 3692
rect 10137 3683 10195 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 12529 3723 12587 3729
rect 12529 3689 12541 3723
rect 12575 3720 12587 3723
rect 12618 3720 12624 3732
rect 12575 3692 12624 3720
rect 12575 3689 12587 3692
rect 12529 3683 12587 3689
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 2556 3624 3280 3652
rect 5905 3655 5963 3661
rect 2556 3612 2562 3624
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 5994 3652 6000 3664
rect 5951 3624 6000 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 6178 3652 6184 3664
rect 6139 3624 6184 3652
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 9030 3652 9036 3664
rect 6788 3624 8892 3652
rect 8991 3624 9036 3652
rect 6788 3612 6794 3624
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 2038 3584 2044 3596
rect 1627 3556 2044 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 2038 3544 2044 3556
rect 2096 3584 2102 3596
rect 2869 3587 2927 3593
rect 2096 3556 2544 3584
rect 2096 3544 2102 3556
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2130 3516 2136 3528
rect 1903 3488 2136 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 1688 3448 1716 3479
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2516 3525 2544 3556
rect 2869 3553 2881 3587
rect 2915 3584 2927 3587
rect 3142 3584 3148 3596
rect 2915 3556 3148 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 4338 3584 4344 3596
rect 4172 3556 4344 3584
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3234 3516 3240 3528
rect 2832 3488 2877 3516
rect 3195 3488 3240 3516
rect 2832 3476 2838 3488
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 4172 3525 4200 3556
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 5442 3584 5448 3596
rect 5355 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3584 5506 3596
rect 6914 3584 6920 3596
rect 5500 3556 6776 3584
rect 6875 3556 6920 3584
rect 5500 3544 5506 3556
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4430 3516 4436 3528
rect 4304 3488 4349 3516
rect 4391 3488 4436 3516
rect 4304 3476 4310 3488
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4580 3488 4905 3516
rect 4580 3476 4586 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 5626 3516 5632 3528
rect 5587 3488 5632 3516
rect 4893 3479 4951 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5868 3488 6009 3516
rect 5868 3476 5874 3488
rect 5997 3485 6009 3488
rect 6043 3485 6055 3519
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 5997 3479 6055 3485
rect 6104 3488 6653 3516
rect 1762 3448 1768 3460
rect 1675 3420 1768 3448
rect 1762 3408 1768 3420
rect 1820 3448 1826 3460
rect 1820 3420 2820 3448
rect 1820 3408 1826 3420
rect 2792 3392 2820 3420
rect 2958 3408 2964 3460
rect 3016 3448 3022 3460
rect 3326 3448 3332 3460
rect 3016 3420 3332 3448
rect 3016 3408 3022 3420
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 4338 3408 4344 3460
rect 4396 3448 4402 3460
rect 4617 3451 4675 3457
rect 4617 3448 4629 3451
rect 4396 3420 4629 3448
rect 4396 3408 4402 3420
rect 4617 3417 4629 3420
rect 4663 3448 4675 3451
rect 4798 3448 4804 3460
rect 4663 3420 4804 3448
rect 4663 3417 4675 3420
rect 4617 3411 4675 3417
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 4982 3408 4988 3460
rect 5040 3448 5046 3460
rect 6104 3448 6132 3488
rect 6641 3485 6653 3488
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 6546 3448 6552 3460
rect 5040 3420 6132 3448
rect 6507 3420 6552 3448
rect 5040 3408 5046 3420
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 2774 3340 2780 3392
rect 2832 3340 2838 3392
rect 3050 3380 3056 3392
rect 3011 3352 3056 3380
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 3510 3380 3516 3392
rect 3200 3352 3516 3380
rect 3200 3340 3206 3352
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 4706 3380 4712 3392
rect 4304 3352 4712 3380
rect 4304 3340 4310 3352
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 5350 3340 5356 3392
rect 5408 3380 5414 3392
rect 5810 3380 5816 3392
rect 5408 3352 5816 3380
rect 5408 3340 5414 3352
rect 5810 3340 5816 3352
rect 5868 3340 5874 3392
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3380 6423 3383
rect 6748 3380 6776 3556
rect 6914 3544 6920 3556
rect 6972 3544 6978 3596
rect 7558 3584 7564 3596
rect 7208 3556 7564 3584
rect 7006 3516 7012 3528
rect 6967 3488 7012 3516
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 7208 3525 7236 3556
rect 7558 3544 7564 3556
rect 7616 3584 7622 3596
rect 8018 3584 8024 3596
rect 7616 3556 8024 3584
rect 7616 3544 7622 3556
rect 8018 3544 8024 3556
rect 8076 3584 8082 3596
rect 8076 3556 8156 3584
rect 8076 3544 8082 3556
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7926 3516 7932 3528
rect 7887 3488 7932 3516
rect 7377 3479 7435 3485
rect 7392 3392 7420 3479
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8128 3525 8156 3556
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 8159 3488 8401 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 8662 3516 8668 3528
rect 8619 3488 8668 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 7558 3448 7564 3460
rect 7519 3420 7564 3448
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 7745 3451 7803 3457
rect 7745 3417 7757 3451
rect 7791 3448 7803 3451
rect 7834 3448 7840 3460
rect 7791 3420 7840 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 7944 3448 7972 3476
rect 8588 3448 8616 3479
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 8754 3448 8760 3460
rect 7944 3420 8616 3448
rect 8715 3420 8760 3448
rect 8754 3408 8760 3420
rect 8812 3408 8818 3460
rect 8864 3448 8892 3624
rect 9030 3612 9036 3624
rect 9088 3612 9094 3664
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 13173 3655 13231 3661
rect 13173 3652 13185 3655
rect 13044 3624 13185 3652
rect 13044 3612 13050 3624
rect 13173 3621 13185 3624
rect 13219 3621 13231 3655
rect 13173 3615 13231 3621
rect 10134 3544 10140 3596
rect 10192 3584 10198 3596
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 10192 3556 10517 3584
rect 10192 3544 10198 3556
rect 10505 3553 10517 3556
rect 10551 3584 10563 3587
rect 11330 3584 11336 3596
rect 10551 3556 11336 3584
rect 10551 3553 10563 3556
rect 10505 3547 10563 3553
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 12710 3516 12716 3528
rect 11914 3488 12716 3516
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 12894 3516 12900 3528
rect 12855 3488 12900 3516
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13078 3516 13084 3528
rect 13039 3488 13084 3516
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 9585 3451 9643 3457
rect 9585 3448 9597 3451
rect 8864 3420 9597 3448
rect 9585 3417 9597 3420
rect 9631 3448 9643 3451
rect 10137 3451 10195 3457
rect 10137 3448 10149 3451
rect 9631 3420 10149 3448
rect 9631 3417 9643 3420
rect 9585 3411 9643 3417
rect 10137 3417 10149 3420
rect 10183 3417 10195 3451
rect 10137 3411 10195 3417
rect 10321 3451 10379 3457
rect 10321 3417 10333 3451
rect 10367 3448 10379 3451
rect 10410 3448 10416 3460
rect 10367 3420 10416 3448
rect 10367 3417 10379 3420
rect 10321 3411 10379 3417
rect 7282 3380 7288 3392
rect 6411 3352 7288 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7374 3340 7380 3392
rect 7432 3340 7438 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 7929 3383 7987 3389
rect 7929 3380 7941 3383
rect 7524 3352 7941 3380
rect 7524 3340 7530 3352
rect 7929 3349 7941 3352
rect 7975 3349 7987 3383
rect 7929 3343 7987 3349
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3380 9551 3383
rect 10042 3380 10048 3392
rect 9539 3352 10048 3380
rect 9539 3349 9551 3352
rect 9493 3343 9551 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 10152 3380 10180 3411
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 10778 3448 10784 3460
rect 10739 3420 10784 3448
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 12621 3451 12679 3457
rect 12621 3417 12633 3451
rect 12667 3417 12679 3451
rect 12802 3448 12808 3460
rect 12763 3420 12808 3448
rect 12621 3411 12679 3417
rect 11146 3380 11152 3392
rect 10152 3352 11152 3380
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 12526 3380 12532 3392
rect 12299 3352 12532 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 12636 3380 12664 3411
rect 12802 3408 12808 3420
rect 12860 3408 12866 3460
rect 13170 3380 13176 3392
rect 12636 3352 13176 3380
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 1104 3290 13892 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 13892 3290
rect 1104 3216 13892 3238
rect 1857 3179 1915 3185
rect 1857 3145 1869 3179
rect 1903 3176 1915 3179
rect 3234 3176 3240 3188
rect 1903 3148 3240 3176
rect 1903 3145 1915 3148
rect 1857 3139 1915 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3329 3179 3387 3185
rect 3329 3145 3341 3179
rect 3375 3176 3387 3179
rect 4522 3176 4528 3188
rect 3375 3148 4528 3176
rect 3375 3145 3387 3148
rect 3329 3139 3387 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 5074 3176 5080 3188
rect 5035 3148 5080 3176
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 5592 3148 6561 3176
rect 5592 3136 5598 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 7377 3179 7435 3185
rect 7377 3176 7389 3179
rect 6696 3148 7389 3176
rect 6696 3136 6702 3148
rect 7377 3145 7389 3148
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8386 3176 8392 3188
rect 8076 3148 8392 3176
rect 8076 3136 8082 3148
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9769 3179 9827 3185
rect 9769 3176 9781 3179
rect 9364 3148 9781 3176
rect 9364 3136 9370 3148
rect 9769 3145 9781 3148
rect 9815 3176 9827 3179
rect 13446 3176 13452 3188
rect 9815 3148 10364 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 2774 3108 2780 3120
rect 1596 3080 2452 3108
rect 2735 3080 2780 3108
rect 1596 3052 1624 3080
rect 2424 3052 2452 3080
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 3789 3111 3847 3117
rect 3789 3108 3801 3111
rect 3436 3080 3801 3108
rect 1578 3040 1584 3052
rect 1491 3012 1584 3040
rect 1578 3000 1584 3012
rect 1636 3000 1642 3052
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 1719 3012 2329 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 1854 2932 1860 2984
rect 1912 2972 1918 2984
rect 2133 2975 2191 2981
rect 2133 2972 2145 2975
rect 1912 2944 2145 2972
rect 1912 2932 1918 2944
rect 2133 2941 2145 2944
rect 2179 2941 2191 2975
rect 2133 2935 2191 2941
rect 2332 2836 2360 3003
rect 2406 3000 2412 3052
rect 2464 3040 2470 3052
rect 2958 3040 2964 3052
rect 2464 3012 2509 3040
rect 2919 3012 2964 3040
rect 2464 3000 2470 3012
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 2682 2972 2688 2984
rect 2643 2944 2688 2972
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 2792 2944 3004 2972
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2904 2651 2907
rect 2792 2904 2820 2944
rect 2639 2876 2820 2904
rect 2976 2904 3004 2944
rect 3050 2932 3056 2984
rect 3108 2972 3114 2984
rect 3160 2972 3188 3003
rect 3108 2944 3188 2972
rect 3108 2932 3114 2944
rect 3436 2904 3464 3080
rect 3789 3077 3801 3080
rect 3835 3077 3847 3111
rect 7561 3111 7619 3117
rect 7561 3108 7573 3111
rect 3789 3071 3847 3077
rect 4172 3080 7573 3108
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3602 3040 3608 3052
rect 3559 3012 3608 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 3697 2975 3755 2981
rect 3697 2941 3709 2975
rect 3743 2972 3755 2975
rect 4062 2972 4068 2984
rect 3743 2944 4068 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 3510 2904 3516 2916
rect 2976 2876 3516 2904
rect 2639 2873 2651 2876
rect 2593 2867 2651 2873
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 4172 2836 4200 3080
rect 7561 3077 7573 3080
rect 7607 3077 7619 3111
rect 7561 3071 7619 3077
rect 8297 3111 8355 3117
rect 8297 3077 8309 3111
rect 8343 3108 8355 3111
rect 8570 3108 8576 3120
rect 8343 3080 8576 3108
rect 8343 3077 8355 3080
rect 8297 3071 8355 3077
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 8754 3068 8760 3120
rect 8812 3068 8818 3120
rect 10336 3117 10364 3148
rect 11164 3148 12112 3176
rect 13407 3148 13452 3176
rect 11164 3120 11192 3148
rect 10321 3111 10379 3117
rect 10321 3077 10333 3111
rect 10367 3077 10379 3111
rect 10321 3071 10379 3077
rect 10410 3068 10416 3120
rect 10468 3108 10474 3120
rect 10505 3111 10563 3117
rect 10505 3108 10517 3111
rect 10468 3080 10517 3108
rect 10468 3068 10474 3080
rect 10505 3077 10517 3080
rect 10551 3077 10563 3111
rect 11146 3108 11152 3120
rect 11107 3080 11152 3108
rect 10505 3071 10563 3077
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 11238 3068 11244 3120
rect 11296 3108 11302 3120
rect 11422 3108 11428 3120
rect 11296 3080 11428 3108
rect 11296 3068 11302 3080
rect 11422 3068 11428 3080
rect 11480 3108 11486 3120
rect 11882 3108 11888 3120
rect 11480 3080 11744 3108
rect 11843 3080 11888 3108
rect 11480 3068 11486 3080
rect 4614 3040 4620 3052
rect 4575 3012 4620 3040
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4798 3040 4804 3052
rect 4759 3012 4804 3040
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5092 2972 5120 3003
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5442 3040 5448 3052
rect 5224 3012 5269 3040
rect 5403 3012 5448 3040
rect 5224 3000 5230 3012
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5994 3040 6000 3052
rect 5955 3012 6000 3040
rect 5721 3003 5779 3009
rect 5350 2972 5356 2984
rect 5092 2944 5356 2972
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 5626 2972 5632 2984
rect 5587 2944 5632 2972
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 4890 2864 4896 2916
rect 4948 2904 4954 2916
rect 5736 2904 5764 3003
rect 5994 3000 6000 3012
rect 6052 3040 6058 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6052 3012 6561 3040
rect 6052 3000 6058 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6788 3012 6929 3040
rect 6788 3000 6794 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 7098 3040 7104 3052
rect 7059 3012 7104 3040
rect 6917 3003 6975 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7374 3040 7380 3052
rect 7239 3012 7380 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7834 3040 7840 3052
rect 7795 3012 7840 3040
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 10962 3040 10968 3052
rect 10923 3012 10968 3040
rect 10962 3000 10968 3012
rect 11020 3000 11026 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 11716 3049 11744 3080
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 12084 3117 12112 3148
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 12069 3111 12127 3117
rect 12069 3077 12081 3111
rect 12115 3077 12127 3111
rect 12069 3071 12127 3077
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12618 3000 12624 3052
rect 12676 3000 12682 3052
rect 13262 3040 13268 3052
rect 13223 3012 13268 3040
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 6362 2972 6368 2984
rect 6323 2944 6368 2972
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 7282 2932 7288 2984
rect 7340 2972 7346 2984
rect 8018 2972 8024 2984
rect 7340 2944 8024 2972
rect 7340 2932 7346 2944
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 11238 2972 11244 2984
rect 10643 2944 11244 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 5994 2904 6000 2916
rect 4948 2876 6000 2904
rect 4948 2864 4954 2876
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 9306 2864 9312 2916
rect 9364 2904 9370 2916
rect 10781 2907 10839 2913
rect 10781 2904 10793 2907
rect 9364 2876 10793 2904
rect 9364 2864 9370 2876
rect 10781 2873 10793 2876
rect 10827 2873 10839 2907
rect 10781 2867 10839 2873
rect 10870 2864 10876 2916
rect 10928 2904 10934 2916
rect 12912 2904 12940 2935
rect 10928 2876 12940 2904
rect 10928 2864 10934 2876
rect 2332 2808 4200 2836
rect 5074 2796 5080 2848
rect 5132 2836 5138 2848
rect 6454 2836 6460 2848
rect 5132 2808 6460 2836
rect 5132 2796 5138 2808
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 10045 2839 10103 2845
rect 10045 2836 10057 2839
rect 10008 2808 10057 2836
rect 10008 2796 10014 2808
rect 10045 2805 10057 2808
rect 10091 2805 10103 2839
rect 10045 2799 10103 2805
rect 1104 2746 13892 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 13892 2746
rect 1104 2672 13892 2694
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 6730 2632 6736 2644
rect 5123 2604 6736 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 7650 2592 7656 2644
rect 7708 2632 7714 2644
rect 7745 2635 7803 2641
rect 7745 2632 7757 2635
rect 7708 2604 7757 2632
rect 7708 2592 7714 2604
rect 7745 2601 7757 2604
rect 7791 2601 7803 2635
rect 7745 2595 7803 2601
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 10962 2632 10968 2644
rect 10735 2604 10968 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11698 2592 11704 2644
rect 11756 2632 11762 2644
rect 11756 2604 12756 2632
rect 11756 2592 11762 2604
rect 4982 2564 4988 2576
rect 3528 2536 4988 2564
rect 2682 2456 2688 2508
rect 2740 2496 2746 2508
rect 3528 2496 3556 2536
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 7466 2564 7472 2576
rect 6748 2536 7472 2564
rect 2740 2468 3556 2496
rect 2740 2456 2746 2468
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 2590 2428 2596 2440
rect 1728 2400 2596 2428
rect 1728 2388 1734 2400
rect 2590 2388 2596 2400
rect 2648 2428 2654 2440
rect 3436 2437 3464 2468
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4798 2496 4804 2508
rect 4120 2468 4165 2496
rect 4759 2468 4804 2496
rect 4120 2456 4126 2468
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5360 2499 5418 2505
rect 5360 2465 5372 2499
rect 5406 2465 5418 2499
rect 5360 2459 5418 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 5718 2496 5724 2508
rect 5675 2468 5724 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 2648 2400 3249 2428
rect 2648 2388 2654 2400
rect 3237 2397 3249 2400
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 3510 2388 3516 2440
rect 3568 2428 3574 2440
rect 3568 2400 3613 2428
rect 3568 2388 3574 2400
rect 2038 2320 2044 2372
rect 2096 2360 2102 2372
rect 3145 2363 3203 2369
rect 3145 2360 3157 2363
rect 2096 2332 3157 2360
rect 2096 2320 2102 2332
rect 3145 2329 3157 2332
rect 3191 2329 3203 2363
rect 3145 2323 3203 2329
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 2774 2292 2780 2304
rect 1903 2264 2780 2292
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 3160 2292 3188 2323
rect 3602 2320 3608 2372
rect 3660 2360 3666 2372
rect 3988 2360 4016 2414
rect 5074 2388 5080 2440
rect 5132 2428 5138 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 5132 2400 5273 2428
rect 5132 2388 5138 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 3660 2332 4016 2360
rect 3660 2320 3666 2332
rect 5368 2292 5396 2459
rect 5718 2456 5724 2468
rect 5776 2456 5782 2508
rect 6748 2414 6776 2536
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 11330 2524 11336 2576
rect 11388 2524 11394 2576
rect 12728 2564 12756 2604
rect 12728 2536 12848 2564
rect 7650 2456 7656 2508
rect 7708 2496 7714 2508
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 7708 2468 7941 2496
rect 7708 2456 7714 2468
rect 7929 2465 7941 2468
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 8110 2456 8116 2508
rect 8168 2496 8174 2508
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8168 2468 8953 2496
rect 8168 2456 8174 2468
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 11348 2496 11376 2524
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 11348 2468 12725 2496
rect 8941 2459 8999 2465
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 7558 2428 7564 2440
rect 7519 2400 7564 2428
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 6932 2332 7297 2360
rect 5810 2292 5816 2304
rect 3160 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 6270 2252 6276 2304
rect 6328 2292 6334 2304
rect 6932 2292 6960 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7285 2323 7343 2329
rect 7374 2320 7380 2372
rect 7432 2360 7438 2372
rect 7760 2360 7788 2391
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7892 2400 8033 2428
rect 7892 2388 7898 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 7432 2332 7788 2360
rect 7432 2320 7438 2332
rect 7926 2320 7932 2372
rect 7984 2360 7990 2372
rect 8312 2360 8340 2391
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8662 2428 8668 2440
rect 8444 2400 8489 2428
rect 8623 2400 8668 2428
rect 8444 2388 8450 2400
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 12820 2437 12848 2536
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2397 12863 2431
rect 13078 2428 13084 2440
rect 13039 2400 13084 2428
rect 12805 2391 12863 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 9214 2360 9220 2372
rect 7984 2332 8340 2360
rect 9175 2332 9220 2360
rect 7984 2320 7990 2332
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 9324 2332 9706 2360
rect 7098 2292 7104 2304
rect 6328 2264 6960 2292
rect 7059 2264 7104 2292
rect 6328 2252 6334 2264
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 8665 2295 8723 2301
rect 8665 2261 8677 2295
rect 8711 2292 8723 2295
rect 9324 2292 9352 2332
rect 11054 2320 11060 2372
rect 11112 2360 11118 2372
rect 12437 2363 12495 2369
rect 11112 2332 11270 2360
rect 11112 2320 11118 2332
rect 12437 2329 12449 2363
rect 12483 2360 12495 2363
rect 13262 2360 13268 2372
rect 12483 2332 13268 2360
rect 12483 2329 12495 2332
rect 12437 2323 12495 2329
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 10962 2292 10968 2304
rect 8711 2264 9352 2292
rect 10923 2264 10968 2292
rect 8711 2261 8723 2264
rect 8665 2255 8723 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 12710 2252 12716 2304
rect 12768 2292 12774 2304
rect 12897 2295 12955 2301
rect 12897 2292 12909 2295
rect 12768 2264 12909 2292
rect 12768 2252 12774 2264
rect 12897 2261 12909 2264
rect 12943 2261 12955 2295
rect 12897 2255 12955 2261
rect 1104 2202 13892 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 13892 2202
rect 1104 2128 13892 2150
rect 1489 2091 1547 2097
rect 1489 2057 1501 2091
rect 1535 2088 1547 2091
rect 2682 2088 2688 2100
rect 1535 2060 2688 2088
rect 1535 2057 1547 2060
rect 1489 2051 1547 2057
rect 2682 2048 2688 2060
rect 2740 2048 2746 2100
rect 3602 2048 3608 2100
rect 3660 2088 3666 2100
rect 3789 2091 3847 2097
rect 3789 2088 3801 2091
rect 3660 2060 3801 2088
rect 3660 2048 3666 2060
rect 3789 2057 3801 2060
rect 3835 2057 3847 2091
rect 4062 2088 4068 2100
rect 4023 2060 4068 2088
rect 3789 2051 3847 2057
rect 4062 2048 4068 2060
rect 4120 2048 4126 2100
rect 7650 2088 7656 2100
rect 4264 2060 7656 2088
rect 4264 2020 4292 2060
rect 7650 2048 7656 2060
rect 7708 2048 7714 2100
rect 9582 2048 9588 2100
rect 9640 2088 9646 2100
rect 10410 2088 10416 2100
rect 9640 2060 10272 2088
rect 10371 2060 10416 2088
rect 9640 2048 9646 2060
rect 3542 1992 4292 2020
rect 4982 1980 4988 2032
rect 5040 1980 5046 2032
rect 5534 2020 5540 2032
rect 5495 1992 5540 2020
rect 5534 1980 5540 1992
rect 5592 1980 5598 2032
rect 6730 2020 6736 2032
rect 5828 1992 6408 2020
rect 6691 1992 6736 2020
rect 5828 1964 5856 1992
rect 1670 1952 1676 1964
rect 1631 1924 1676 1952
rect 1670 1912 1676 1924
rect 1728 1912 1734 1964
rect 1854 1952 1860 1964
rect 1815 1924 1860 1952
rect 1854 1912 1860 1924
rect 1912 1912 1918 1964
rect 2038 1952 2044 1964
rect 1999 1924 2044 1952
rect 2038 1912 2044 1924
rect 2096 1912 2102 1964
rect 5810 1912 5816 1964
rect 5868 1952 5874 1964
rect 6181 1955 6239 1961
rect 5868 1924 5913 1952
rect 5868 1912 5874 1924
rect 6181 1921 6193 1955
rect 6227 1921 6239 1955
rect 6181 1915 6239 1921
rect 2317 1887 2375 1893
rect 2317 1853 2329 1887
rect 2363 1884 2375 1887
rect 3326 1884 3332 1896
rect 2363 1856 3332 1884
rect 2363 1853 2375 1856
rect 2317 1847 2375 1853
rect 3326 1844 3332 1856
rect 3384 1844 3390 1896
rect 1857 1751 1915 1757
rect 1857 1717 1869 1751
rect 1903 1748 1915 1751
rect 2498 1748 2504 1760
rect 1903 1720 2504 1748
rect 1903 1717 1915 1720
rect 1857 1711 1915 1717
rect 2498 1708 2504 1720
rect 2556 1708 2562 1760
rect 5994 1748 6000 1760
rect 5955 1720 6000 1748
rect 5994 1708 6000 1720
rect 6052 1708 6058 1760
rect 6196 1748 6224 1915
rect 6380 1884 6408 1992
rect 6730 1980 6736 1992
rect 6788 1980 6794 2032
rect 7742 1980 7748 2032
rect 7800 1980 7806 2032
rect 9674 1980 9680 2032
rect 9732 1980 9738 2032
rect 8018 1912 8024 1964
rect 8076 1952 8082 1964
rect 8665 1955 8723 1961
rect 8665 1952 8677 1955
rect 8076 1924 8677 1952
rect 8076 1912 8082 1924
rect 8665 1921 8677 1924
rect 8711 1921 8723 1955
rect 10244 1952 10272 2060
rect 10410 2048 10416 2060
rect 10468 2048 10474 2100
rect 11054 2088 11060 2100
rect 11015 2060 11060 2088
rect 11054 2048 11060 2060
rect 11112 2048 11118 2100
rect 11238 2048 11244 2100
rect 11296 2048 11302 2100
rect 11422 2048 11428 2100
rect 11480 2088 11486 2100
rect 13078 2088 13084 2100
rect 11480 2060 13084 2088
rect 11480 2048 11486 2060
rect 13078 2048 13084 2060
rect 13136 2048 13142 2100
rect 13262 2088 13268 2100
rect 13223 2060 13268 2088
rect 13262 2048 13268 2060
rect 13320 2048 13326 2100
rect 11256 2020 11284 2048
rect 11790 2020 11796 2032
rect 11256 1992 11796 2020
rect 11790 1980 11796 1992
rect 11848 1980 11854 2032
rect 11882 1980 11888 2032
rect 11940 2020 11946 2032
rect 11940 1992 12282 2020
rect 11940 1980 11946 1992
rect 10873 1955 10931 1961
rect 10873 1952 10885 1955
rect 10244 1924 10885 1952
rect 8665 1915 8723 1921
rect 10873 1921 10885 1924
rect 10919 1921 10931 1955
rect 10873 1915 10931 1921
rect 10965 1955 11023 1961
rect 10965 1921 10977 1955
rect 11011 1921 11023 1955
rect 11238 1952 11244 1964
rect 11199 1924 11244 1952
rect 10965 1915 11023 1921
rect 6457 1887 6515 1893
rect 6457 1884 6469 1887
rect 6380 1856 6469 1884
rect 6457 1853 6469 1856
rect 6503 1884 6515 1887
rect 7282 1884 7288 1896
rect 6503 1856 7288 1884
rect 6503 1853 6515 1856
rect 6457 1847 6515 1853
rect 7282 1844 7288 1856
rect 7340 1844 7346 1896
rect 7374 1844 7380 1896
rect 7432 1884 7438 1896
rect 8205 1887 8263 1893
rect 8205 1884 8217 1887
rect 7432 1856 8217 1884
rect 7432 1844 7438 1856
rect 8205 1853 8217 1856
rect 8251 1853 8263 1887
rect 8938 1884 8944 1896
rect 8899 1856 8944 1884
rect 8205 1847 8263 1853
rect 8938 1844 8944 1856
rect 8996 1844 9002 1896
rect 10980 1884 11008 1915
rect 11238 1912 11244 1924
rect 11296 1912 11302 1964
rect 11330 1912 11336 1964
rect 11388 1952 11394 1964
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 11388 1924 11529 1952
rect 11388 1912 11394 1924
rect 11517 1921 11529 1924
rect 11563 1921 11575 1955
rect 11517 1915 11575 1921
rect 11054 1884 11060 1896
rect 10704 1856 11060 1884
rect 7466 1748 7472 1760
rect 6196 1720 7472 1748
rect 7466 1708 7472 1720
rect 7524 1708 7530 1760
rect 7926 1708 7932 1760
rect 7984 1748 7990 1760
rect 10704 1757 10732 1856
rect 11054 1844 11060 1856
rect 11112 1844 11118 1896
rect 11793 1887 11851 1893
rect 11793 1884 11805 1887
rect 11164 1856 11805 1884
rect 11164 1828 11192 1856
rect 11793 1853 11805 1856
rect 11839 1853 11851 1887
rect 11793 1847 11851 1853
rect 11146 1776 11152 1828
rect 11204 1776 11210 1828
rect 10689 1751 10747 1757
rect 10689 1748 10701 1751
rect 7984 1720 10701 1748
rect 7984 1708 7990 1720
rect 10689 1717 10701 1720
rect 10735 1717 10747 1751
rect 10689 1711 10747 1717
rect 1104 1658 13892 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 13892 1658
rect 1104 1584 13892 1606
rect 3326 1544 3332 1556
rect 3287 1516 3332 1544
rect 3326 1504 3332 1516
rect 3384 1504 3390 1556
rect 7466 1504 7472 1556
rect 7524 1544 7530 1556
rect 9033 1547 9091 1553
rect 7524 1516 7880 1544
rect 7524 1504 7530 1516
rect 2866 1476 2872 1488
rect 2827 1448 2872 1476
rect 2866 1436 2872 1448
rect 2924 1436 2930 1488
rect 5074 1436 5080 1488
rect 5132 1476 5138 1488
rect 6917 1479 6975 1485
rect 6917 1476 6929 1479
rect 5132 1448 6929 1476
rect 5132 1436 5138 1448
rect 6917 1445 6929 1448
rect 6963 1445 6975 1479
rect 7742 1476 7748 1488
rect 7703 1448 7748 1476
rect 6917 1439 6975 1445
rect 7742 1436 7748 1448
rect 7800 1436 7806 1488
rect 7852 1476 7880 1516
rect 9033 1513 9045 1547
rect 9079 1544 9091 1547
rect 9214 1544 9220 1556
rect 9079 1516 9220 1544
rect 9079 1513 9091 1516
rect 9033 1507 9091 1513
rect 9214 1504 9220 1516
rect 9272 1504 9278 1556
rect 7852 1448 11836 1476
rect 11808 1420 11836 1448
rect 3602 1368 3608 1420
rect 3660 1408 3666 1420
rect 4433 1411 4491 1417
rect 3660 1380 4292 1408
rect 3660 1368 3666 1380
rect 1394 1340 1400 1352
rect 1355 1312 1400 1340
rect 1394 1300 1400 1312
rect 1452 1300 1458 1352
rect 3513 1343 3571 1349
rect 3513 1309 3525 1343
rect 3559 1340 3571 1343
rect 3863 1343 3921 1349
rect 3863 1340 3875 1343
rect 3559 1312 3875 1340
rect 3559 1309 3571 1312
rect 3513 1303 3571 1309
rect 3863 1309 3875 1312
rect 3909 1309 3921 1343
rect 3863 1303 3921 1309
rect 4062 1232 4068 1284
rect 4120 1272 4126 1284
rect 4157 1275 4215 1281
rect 4157 1272 4169 1275
rect 4120 1244 4169 1272
rect 4120 1232 4126 1244
rect 4157 1241 4169 1244
rect 4203 1241 4215 1275
rect 4264 1272 4292 1380
rect 4433 1377 4445 1411
rect 4479 1408 4491 1411
rect 5994 1408 6000 1420
rect 4479 1380 6000 1408
rect 4479 1377 4491 1380
rect 4433 1371 4491 1377
rect 5994 1368 6000 1380
rect 6052 1368 6058 1420
rect 6181 1411 6239 1417
rect 6181 1377 6193 1411
rect 6227 1408 6239 1411
rect 6362 1408 6368 1420
rect 6227 1380 6368 1408
rect 6227 1377 6239 1380
rect 6181 1371 6239 1377
rect 6362 1368 6368 1380
rect 6420 1368 6426 1420
rect 7377 1411 7435 1417
rect 7377 1408 7389 1411
rect 7208 1380 7389 1408
rect 4706 1340 4712 1352
rect 4667 1312 4712 1340
rect 4706 1300 4712 1312
rect 4764 1300 4770 1352
rect 4798 1300 4804 1352
rect 4856 1340 4862 1352
rect 4982 1340 4988 1352
rect 4856 1312 4901 1340
rect 4943 1312 4988 1340
rect 4856 1300 4862 1312
rect 4982 1300 4988 1312
rect 5040 1300 5046 1352
rect 5537 1343 5595 1349
rect 5537 1309 5549 1343
rect 5583 1340 5595 1343
rect 5626 1340 5632 1352
rect 5583 1312 5632 1340
rect 5583 1309 5595 1312
rect 5537 1303 5595 1309
rect 4341 1275 4399 1281
rect 4341 1272 4353 1275
rect 4264 1244 4353 1272
rect 4157 1235 4215 1241
rect 4341 1241 4353 1244
rect 4387 1241 4399 1275
rect 4341 1235 4399 1241
rect 4172 1204 4200 1235
rect 5552 1204 5580 1303
rect 5626 1300 5632 1312
rect 5684 1300 5690 1352
rect 5813 1343 5871 1349
rect 5813 1309 5825 1343
rect 5859 1340 5871 1343
rect 6733 1343 6791 1349
rect 5859 1312 6592 1340
rect 5859 1309 5871 1312
rect 5813 1303 5871 1309
rect 6564 1213 6592 1312
rect 6733 1309 6745 1343
rect 6779 1340 6791 1343
rect 7098 1340 7104 1352
rect 6779 1312 7104 1340
rect 6779 1309 6791 1312
rect 6733 1303 6791 1309
rect 7098 1300 7104 1312
rect 7156 1300 7162 1352
rect 4172 1176 5580 1204
rect 6549 1207 6607 1213
rect 6549 1173 6561 1207
rect 6595 1204 6607 1207
rect 7208 1204 7236 1380
rect 7377 1377 7389 1380
rect 7423 1408 7435 1411
rect 7558 1408 7564 1420
rect 7423 1380 7564 1408
rect 7423 1377 7435 1380
rect 7377 1371 7435 1377
rect 7558 1368 7564 1380
rect 7616 1368 7622 1420
rect 7834 1408 7840 1420
rect 7760 1380 7840 1408
rect 7466 1340 7472 1352
rect 7427 1312 7472 1340
rect 7466 1300 7472 1312
rect 7524 1300 7530 1352
rect 7760 1349 7788 1380
rect 7834 1368 7840 1380
rect 7892 1368 7898 1420
rect 8662 1368 8668 1420
rect 8720 1408 8726 1420
rect 9674 1408 9680 1420
rect 8720 1380 9536 1408
rect 9635 1380 9680 1408
rect 8720 1368 8726 1380
rect 7745 1343 7803 1349
rect 7745 1309 7757 1343
rect 7791 1309 7803 1343
rect 7926 1340 7932 1352
rect 7887 1312 7932 1340
rect 7745 1303 7803 1309
rect 7374 1272 7380 1284
rect 7335 1244 7380 1272
rect 7374 1232 7380 1244
rect 7432 1232 7438 1284
rect 7760 1272 7788 1303
rect 7926 1300 7932 1312
rect 7984 1300 7990 1352
rect 8573 1343 8631 1349
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 9030 1340 9036 1352
rect 8619 1312 9036 1340
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 9030 1300 9036 1312
rect 9088 1300 9094 1352
rect 9214 1340 9220 1352
rect 9175 1312 9220 1340
rect 9214 1300 9220 1312
rect 9272 1300 9278 1352
rect 9398 1340 9404 1352
rect 9359 1312 9404 1340
rect 9398 1300 9404 1312
rect 9456 1300 9462 1352
rect 9508 1349 9536 1380
rect 9674 1368 9680 1380
rect 9732 1368 9738 1420
rect 11238 1408 11244 1420
rect 10980 1380 11244 1408
rect 9493 1343 9551 1349
rect 9493 1309 9505 1343
rect 9539 1309 9551 1343
rect 9493 1303 9551 1309
rect 9950 1300 9956 1352
rect 10008 1340 10014 1352
rect 10045 1343 10103 1349
rect 10045 1340 10057 1343
rect 10008 1312 10057 1340
rect 10008 1300 10014 1312
rect 10045 1309 10057 1312
rect 10091 1309 10103 1343
rect 10980 1340 11008 1380
rect 11238 1368 11244 1380
rect 11296 1408 11302 1420
rect 11296 1380 11744 1408
rect 11296 1368 11302 1380
rect 10045 1303 10103 1309
rect 10888 1312 11008 1340
rect 10888 1272 10916 1312
rect 11054 1300 11060 1352
rect 11112 1340 11118 1352
rect 11514 1340 11520 1352
rect 11112 1312 11520 1340
rect 11112 1300 11118 1312
rect 11514 1300 11520 1312
rect 11572 1300 11578 1352
rect 11716 1349 11744 1380
rect 11790 1368 11796 1420
rect 11848 1408 11854 1420
rect 12069 1411 12127 1417
rect 12069 1408 12081 1411
rect 11848 1380 12081 1408
rect 11848 1368 11854 1380
rect 12069 1377 12081 1380
rect 12115 1377 12127 1411
rect 12069 1371 12127 1377
rect 11701 1343 11759 1349
rect 11701 1309 11713 1343
rect 11747 1309 11759 1343
rect 11882 1340 11888 1352
rect 11843 1312 11888 1340
rect 11701 1303 11759 1309
rect 11882 1300 11888 1312
rect 11940 1300 11946 1352
rect 12618 1340 12624 1352
rect 12579 1312 12624 1340
rect 12618 1300 12624 1312
rect 12676 1300 12682 1352
rect 12713 1343 12771 1349
rect 12713 1309 12725 1343
rect 12759 1309 12771 1343
rect 12713 1303 12771 1309
rect 7760 1244 10916 1272
rect 10962 1232 10968 1284
rect 11020 1272 11026 1284
rect 12728 1272 12756 1303
rect 11020 1244 12756 1272
rect 11020 1232 11026 1244
rect 6595 1176 7236 1204
rect 8389 1207 8447 1213
rect 6595 1173 6607 1176
rect 6549 1167 6607 1173
rect 8389 1173 8401 1207
rect 8435 1204 8447 1207
rect 8570 1204 8576 1216
rect 8435 1176 8576 1204
rect 8435 1173 8447 1176
rect 8389 1167 8447 1173
rect 8570 1164 8576 1176
rect 8628 1164 8634 1216
rect 8938 1164 8944 1216
rect 8996 1204 9002 1216
rect 9861 1207 9919 1213
rect 9861 1204 9873 1207
rect 8996 1176 9873 1204
rect 8996 1164 9002 1176
rect 9861 1173 9873 1176
rect 9907 1173 9919 1207
rect 9861 1167 9919 1173
rect 11146 1164 11152 1216
rect 11204 1204 11210 1216
rect 11241 1207 11299 1213
rect 11241 1204 11253 1207
rect 11204 1176 11253 1204
rect 11204 1164 11210 1176
rect 11241 1173 11253 1176
rect 11287 1173 11299 1207
rect 11241 1167 11299 1173
rect 1104 1114 13892 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 13892 1114
rect 1104 1040 13892 1062
<< via1 >>
rect 9312 13880 9364 13932
rect 14372 13880 14424 13932
rect 8760 13812 8812 13864
rect 11520 13812 11572 13864
rect 7012 13744 7064 13796
rect 13360 13744 13412 13796
rect 9036 13676 9088 13728
rect 11612 13676 11664 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 10784 13472 10836 13524
rect 2872 13404 2924 13456
rect 7564 13404 7616 13456
rect 7656 13447 7708 13456
rect 7656 13413 7665 13447
rect 7665 13413 7699 13447
rect 7699 13413 7708 13447
rect 7656 13404 7708 13413
rect 9036 13404 9088 13456
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2044 13243 2096 13252
rect 1400 13175 1452 13184
rect 1400 13141 1409 13175
rect 1409 13141 1443 13175
rect 1443 13141 1452 13175
rect 2044 13209 2053 13243
rect 2053 13209 2087 13243
rect 2087 13209 2096 13243
rect 3516 13268 3568 13320
rect 4160 13268 4212 13320
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 5080 13311 5132 13320
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 6184 13268 6236 13320
rect 2688 13243 2740 13252
rect 2044 13200 2096 13209
rect 2688 13209 2697 13243
rect 2697 13209 2731 13243
rect 2731 13209 2740 13243
rect 2688 13200 2740 13209
rect 2780 13243 2832 13252
rect 2780 13209 2789 13243
rect 2789 13209 2823 13243
rect 2823 13209 2832 13243
rect 2780 13200 2832 13209
rect 3056 13200 3108 13252
rect 3884 13200 3936 13252
rect 4804 13200 4856 13252
rect 5632 13243 5684 13252
rect 5632 13209 5641 13243
rect 5641 13209 5675 13243
rect 5675 13209 5684 13243
rect 5632 13200 5684 13209
rect 1400 13132 1452 13141
rect 3148 13132 3200 13184
rect 4988 13132 5040 13184
rect 5448 13132 5500 13184
rect 9312 13336 9364 13388
rect 11152 13336 11204 13388
rect 11612 13336 11664 13388
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 7380 13268 7432 13320
rect 7564 13268 7616 13320
rect 8116 13268 8168 13320
rect 8760 13311 8812 13320
rect 7288 13243 7340 13252
rect 7012 13132 7064 13184
rect 7288 13209 7297 13243
rect 7297 13209 7331 13243
rect 7331 13209 7340 13243
rect 7288 13200 7340 13209
rect 7932 13243 7984 13252
rect 7932 13209 7941 13243
rect 7941 13209 7975 13243
rect 7975 13209 7984 13243
rect 7932 13200 7984 13209
rect 8024 13243 8076 13252
rect 8024 13209 8033 13243
rect 8033 13209 8067 13243
rect 8067 13209 8076 13243
rect 8024 13200 8076 13209
rect 7564 13132 7616 13184
rect 8760 13277 8769 13311
rect 8769 13277 8803 13311
rect 8803 13277 8812 13311
rect 8760 13268 8812 13277
rect 9588 13311 9640 13320
rect 9588 13277 9597 13311
rect 9597 13277 9631 13311
rect 9631 13277 9640 13311
rect 9588 13268 9640 13277
rect 10232 13268 10284 13320
rect 10416 13268 10468 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11060 13268 11112 13320
rect 10324 13243 10376 13252
rect 8576 13132 8628 13184
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 10324 13209 10333 13243
rect 10333 13209 10367 13243
rect 10367 13209 10376 13243
rect 10324 13200 10376 13209
rect 10692 13132 10744 13184
rect 10784 13132 10836 13184
rect 11244 13200 11296 13252
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12808 13311 12860 13320
rect 12164 13268 12216 13277
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 12900 13268 12952 13320
rect 11520 13200 11572 13252
rect 12624 13243 12676 13252
rect 12624 13209 12633 13243
rect 12633 13209 12667 13243
rect 12667 13209 12676 13243
rect 12624 13200 12676 13209
rect 13268 13243 13320 13252
rect 13268 13209 13277 13243
rect 13277 13209 13311 13243
rect 13311 13209 13320 13243
rect 13268 13200 13320 13209
rect 13176 13132 13228 13184
rect 13728 13132 13780 13184
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 2780 12928 2832 12980
rect 7656 12928 7708 12980
rect 9496 12928 9548 12980
rect 9588 12928 9640 12980
rect 1952 12860 2004 12912
rect 5264 12860 5316 12912
rect 6184 12903 6236 12912
rect 6184 12869 6193 12903
rect 6193 12869 6227 12903
rect 6227 12869 6236 12903
rect 6184 12860 6236 12869
rect 7012 12860 7064 12912
rect 8024 12860 8076 12912
rect 10048 12903 10100 12912
rect 2596 12835 2648 12844
rect 2596 12801 2605 12835
rect 2605 12801 2639 12835
rect 2639 12801 2648 12835
rect 2596 12792 2648 12801
rect 3056 12792 3108 12844
rect 3424 12792 3476 12844
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 5080 12792 5132 12844
rect 5448 12792 5500 12844
rect 6368 12835 6420 12844
rect 6368 12801 6377 12835
rect 6377 12801 6411 12835
rect 6411 12801 6420 12835
rect 6368 12792 6420 12801
rect 7196 12792 7248 12844
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 10048 12869 10057 12903
rect 10057 12869 10091 12903
rect 10091 12869 10100 12903
rect 10048 12860 10100 12869
rect 10324 12860 10376 12912
rect 10784 12928 10836 12980
rect 10968 12928 11020 12980
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 10692 12860 10744 12912
rect 11888 12860 11940 12912
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 2228 12699 2280 12708
rect 2228 12665 2237 12699
rect 2237 12665 2271 12699
rect 2271 12665 2280 12699
rect 2228 12656 2280 12665
rect 3516 12656 3568 12708
rect 3884 12656 3936 12708
rect 7656 12699 7708 12708
rect 7656 12665 7665 12699
rect 7665 12665 7699 12699
rect 7699 12665 7708 12699
rect 7656 12656 7708 12665
rect 5356 12588 5408 12640
rect 9496 12724 9548 12776
rect 10232 12792 10284 12844
rect 10784 12792 10836 12844
rect 9312 12656 9364 12708
rect 12164 12792 12216 12844
rect 12624 12860 12676 12912
rect 9680 12588 9732 12640
rect 9956 12588 10008 12640
rect 10140 12588 10192 12640
rect 12900 12588 12952 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 4160 12384 4212 12436
rect 4988 12384 5040 12436
rect 5632 12384 5684 12436
rect 2688 12316 2740 12368
rect 3424 12359 3476 12368
rect 2044 12180 2096 12232
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3424 12325 3433 12359
rect 3433 12325 3467 12359
rect 3467 12325 3476 12359
rect 3424 12316 3476 12325
rect 4896 12316 4948 12368
rect 7656 12316 7708 12368
rect 8852 12384 8904 12436
rect 10692 12384 10744 12436
rect 4988 12248 5040 12300
rect 6552 12248 6604 12300
rect 7288 12248 7340 12300
rect 7840 12248 7892 12300
rect 8576 12291 8628 12300
rect 4804 12223 4856 12232
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 5540 12180 5592 12232
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 7196 12180 7248 12232
rect 7564 12180 7616 12232
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 8944 12248 8996 12300
rect 9772 12316 9824 12368
rect 10048 12316 10100 12368
rect 10324 12316 10376 12368
rect 11336 12316 11388 12368
rect 9220 12223 9272 12232
rect 5080 12155 5132 12164
rect 5080 12121 5089 12155
rect 5089 12121 5123 12155
rect 5123 12121 5132 12155
rect 5080 12112 5132 12121
rect 3332 12044 3384 12096
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 3608 12044 3660 12053
rect 4988 12044 5040 12096
rect 5724 12112 5776 12164
rect 5908 12155 5960 12164
rect 5908 12121 5917 12155
rect 5917 12121 5951 12155
rect 5951 12121 5960 12155
rect 5908 12112 5960 12121
rect 6092 12155 6144 12164
rect 6092 12121 6101 12155
rect 6101 12121 6135 12155
rect 6135 12121 6144 12155
rect 6092 12112 6144 12121
rect 6644 12112 6696 12164
rect 7380 12112 7432 12164
rect 9220 12189 9224 12223
rect 9224 12189 9258 12223
rect 9258 12189 9272 12223
rect 9220 12180 9272 12189
rect 9956 12248 10008 12300
rect 11704 12248 11756 12300
rect 9496 12180 9548 12232
rect 9772 12180 9824 12232
rect 10692 12180 10744 12232
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 11244 12180 11296 12232
rect 11520 12180 11572 12232
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 6184 12044 6236 12096
rect 7656 12044 7708 12096
rect 8024 12044 8076 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 11060 12112 11112 12164
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 12348 12155 12400 12164
rect 12348 12121 12357 12155
rect 12357 12121 12391 12155
rect 12391 12121 12400 12155
rect 12348 12112 12400 12121
rect 13452 12155 13504 12164
rect 13452 12121 13461 12155
rect 13461 12121 13495 12155
rect 13495 12121 13504 12155
rect 13452 12112 13504 12121
rect 12072 12044 12124 12096
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 2228 11815 2280 11824
rect 2228 11781 2237 11815
rect 2237 11781 2271 11815
rect 2271 11781 2280 11815
rect 2228 11772 2280 11781
rect 2596 11815 2648 11824
rect 2596 11781 2605 11815
rect 2605 11781 2639 11815
rect 2639 11781 2648 11815
rect 2596 11772 2648 11781
rect 3608 11772 3660 11824
rect 1768 11704 1820 11756
rect 2688 11704 2740 11756
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 3424 11704 3476 11756
rect 3792 11704 3844 11756
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 4804 11772 4856 11824
rect 3976 11704 4028 11713
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 6184 11840 6236 11892
rect 6276 11840 6328 11892
rect 6552 11840 6604 11892
rect 7840 11840 7892 11892
rect 7932 11840 7984 11892
rect 8024 11840 8076 11892
rect 6092 11772 6144 11824
rect 6368 11772 6420 11824
rect 5264 11747 5316 11756
rect 5264 11713 5268 11747
rect 5268 11713 5302 11747
rect 5302 11713 5316 11747
rect 5264 11704 5316 11713
rect 1400 11611 1452 11620
rect 1400 11577 1409 11611
rect 1409 11577 1443 11611
rect 1443 11577 1452 11611
rect 1400 11568 1452 11577
rect 2872 11636 2924 11688
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 4620 11568 4672 11620
rect 4804 11636 4856 11688
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 6460 11704 6512 11756
rect 6644 11747 6696 11756
rect 6644 11713 6653 11747
rect 6653 11713 6687 11747
rect 6687 11713 6696 11747
rect 8208 11772 8260 11824
rect 6644 11704 6696 11713
rect 5724 11636 5776 11688
rect 6552 11636 6604 11688
rect 6736 11636 6788 11688
rect 7472 11704 7524 11756
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 8760 11840 8812 11892
rect 10508 11840 10560 11892
rect 11428 11840 11480 11892
rect 11520 11840 11572 11892
rect 8852 11772 8904 11824
rect 9128 11772 9180 11824
rect 8484 11747 8536 11756
rect 8484 11713 8493 11747
rect 8493 11713 8527 11747
rect 8527 11713 8536 11747
rect 8484 11704 8536 11713
rect 9404 11747 9456 11756
rect 7840 11636 7892 11688
rect 8852 11636 8904 11688
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 10232 11815 10284 11824
rect 10232 11781 10241 11815
rect 10241 11781 10275 11815
rect 10275 11781 10284 11815
rect 10232 11772 10284 11781
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 9312 11679 9364 11688
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 10140 11704 10192 11756
rect 11244 11704 11296 11756
rect 11520 11704 11572 11756
rect 11796 11704 11848 11756
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 12808 11704 12860 11756
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 9312 11636 9364 11645
rect 3608 11500 3660 11552
rect 5356 11500 5408 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6000 11500 6052 11552
rect 7564 11543 7616 11552
rect 7564 11509 7573 11543
rect 7573 11509 7607 11543
rect 7607 11509 7616 11543
rect 7564 11500 7616 11509
rect 7932 11500 7984 11552
rect 9036 11500 9088 11552
rect 9496 11500 9548 11552
rect 10600 11636 10652 11688
rect 11152 11636 11204 11688
rect 12164 11636 12216 11688
rect 10508 11568 10560 11620
rect 12348 11568 12400 11620
rect 13268 11611 13320 11620
rect 13268 11577 13277 11611
rect 13277 11577 13311 11611
rect 13311 11577 13320 11611
rect 13268 11568 13320 11577
rect 10876 11500 10928 11552
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 11980 11500 12032 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 5264 11296 5316 11348
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 6920 11296 6972 11348
rect 7564 11296 7616 11348
rect 7932 11296 7984 11348
rect 8668 11296 8720 11348
rect 9036 11296 9088 11348
rect 10968 11296 11020 11348
rect 11520 11339 11572 11348
rect 11520 11305 11529 11339
rect 11529 11305 11563 11339
rect 11563 11305 11572 11339
rect 11520 11296 11572 11305
rect 11888 11296 11940 11348
rect 2688 11228 2740 11280
rect 1400 11160 1452 11212
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 3608 11203 3660 11212
rect 3608 11169 3617 11203
rect 3617 11169 3651 11203
rect 3651 11169 3660 11203
rect 3608 11160 3660 11169
rect 5172 11228 5224 11280
rect 6184 11228 6236 11280
rect 6276 11228 6328 11280
rect 7012 11228 7064 11280
rect 7288 11271 7340 11280
rect 7288 11237 7297 11271
rect 7297 11237 7331 11271
rect 7331 11237 7340 11271
rect 7288 11228 7340 11237
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 4896 11160 4948 11212
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 5356 11135 5408 11144
rect 5356 11101 5370 11135
rect 5370 11101 5404 11135
rect 5404 11101 5408 11135
rect 5908 11135 5960 11144
rect 5356 11092 5408 11101
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6460 11160 6512 11212
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6828 11135 6880 11144
rect 6644 11092 6696 11101
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 7564 11160 7616 11212
rect 9680 11228 9732 11280
rect 10140 11228 10192 11280
rect 10876 11228 10928 11280
rect 8208 11160 8260 11212
rect 9956 11160 10008 11212
rect 3608 11024 3660 11076
rect 3792 11067 3844 11076
rect 3792 11033 3801 11067
rect 3801 11033 3835 11067
rect 3835 11033 3844 11067
rect 3792 11024 3844 11033
rect 5172 11067 5224 11076
rect 5172 11033 5181 11067
rect 5181 11033 5215 11067
rect 5215 11033 5224 11067
rect 5172 11024 5224 11033
rect 5264 11067 5316 11076
rect 5264 11033 5273 11067
rect 5273 11033 5307 11067
rect 5307 11033 5316 11067
rect 5264 11024 5316 11033
rect 1952 10956 2004 11008
rect 3148 10956 3200 11008
rect 5448 10956 5500 11008
rect 6736 11024 6788 11076
rect 7472 11092 7524 11144
rect 7932 11135 7984 11144
rect 7932 11101 7981 11135
rect 7981 11101 7984 11135
rect 7932 11092 7984 11101
rect 9220 11092 9272 11144
rect 10140 11092 10192 11144
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10508 11135 10560 11144
rect 10232 11092 10284 11101
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 6552 10956 6604 11008
rect 6828 10956 6880 11008
rect 7288 11024 7340 11076
rect 7932 10956 7984 11008
rect 8760 11067 8812 11076
rect 8760 11033 8769 11067
rect 8769 11033 8803 11067
rect 8803 11033 8812 11067
rect 8760 11024 8812 11033
rect 8944 11067 8996 11076
rect 8944 11033 8953 11067
rect 8953 11033 8987 11067
rect 8987 11033 8996 11067
rect 8944 11024 8996 11033
rect 9680 11067 9732 11076
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 9680 11033 9689 11067
rect 9689 11033 9723 11067
rect 9723 11033 9732 11067
rect 9680 11024 9732 11033
rect 9864 11067 9916 11076
rect 9864 11033 9873 11067
rect 9873 11033 9907 11067
rect 9907 11033 9916 11067
rect 9864 11024 9916 11033
rect 10048 11067 10100 11076
rect 10048 11033 10057 11067
rect 10057 11033 10091 11067
rect 10091 11033 10100 11067
rect 10048 11024 10100 11033
rect 11060 11135 11112 11144
rect 11060 11101 11083 11135
rect 11083 11101 11112 11135
rect 11060 11092 11112 11101
rect 11980 11228 12032 11280
rect 12072 11160 12124 11212
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12992 11160 13044 11212
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 13268 11092 13320 11144
rect 11796 11067 11848 11076
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 12072 11067 12124 11076
rect 12072 11033 12081 11067
rect 12081 11033 12115 11067
rect 12115 11033 12124 11067
rect 12072 11024 12124 11033
rect 13084 11067 13136 11076
rect 13084 11033 13093 11067
rect 13093 11033 13127 11067
rect 13127 11033 13136 11067
rect 13084 11024 13136 11033
rect 13636 11024 13688 11076
rect 9588 10956 9640 11008
rect 10324 10956 10376 11008
rect 10600 10956 10652 11008
rect 11336 10956 11388 11008
rect 13360 10956 13412 11008
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 3700 10752 3752 10804
rect 2320 10616 2372 10668
rect 2872 10616 2924 10668
rect 3332 10659 3384 10668
rect 3332 10625 3336 10659
rect 3336 10625 3370 10659
rect 3370 10625 3384 10659
rect 3332 10616 3384 10625
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 3608 10616 3660 10668
rect 572 10548 624 10600
rect 2688 10523 2740 10532
rect 2688 10489 2697 10523
rect 2697 10489 2731 10523
rect 2731 10489 2740 10523
rect 2688 10480 2740 10489
rect 5356 10752 5408 10804
rect 6460 10752 6512 10804
rect 4896 10684 4948 10736
rect 5264 10727 5316 10736
rect 5264 10693 5273 10727
rect 5273 10693 5307 10727
rect 5307 10693 5316 10727
rect 5264 10684 5316 10693
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 6092 10616 6144 10668
rect 6276 10616 6328 10668
rect 8116 10752 8168 10804
rect 8484 10752 8536 10804
rect 9496 10684 9548 10736
rect 5264 10480 5316 10532
rect 6552 10548 6604 10600
rect 7380 10548 7432 10600
rect 7932 10659 7984 10668
rect 7932 10625 7941 10659
rect 7941 10625 7975 10659
rect 7975 10625 7984 10659
rect 7932 10616 7984 10625
rect 6920 10480 6972 10532
rect 7104 10480 7156 10532
rect 8024 10548 8076 10600
rect 8116 10523 8168 10532
rect 3056 10412 3108 10464
rect 3516 10412 3568 10464
rect 6460 10412 6512 10464
rect 6736 10412 6788 10464
rect 7472 10412 7524 10464
rect 8116 10489 8125 10523
rect 8125 10489 8159 10523
rect 8159 10489 8168 10523
rect 8392 10548 8444 10600
rect 9036 10616 9088 10668
rect 9588 10616 9640 10668
rect 10048 10752 10100 10804
rect 10692 10752 10744 10804
rect 10968 10727 11020 10736
rect 10968 10693 10977 10727
rect 10977 10693 11011 10727
rect 11011 10693 11020 10727
rect 10968 10684 11020 10693
rect 11152 10752 11204 10804
rect 11336 10752 11388 10804
rect 11428 10752 11480 10804
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 8116 10480 8168 10489
rect 8300 10412 8352 10464
rect 8392 10412 8444 10464
rect 9128 10412 9180 10464
rect 9956 10548 10008 10600
rect 10600 10616 10652 10668
rect 10692 10659 10744 10668
rect 10692 10625 10741 10659
rect 10741 10625 10744 10659
rect 10692 10616 10744 10625
rect 12164 10684 12216 10736
rect 11980 10659 12032 10668
rect 11980 10625 11989 10659
rect 11989 10625 12023 10659
rect 12023 10625 12032 10659
rect 11980 10616 12032 10625
rect 12624 10616 12676 10668
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 12072 10548 12124 10600
rect 10600 10523 10652 10532
rect 10600 10489 10609 10523
rect 10609 10489 10643 10523
rect 10643 10489 10652 10523
rect 10600 10480 10652 10489
rect 11060 10480 11112 10532
rect 11336 10480 11388 10532
rect 13084 10480 13136 10532
rect 9680 10412 9732 10464
rect 11152 10412 11204 10464
rect 11428 10412 11480 10464
rect 11796 10412 11848 10464
rect 13176 10412 13228 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 6276 10208 6328 10260
rect 6460 10251 6512 10260
rect 6460 10217 6469 10251
rect 6469 10217 6503 10251
rect 6503 10217 6512 10251
rect 6460 10208 6512 10217
rect 8116 10208 8168 10260
rect 8300 10208 8352 10260
rect 5080 10183 5132 10192
rect 5080 10149 5089 10183
rect 5089 10149 5123 10183
rect 5123 10149 5132 10183
rect 5080 10140 5132 10149
rect 5724 10183 5776 10192
rect 5724 10149 5733 10183
rect 5733 10149 5767 10183
rect 5767 10149 5776 10183
rect 5724 10140 5776 10149
rect 6184 10140 6236 10192
rect 7564 10140 7616 10192
rect 8484 10140 8536 10192
rect 8576 10140 8628 10192
rect 9128 10208 9180 10260
rect 9680 10208 9732 10260
rect 10048 10208 10100 10260
rect 2688 10047 2740 10056
rect 1952 9979 2004 9988
rect 1952 9945 1961 9979
rect 1961 9945 1995 9979
rect 1995 9945 2004 9979
rect 1952 9936 2004 9945
rect 2688 10013 2697 10047
rect 2697 10013 2731 10047
rect 2731 10013 2740 10047
rect 2688 10004 2740 10013
rect 3240 10004 3292 10056
rect 5172 10072 5224 10124
rect 3976 10004 4028 10056
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6368 10072 6420 10124
rect 6276 10004 6328 10056
rect 7288 10072 7340 10124
rect 6828 10004 6880 10056
rect 2872 9936 2924 9988
rect 6092 9979 6144 9988
rect 6092 9945 6101 9979
rect 6101 9945 6135 9979
rect 6135 9945 6144 9979
rect 6092 9936 6144 9945
rect 6552 9936 6604 9988
rect 6644 9979 6696 9988
rect 6644 9945 6653 9979
rect 6653 9945 6687 9979
rect 6687 9945 6696 9979
rect 6644 9936 6696 9945
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 2964 9911 3016 9920
rect 2964 9877 2973 9911
rect 2973 9877 3007 9911
rect 3007 9877 3016 9911
rect 2964 9868 3016 9877
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 3240 9868 3292 9920
rect 5448 9911 5500 9920
rect 5448 9877 5457 9911
rect 5457 9877 5491 9911
rect 5491 9877 5500 9911
rect 5448 9868 5500 9877
rect 5724 9868 5776 9920
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 7932 10004 7984 10056
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 8484 10047 8536 10090
rect 8484 10038 8493 10047
rect 8493 10038 8527 10047
rect 8527 10038 8536 10047
rect 9864 10072 9916 10124
rect 10048 10072 10100 10124
rect 10140 10072 10192 10124
rect 7012 9936 7064 9988
rect 7288 9936 7340 9988
rect 8116 9936 8168 9988
rect 9588 10004 9640 10056
rect 9036 9936 9088 9988
rect 7196 9868 7248 9920
rect 7564 9911 7616 9920
rect 7564 9877 7573 9911
rect 7573 9877 7607 9911
rect 7607 9877 7616 9911
rect 7564 9868 7616 9877
rect 9128 9868 9180 9920
rect 9312 9868 9364 9920
rect 10048 9868 10100 9920
rect 10416 10004 10468 10056
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 10968 10072 11020 10124
rect 11980 10072 12032 10124
rect 11612 10004 11664 10056
rect 13176 10208 13228 10260
rect 10600 9979 10652 9988
rect 10600 9945 10609 9979
rect 10609 9945 10643 9979
rect 10643 9945 10652 9979
rect 10600 9936 10652 9945
rect 10784 9936 10836 9988
rect 11428 9936 11480 9988
rect 12716 10004 12768 10056
rect 12900 9936 12952 9988
rect 10416 9868 10468 9920
rect 10692 9868 10744 9920
rect 12440 9868 12492 9920
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 3424 9664 3476 9716
rect 4896 9707 4948 9716
rect 4896 9673 4905 9707
rect 4905 9673 4939 9707
rect 4939 9673 4948 9707
rect 4896 9664 4948 9673
rect 6552 9664 6604 9716
rect 7840 9664 7892 9716
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 1676 9596 1728 9648
rect 1952 9639 2004 9648
rect 1952 9605 1961 9639
rect 1961 9605 1995 9639
rect 1995 9605 2004 9639
rect 1952 9596 2004 9605
rect 2872 9596 2924 9648
rect 5080 9596 5132 9648
rect 5448 9596 5500 9648
rect 6368 9639 6420 9648
rect 6368 9605 6377 9639
rect 6377 9605 6411 9639
rect 6411 9605 6420 9639
rect 6368 9596 6420 9605
rect 6644 9596 6696 9648
rect 7288 9639 7340 9648
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 3424 9528 3476 9580
rect 3976 9571 4028 9580
rect 3976 9537 3985 9571
rect 3985 9537 4019 9571
rect 4019 9537 4028 9571
rect 3976 9528 4028 9537
rect 4896 9528 4948 9580
rect 6000 9528 6052 9580
rect 6460 9528 6512 9580
rect 7288 9605 7297 9639
rect 7297 9605 7331 9639
rect 7331 9605 7340 9639
rect 7288 9596 7340 9605
rect 2688 9460 2740 9512
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 3332 9392 3384 9444
rect 5264 9435 5316 9444
rect 5264 9401 5273 9435
rect 5273 9401 5307 9435
rect 5307 9401 5316 9435
rect 5264 9392 5316 9401
rect 6092 9460 6144 9512
rect 7104 9528 7156 9580
rect 6736 9392 6788 9444
rect 6828 9392 6880 9444
rect 8300 9639 8352 9648
rect 8300 9605 8309 9639
rect 8309 9605 8343 9639
rect 8343 9605 8352 9639
rect 8944 9664 8996 9716
rect 9956 9664 10008 9716
rect 10232 9664 10284 9716
rect 8300 9596 8352 9605
rect 8392 9571 8444 9580
rect 8392 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8444 9571
rect 8392 9528 8444 9537
rect 8760 9528 8812 9580
rect 8300 9460 8352 9512
rect 9128 9528 9180 9580
rect 9588 9571 9640 9580
rect 9588 9537 9597 9571
rect 9597 9537 9631 9571
rect 9631 9537 9640 9571
rect 9588 9528 9640 9537
rect 9772 9528 9824 9580
rect 9956 9571 10008 9580
rect 9956 9537 9975 9571
rect 9975 9537 10008 9571
rect 9956 9528 10008 9537
rect 10324 9596 10376 9648
rect 11060 9596 11112 9648
rect 11244 9596 11296 9648
rect 11612 9596 11664 9648
rect 10508 9528 10560 9580
rect 9680 9460 9732 9512
rect 11428 9528 11480 9580
rect 11704 9528 11756 9580
rect 1860 9324 1912 9376
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 8668 9392 8720 9444
rect 8852 9392 8904 9444
rect 8944 9324 8996 9376
rect 12808 9460 12860 9512
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 11152 9392 11204 9444
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 10784 9324 10836 9376
rect 12624 9324 12676 9376
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 1768 9120 1820 9172
rect 2688 9120 2740 9172
rect 3608 9163 3660 9172
rect 3608 9129 3617 9163
rect 3617 9129 3651 9163
rect 3651 9129 3660 9163
rect 3608 9120 3660 9129
rect 6184 9163 6236 9172
rect 6184 9129 6193 9163
rect 6193 9129 6227 9163
rect 6227 9129 6236 9163
rect 6184 9120 6236 9129
rect 6460 9163 6512 9172
rect 6460 9129 6469 9163
rect 6469 9129 6503 9163
rect 6503 9129 6512 9163
rect 6460 9120 6512 9129
rect 7104 9120 7156 9172
rect 7656 9120 7708 9172
rect 7840 9120 7892 9172
rect 8668 9120 8720 9172
rect 8760 9120 8812 9172
rect 10048 9120 10100 9172
rect 12808 9163 12860 9172
rect 6920 9052 6972 9104
rect 7196 9052 7248 9104
rect 7564 9052 7616 9104
rect 2780 8984 2832 9036
rect 2964 8984 3016 9036
rect 3976 8984 4028 9036
rect 3332 8959 3384 8968
rect 3332 8925 3341 8959
rect 3341 8925 3375 8959
rect 3375 8925 3384 8959
rect 3332 8916 3384 8925
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 5632 8916 5684 8968
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6828 8916 6880 8968
rect 7472 8959 7524 8968
rect 3056 8848 3108 8900
rect 3424 8891 3476 8900
rect 3424 8857 3433 8891
rect 3433 8857 3467 8891
rect 3467 8857 3476 8891
rect 3424 8848 3476 8857
rect 4896 8891 4948 8900
rect 4896 8857 4905 8891
rect 4905 8857 4939 8891
rect 4939 8857 4948 8891
rect 4896 8848 4948 8857
rect 4988 8891 5040 8900
rect 4988 8857 4997 8891
rect 4997 8857 5031 8891
rect 5031 8857 5040 8891
rect 5264 8891 5316 8900
rect 4988 8848 5040 8857
rect 5264 8857 5273 8891
rect 5273 8857 5307 8891
rect 5307 8857 5316 8891
rect 5264 8848 5316 8857
rect 6368 8848 6420 8900
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 7840 8916 7892 8968
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 7196 8891 7248 8900
rect 7196 8857 7205 8891
rect 7205 8857 7239 8891
rect 7239 8857 7248 8891
rect 7196 8848 7248 8857
rect 8760 8984 8812 9036
rect 9496 9052 9548 9104
rect 9772 9052 9824 9104
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 10692 9095 10744 9104
rect 10692 9061 10701 9095
rect 10701 9061 10735 9095
rect 10735 9061 10744 9095
rect 10692 9052 10744 9061
rect 11152 9095 11204 9104
rect 11152 9061 11161 9095
rect 11161 9061 11195 9095
rect 11195 9061 11204 9095
rect 11152 9052 11204 9061
rect 9036 8916 9088 8968
rect 9680 8984 9732 9036
rect 11244 8984 11296 9036
rect 9220 8925 9230 8946
rect 9230 8925 9264 8946
rect 9264 8925 9272 8946
rect 9220 8894 9272 8925
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 10140 8916 10192 8968
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 11060 8916 11112 8968
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2780 8780 2832 8832
rect 6644 8780 6696 8832
rect 8852 8780 8904 8832
rect 9956 8848 10008 8900
rect 12072 8848 12124 8900
rect 12532 8848 12584 8900
rect 13544 8848 13596 8900
rect 10048 8780 10100 8832
rect 10416 8780 10468 8832
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 4988 8576 5040 8628
rect 3332 8508 3384 8560
rect 7840 8576 7892 8628
rect 8576 8576 8628 8628
rect 9036 8619 9088 8628
rect 9036 8585 9045 8619
rect 9045 8585 9079 8619
rect 9079 8585 9088 8619
rect 9036 8576 9088 8585
rect 9496 8576 9548 8628
rect 10232 8576 10284 8628
rect 10968 8576 11020 8628
rect 7288 8508 7340 8560
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2688 8372 2740 8424
rect 3976 8440 4028 8492
rect 4436 8440 4488 8492
rect 5632 8440 5684 8492
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 6828 8440 6880 8492
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 8116 8508 8168 8560
rect 9404 8508 9456 8560
rect 8576 8483 8628 8492
rect 8576 8449 8585 8483
rect 8585 8449 8619 8483
rect 8619 8449 8628 8483
rect 8576 8440 8628 8449
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9128 8440 9180 8492
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9496 8483 9548 8492
rect 9312 8440 9364 8449
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9864 8508 9916 8560
rect 9680 8440 9732 8492
rect 10692 8483 10744 8492
rect 10692 8449 10695 8483
rect 10695 8449 10729 8483
rect 10729 8449 10744 8483
rect 10968 8483 11020 8492
rect 10692 8440 10744 8449
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 6092 8372 6144 8424
rect 9772 8372 9824 8424
rect 10048 8415 10100 8424
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 10324 8372 10376 8424
rect 4896 8304 4948 8356
rect 6920 8347 6972 8356
rect 6920 8313 6929 8347
rect 6929 8313 6963 8347
rect 6963 8313 6972 8347
rect 6920 8304 6972 8313
rect 8024 8304 8076 8356
rect 9220 8304 9272 8356
rect 12716 8576 12768 8628
rect 13452 8576 13504 8628
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 3240 8236 3292 8288
rect 6368 8236 6420 8288
rect 7472 8236 7524 8288
rect 8760 8236 8812 8288
rect 8944 8236 8996 8288
rect 9312 8236 9364 8288
rect 11704 8347 11756 8356
rect 11704 8313 11713 8347
rect 11713 8313 11747 8347
rect 11747 8313 11756 8347
rect 12900 8508 12952 8560
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12808 8440 12860 8492
rect 12900 8372 12952 8424
rect 13176 8372 13228 8424
rect 13452 8440 13504 8492
rect 11704 8304 11756 8313
rect 12072 8304 12124 8356
rect 12164 8304 12216 8356
rect 12808 8304 12860 8356
rect 10232 8236 10284 8288
rect 10508 8279 10560 8288
rect 10508 8245 10517 8279
rect 10517 8245 10551 8279
rect 10551 8245 10560 8279
rect 10508 8236 10560 8245
rect 11060 8236 11112 8288
rect 13728 8236 13780 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 3700 8032 3752 8084
rect 4620 8032 4672 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 8668 8032 8720 8084
rect 9404 8075 9456 8084
rect 9404 8041 9413 8075
rect 9413 8041 9447 8075
rect 9447 8041 9456 8075
rect 9404 8032 9456 8041
rect 10784 8032 10836 8084
rect 1676 8007 1728 8016
rect 1676 7973 1685 8007
rect 1685 7973 1719 8007
rect 1719 7973 1728 8007
rect 1676 7964 1728 7973
rect 3884 7964 3936 8016
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 1768 7828 1820 7880
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 3976 7896 4028 7948
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 1952 7692 2004 7744
rect 2780 7803 2832 7812
rect 2780 7769 2789 7803
rect 2789 7769 2823 7803
rect 2823 7769 2832 7803
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3884 7871 3936 7880
rect 3240 7828 3292 7837
rect 2780 7760 2832 7769
rect 3056 7760 3108 7812
rect 3884 7837 3893 7871
rect 3893 7837 3927 7871
rect 3927 7837 3936 7871
rect 3884 7828 3936 7837
rect 4712 7896 4764 7948
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 7840 7964 7892 8016
rect 9036 8007 9088 8016
rect 7656 7896 7708 7948
rect 9036 7973 9045 8007
rect 9045 7973 9079 8007
rect 9079 7973 9088 8007
rect 9036 7964 9088 7973
rect 9220 7964 9272 8016
rect 11244 8007 11296 8016
rect 11244 7973 11253 8007
rect 11253 7973 11287 8007
rect 11287 7973 11296 8007
rect 11244 7964 11296 7973
rect 11980 7964 12032 8016
rect 13084 7964 13136 8016
rect 4804 7828 4856 7837
rect 5448 7871 5500 7880
rect 3792 7760 3844 7812
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 6184 7828 6236 7880
rect 7472 7828 7524 7880
rect 5356 7760 5408 7812
rect 5816 7760 5868 7812
rect 6828 7760 6880 7812
rect 7932 7803 7984 7812
rect 7932 7769 7941 7803
rect 7941 7769 7975 7803
rect 7975 7769 7984 7803
rect 9312 7828 9364 7880
rect 10048 7896 10100 7948
rect 9680 7828 9732 7880
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 10968 7896 11020 7948
rect 11336 7896 11388 7948
rect 9864 7828 9916 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 11060 7828 11112 7880
rect 11520 7828 11572 7880
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 7932 7760 7984 7769
rect 10600 7760 10652 7812
rect 11888 7760 11940 7812
rect 12072 7803 12124 7812
rect 12072 7769 12081 7803
rect 12081 7769 12115 7803
rect 12115 7769 12124 7803
rect 12072 7760 12124 7769
rect 2596 7735 2648 7744
rect 2596 7701 2605 7735
rect 2605 7701 2639 7735
rect 2639 7701 2648 7735
rect 2596 7692 2648 7701
rect 4068 7735 4120 7744
rect 4068 7701 4077 7735
rect 4077 7701 4111 7735
rect 4111 7701 4120 7735
rect 4068 7692 4120 7701
rect 5540 7692 5592 7744
rect 5908 7735 5960 7744
rect 5908 7701 5917 7735
rect 5917 7701 5951 7735
rect 5951 7701 5960 7735
rect 5908 7692 5960 7701
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 7472 7692 7524 7744
rect 8116 7692 8168 7744
rect 8760 7692 8812 7744
rect 9128 7692 9180 7744
rect 10232 7692 10284 7744
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 11152 7692 11204 7744
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 12624 7692 12676 7744
rect 13360 7692 13412 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 1492 7488 1544 7540
rect 2136 7488 2188 7540
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 3884 7488 3936 7540
rect 7288 7488 7340 7540
rect 6920 7420 6972 7472
rect 8116 7488 8168 7540
rect 8208 7488 8260 7540
rect 9220 7531 9272 7540
rect 9220 7497 9229 7531
rect 9229 7497 9263 7531
rect 9263 7497 9272 7531
rect 9220 7488 9272 7497
rect 4068 7352 4120 7404
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 3516 7284 3568 7336
rect 3976 7284 4028 7336
rect 5356 7352 5408 7404
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 8760 7395 8812 7404
rect 8760 7361 8783 7395
rect 8783 7361 8812 7395
rect 5264 7284 5316 7336
rect 8300 7284 8352 7336
rect 8760 7352 8812 7361
rect 9128 7352 9180 7404
rect 9404 7352 9456 7404
rect 10416 7488 10468 7540
rect 10508 7488 10560 7540
rect 10232 7420 10284 7472
rect 10140 7352 10192 7404
rect 9864 7284 9916 7336
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 11704 7488 11756 7540
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 12164 7395 12216 7404
rect 11888 7352 11940 7361
rect 12164 7361 12173 7395
rect 12173 7361 12207 7395
rect 12207 7361 12216 7395
rect 12164 7352 12216 7361
rect 11704 7284 11756 7336
rect 12072 7327 12124 7336
rect 12072 7293 12081 7327
rect 12081 7293 12115 7327
rect 12115 7293 12124 7327
rect 12072 7284 12124 7293
rect 12532 7284 12584 7336
rect 12992 7327 13044 7336
rect 12992 7293 13001 7327
rect 13001 7293 13035 7327
rect 13035 7293 13044 7327
rect 12992 7284 13044 7293
rect 4804 7216 4856 7268
rect 6828 7216 6880 7268
rect 10416 7259 10468 7268
rect 10416 7225 10429 7259
rect 10429 7225 10463 7259
rect 10463 7225 10468 7259
rect 10416 7216 10468 7225
rect 2964 7148 3016 7200
rect 4620 7148 4672 7200
rect 12808 7216 12860 7268
rect 13176 7216 13228 7268
rect 11612 7191 11664 7200
rect 11612 7157 11621 7191
rect 11621 7157 11655 7191
rect 11655 7157 11664 7191
rect 11612 7148 11664 7157
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 3516 6987 3568 6996
rect 3516 6953 3525 6987
rect 3525 6953 3559 6987
rect 3559 6953 3568 6987
rect 3516 6944 3568 6953
rect 5540 6944 5592 6996
rect 6828 6944 6880 6996
rect 9956 6944 10008 6996
rect 10416 6944 10468 6996
rect 10968 6944 11020 6996
rect 11612 6944 11664 6996
rect 12624 6987 12676 6996
rect 12624 6953 12633 6987
rect 12633 6953 12667 6987
rect 12667 6953 12676 6987
rect 12624 6944 12676 6953
rect 11060 6876 11112 6928
rect 2964 6808 3016 6860
rect 5264 6808 5316 6860
rect 7932 6808 7984 6860
rect 3424 6740 3476 6792
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 6368 6783 6420 6792
rect 2688 6672 2740 6724
rect 2964 6715 3016 6724
rect 2964 6681 2973 6715
rect 2973 6681 3007 6715
rect 3007 6681 3016 6715
rect 2964 6672 3016 6681
rect 4252 6715 4304 6724
rect 4252 6681 4261 6715
rect 4261 6681 4295 6715
rect 4295 6681 4304 6715
rect 4252 6672 4304 6681
rect 5632 6604 5684 6656
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 7012 6672 7064 6724
rect 7288 6672 7340 6724
rect 10324 6808 10376 6860
rect 12072 6808 12124 6860
rect 9128 6740 9180 6792
rect 9864 6740 9916 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 12992 6808 13044 6860
rect 13176 6851 13228 6860
rect 13176 6817 13185 6851
rect 13185 6817 13219 6851
rect 13219 6817 13228 6851
rect 13176 6808 13228 6817
rect 12716 6740 12768 6792
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 8300 6672 8352 6724
rect 10416 6672 10468 6724
rect 11060 6672 11112 6724
rect 7104 6604 7156 6656
rect 8116 6604 8168 6656
rect 9312 6604 9364 6656
rect 10324 6647 10376 6656
rect 10324 6613 10333 6647
rect 10333 6613 10367 6647
rect 10367 6613 10376 6647
rect 10324 6604 10376 6613
rect 11796 6604 11848 6656
rect 12164 6604 12216 6656
rect 13360 6672 13412 6724
rect 13084 6647 13136 6656
rect 13084 6613 13093 6647
rect 13093 6613 13127 6647
rect 13127 6613 13136 6647
rect 13268 6647 13320 6656
rect 13084 6604 13136 6613
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 1768 6400 1820 6452
rect 1492 6332 1544 6384
rect 2964 6400 3016 6452
rect 4252 6400 4304 6452
rect 6920 6400 6972 6452
rect 7288 6443 7340 6452
rect 7288 6409 7297 6443
rect 7297 6409 7331 6443
rect 7331 6409 7340 6443
rect 7288 6400 7340 6409
rect 9128 6400 9180 6452
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 1768 6264 1820 6316
rect 2228 6264 2280 6316
rect 2872 6264 2924 6316
rect 3700 6264 3752 6316
rect 4620 6332 4672 6384
rect 1860 6128 1912 6180
rect 3056 6128 3108 6180
rect 3424 6171 3476 6180
rect 3424 6137 3433 6171
rect 3433 6137 3467 6171
rect 3467 6137 3476 6171
rect 3424 6128 3476 6137
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 4068 6128 4120 6180
rect 1492 6060 1544 6112
rect 3700 6060 3752 6112
rect 5448 6264 5500 6316
rect 6184 6264 6236 6316
rect 6368 6264 6420 6316
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 7104 6264 7156 6316
rect 7748 6264 7800 6316
rect 9128 6264 9180 6316
rect 10324 6400 10376 6452
rect 10784 6400 10836 6452
rect 9864 6375 9916 6384
rect 9864 6341 9873 6375
rect 9873 6341 9907 6375
rect 9907 6341 9916 6375
rect 9864 6332 9916 6341
rect 10416 6332 10468 6384
rect 9680 6264 9732 6316
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10192 6307
rect 10140 6264 10192 6273
rect 7288 6196 7340 6248
rect 8024 6196 8076 6248
rect 8116 6196 8168 6248
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 10508 6239 10560 6248
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10968 6332 11020 6384
rect 11888 6400 11940 6452
rect 12900 6400 12952 6452
rect 13728 6400 13780 6452
rect 11428 6332 11480 6384
rect 11520 6307 11572 6316
rect 11520 6273 11529 6307
rect 11529 6273 11563 6307
rect 11563 6273 11572 6307
rect 11520 6264 11572 6273
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 13636 6332 13688 6384
rect 11888 6264 11940 6316
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 13176 6264 13228 6316
rect 10508 6196 10560 6205
rect 4712 6060 4764 6112
rect 4896 6060 4948 6112
rect 5632 6128 5684 6180
rect 6920 6128 6972 6180
rect 7012 6128 7064 6180
rect 9864 6128 9916 6180
rect 10600 6128 10652 6180
rect 12900 6171 12952 6180
rect 12900 6137 12909 6171
rect 12909 6137 12943 6171
rect 12943 6137 12952 6171
rect 12900 6128 12952 6137
rect 5356 6060 5408 6112
rect 7196 6060 7248 6112
rect 9772 6060 9824 6112
rect 10048 6060 10100 6112
rect 10508 6060 10560 6112
rect 12624 6103 12676 6112
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 12624 6060 12676 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 2872 5856 2924 5908
rect 4160 5856 4212 5908
rect 1584 5788 1636 5840
rect 2320 5788 2372 5840
rect 1492 5695 1544 5704
rect 1492 5661 1501 5695
rect 1501 5661 1535 5695
rect 1535 5661 1544 5695
rect 1492 5652 1544 5661
rect 1860 5652 1912 5704
rect 1676 5584 1728 5636
rect 2320 5695 2372 5704
rect 2320 5661 2330 5695
rect 2330 5661 2364 5695
rect 2364 5661 2372 5695
rect 2688 5695 2740 5704
rect 2320 5652 2372 5661
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 4988 5856 5040 5908
rect 4620 5720 4672 5772
rect 6092 5856 6144 5908
rect 6920 5720 6972 5772
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4712 5695 4764 5704
rect 4528 5652 4580 5661
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4896 5695 4948 5704
rect 4896 5661 4905 5695
rect 4905 5661 4939 5695
rect 4939 5661 4948 5695
rect 4896 5652 4948 5661
rect 5448 5695 5500 5704
rect 2872 5584 2924 5636
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 7196 5652 7248 5704
rect 9680 5856 9732 5908
rect 12532 5856 12584 5908
rect 12716 5856 12768 5908
rect 1952 5516 2004 5568
rect 2228 5516 2280 5568
rect 3056 5516 3108 5568
rect 3884 5559 3936 5568
rect 3884 5525 3893 5559
rect 3893 5525 3927 5559
rect 3927 5525 3936 5559
rect 3884 5516 3936 5525
rect 4160 5516 4212 5568
rect 6460 5584 6512 5636
rect 7104 5584 7156 5636
rect 8852 5652 8904 5704
rect 10324 5720 10376 5772
rect 9956 5652 10008 5704
rect 10048 5652 10100 5704
rect 12072 5720 12124 5772
rect 12992 5720 13044 5772
rect 12808 5652 12860 5704
rect 12072 5584 12124 5636
rect 6092 5516 6144 5568
rect 7748 5516 7800 5568
rect 8852 5516 8904 5568
rect 10232 5516 10284 5568
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 12808 5516 12860 5568
rect 13268 5516 13320 5568
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 4160 5312 4212 5364
rect 5448 5312 5500 5364
rect 3884 5287 3936 5296
rect 3884 5253 3893 5287
rect 3893 5253 3927 5287
rect 3927 5253 3936 5287
rect 3884 5244 3936 5253
rect 4804 5244 4856 5296
rect 2412 5219 2464 5228
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 3976 5176 4028 5228
rect 8116 5312 8168 5364
rect 9864 5355 9916 5364
rect 6460 5244 6512 5296
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 7104 5244 7156 5296
rect 7840 5244 7892 5296
rect 5908 5176 5960 5185
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 9864 5321 9873 5355
rect 9873 5321 9907 5355
rect 9907 5321 9916 5355
rect 9864 5312 9916 5321
rect 9956 5244 10008 5296
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 9864 5176 9916 5228
rect 10324 5312 10376 5364
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 10232 5244 10284 5296
rect 11244 5244 11296 5296
rect 11704 5244 11756 5296
rect 11796 5244 11848 5296
rect 2780 5108 2832 5117
rect 3792 5108 3844 5160
rect 1952 5040 2004 5092
rect 2228 5040 2280 5092
rect 3884 4972 3936 5024
rect 4528 5040 4580 5092
rect 10324 5151 10376 5160
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 11520 5176 11572 5228
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 12716 5176 12768 5228
rect 12992 5219 13044 5228
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 12624 5151 12676 5160
rect 9312 5083 9364 5092
rect 9312 5049 9321 5083
rect 9321 5049 9355 5083
rect 9355 5049 9364 5083
rect 9312 5040 9364 5049
rect 9404 5040 9456 5092
rect 10048 5040 10100 5092
rect 4896 4972 4948 5024
rect 9220 4972 9272 5024
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 13084 5108 13136 5160
rect 12716 5083 12768 5092
rect 12716 5049 12725 5083
rect 12725 5049 12759 5083
rect 12759 5049 12768 5083
rect 12716 5040 12768 5049
rect 12532 4972 12584 5024
rect 12624 4972 12676 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 2136 4743 2188 4752
rect 2136 4709 2145 4743
rect 2145 4709 2179 4743
rect 2179 4709 2188 4743
rect 2136 4700 2188 4709
rect 5908 4768 5960 4820
rect 6920 4768 6972 4820
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 3332 4632 3384 4684
rect 3608 4632 3660 4684
rect 1492 4496 1544 4548
rect 2780 4564 2832 4616
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 3056 4607 3108 4616
rect 2872 4564 2924 4573
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3792 4607 3844 4616
rect 3148 4564 3200 4573
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 3976 4564 4028 4616
rect 4712 4632 4764 4684
rect 4896 4632 4948 4684
rect 7104 4700 7156 4752
rect 4896 4539 4948 4548
rect 4896 4505 4905 4539
rect 4905 4505 4939 4539
rect 4939 4505 4948 4539
rect 4896 4496 4948 4505
rect 5724 4539 5776 4548
rect 5724 4505 5733 4539
rect 5733 4505 5767 4539
rect 5767 4505 5776 4539
rect 5724 4496 5776 4505
rect 7288 4632 7340 4684
rect 10324 4768 10376 4820
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 7840 4700 7892 4752
rect 13268 4700 13320 4752
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 7196 4607 7248 4616
rect 6644 4564 6696 4573
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 9128 4632 9180 4684
rect 9220 4607 9272 4616
rect 6000 4539 6052 4548
rect 6000 4505 6009 4539
rect 6009 4505 6043 4539
rect 6043 4505 6052 4539
rect 6000 4496 6052 4505
rect 6184 4539 6236 4548
rect 6184 4505 6193 4539
rect 6193 4505 6227 4539
rect 6227 4505 6236 4539
rect 6184 4496 6236 4505
rect 7104 4496 7156 4548
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 10784 4632 10836 4684
rect 11796 4632 11848 4684
rect 9404 4564 9456 4616
rect 12716 4564 12768 4616
rect 13360 4564 13412 4616
rect 8668 4496 8720 4548
rect 9772 4539 9824 4548
rect 9772 4505 9781 4539
rect 9781 4505 9815 4539
rect 9815 4505 9824 4539
rect 9772 4496 9824 4505
rect 10232 4496 10284 4548
rect 13728 4496 13780 4548
rect 2044 4428 2096 4480
rect 2688 4428 2740 4480
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 4436 4428 4488 4480
rect 4988 4428 5040 4480
rect 7380 4428 7432 4480
rect 9588 4428 9640 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 3148 4224 3200 4276
rect 3884 4224 3936 4276
rect 1492 4199 1544 4208
rect 1492 4165 1501 4199
rect 1501 4165 1535 4199
rect 1535 4165 1544 4199
rect 1492 4156 1544 4165
rect 2872 4156 2924 4208
rect 3608 4156 3660 4208
rect 1768 4088 1820 4140
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 3056 4088 3108 4140
rect 3148 4088 3200 4140
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 3608 3952 3660 4004
rect 4988 4156 5040 4208
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4896 4088 4948 4140
rect 5172 4088 5224 4140
rect 6368 4156 6420 4208
rect 6920 4156 6972 4208
rect 9496 4224 9548 4276
rect 9772 4224 9824 4276
rect 10416 4224 10468 4276
rect 11060 4267 11112 4276
rect 11060 4233 11069 4267
rect 11069 4233 11103 4267
rect 11103 4233 11112 4267
rect 11060 4224 11112 4233
rect 11244 4224 11296 4276
rect 9404 4156 9456 4208
rect 5908 4088 5960 4140
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 8576 4088 8628 4140
rect 11888 4156 11940 4208
rect 5080 4020 5132 4072
rect 5724 4020 5776 4072
rect 6736 4020 6788 4072
rect 7288 4020 7340 4072
rect 5264 3952 5316 4004
rect 6552 3952 6604 4004
rect 9772 4020 9824 4072
rect 10784 4088 10836 4140
rect 11244 4131 11296 4140
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 2964 3884 3016 3893
rect 4620 3884 4672 3936
rect 6644 3884 6696 3936
rect 6828 3884 6880 3936
rect 9220 3884 9272 3936
rect 11244 4097 11253 4131
rect 11253 4097 11287 4131
rect 11287 4097 11296 4131
rect 11244 4088 11296 4097
rect 11336 4020 11388 4072
rect 13452 4020 13504 4072
rect 13176 3952 13228 4004
rect 11520 3884 11572 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 1952 3680 2004 3732
rect 2872 3680 2924 3732
rect 3516 3723 3568 3732
rect 1676 3612 1728 3664
rect 2504 3612 2556 3664
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 5632 3680 5684 3732
rect 7012 3680 7064 3732
rect 7932 3680 7984 3732
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 10048 3680 10100 3732
rect 10968 3680 11020 3732
rect 12624 3680 12676 3732
rect 6000 3612 6052 3664
rect 6184 3655 6236 3664
rect 6184 3621 6193 3655
rect 6193 3621 6227 3655
rect 6227 3621 6236 3655
rect 6184 3612 6236 3621
rect 6736 3612 6788 3664
rect 9036 3655 9088 3664
rect 2044 3544 2096 3596
rect 2136 3476 2188 3528
rect 3148 3544 3200 3596
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 3240 3519 3292 3528
rect 2780 3476 2832 3485
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 4344 3544 4396 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 6920 3587 6972 3596
rect 5448 3544 5500 3553
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4436 3519 4488 3528
rect 4252 3476 4304 3485
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 5816 3476 5868 3528
rect 1768 3408 1820 3460
rect 2964 3408 3016 3460
rect 3332 3408 3384 3460
rect 4344 3408 4396 3460
rect 4804 3408 4856 3460
rect 4988 3408 5040 3460
rect 6552 3451 6604 3460
rect 6552 3417 6561 3451
rect 6561 3417 6595 3451
rect 6595 3417 6604 3451
rect 6552 3408 6604 3417
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 2780 3340 2832 3392
rect 3056 3383 3108 3392
rect 3056 3349 3065 3383
rect 3065 3349 3099 3383
rect 3099 3349 3108 3383
rect 3056 3340 3108 3349
rect 3148 3340 3200 3392
rect 3516 3340 3568 3392
rect 4252 3340 4304 3392
rect 4712 3383 4764 3392
rect 4712 3349 4721 3383
rect 4721 3349 4755 3383
rect 4755 3349 4764 3383
rect 4712 3340 4764 3349
rect 5356 3340 5408 3392
rect 5816 3340 5868 3392
rect 6920 3553 6929 3587
rect 6929 3553 6963 3587
rect 6963 3553 6972 3587
rect 6920 3544 6972 3553
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 7564 3544 7616 3596
rect 8024 3544 8076 3596
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 7564 3451 7616 3460
rect 7564 3417 7573 3451
rect 7573 3417 7607 3451
rect 7607 3417 7616 3451
rect 7564 3408 7616 3417
rect 7840 3408 7892 3460
rect 8668 3476 8720 3528
rect 8760 3451 8812 3460
rect 8760 3417 8769 3451
rect 8769 3417 8803 3451
rect 8803 3417 8812 3451
rect 8760 3408 8812 3417
rect 9036 3621 9045 3655
rect 9045 3621 9079 3655
rect 9079 3621 9088 3655
rect 9036 3612 9088 3621
rect 12992 3612 13044 3664
rect 10140 3544 10192 3596
rect 11336 3544 11388 3596
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 12716 3476 12768 3528
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 7288 3340 7340 3392
rect 7380 3340 7432 3392
rect 7472 3340 7524 3392
rect 10048 3340 10100 3392
rect 10416 3408 10468 3460
rect 10784 3451 10836 3460
rect 10784 3417 10793 3451
rect 10793 3417 10827 3451
rect 10827 3417 10836 3451
rect 10784 3408 10836 3417
rect 12808 3451 12860 3460
rect 11152 3340 11204 3392
rect 12532 3340 12584 3392
rect 12808 3417 12817 3451
rect 12817 3417 12851 3451
rect 12851 3417 12860 3451
rect 12808 3408 12860 3417
rect 13176 3340 13228 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 3240 3136 3292 3188
rect 4528 3136 4580 3188
rect 5080 3179 5132 3188
rect 5080 3145 5089 3179
rect 5089 3145 5123 3179
rect 5123 3145 5132 3179
rect 5080 3136 5132 3145
rect 5540 3136 5592 3188
rect 6644 3136 6696 3188
rect 8024 3136 8076 3188
rect 8392 3136 8444 3188
rect 9312 3136 9364 3188
rect 13452 3179 13504 3188
rect 2780 3111 2832 3120
rect 2780 3077 2789 3111
rect 2789 3077 2823 3111
rect 2823 3077 2832 3111
rect 2780 3068 2832 3077
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 1860 2932 1912 2984
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2964 3043 3016 3052
rect 2412 3000 2464 3009
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 2688 2975 2740 2984
rect 2688 2941 2697 2975
rect 2697 2941 2731 2975
rect 2731 2941 2740 2975
rect 2688 2932 2740 2941
rect 3056 2932 3108 2984
rect 3608 3000 3660 3052
rect 4068 2932 4120 2984
rect 3516 2864 3568 2916
rect 8576 3068 8628 3120
rect 8760 3068 8812 3120
rect 10416 3068 10468 3120
rect 11152 3111 11204 3120
rect 11152 3077 11161 3111
rect 11161 3077 11195 3111
rect 11195 3077 11204 3111
rect 11152 3068 11204 3077
rect 11244 3068 11296 3120
rect 11428 3068 11480 3120
rect 11888 3111 11940 3120
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5448 3043 5500 3052
rect 5172 3000 5224 3009
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 6000 3043 6052 3052
rect 5356 2932 5408 2984
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 4896 2864 4948 2916
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 6736 3000 6788 3052
rect 7104 3043 7156 3052
rect 7104 3009 7113 3043
rect 7113 3009 7147 3043
rect 7147 3009 7156 3043
rect 7104 3000 7156 3009
rect 7380 3000 7432 3052
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 11888 3077 11897 3111
rect 11897 3077 11931 3111
rect 11931 3077 11940 3111
rect 11888 3068 11940 3077
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 12624 3000 12676 3052
rect 13268 3043 13320 3052
rect 13268 3009 13277 3043
rect 13277 3009 13311 3043
rect 13311 3009 13320 3043
rect 13268 3000 13320 3009
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 7288 2932 7340 2984
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 11244 2932 11296 2984
rect 6000 2864 6052 2916
rect 9312 2864 9364 2916
rect 10876 2864 10928 2916
rect 5080 2796 5132 2848
rect 6460 2796 6512 2848
rect 9956 2796 10008 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 6736 2592 6788 2644
rect 7656 2592 7708 2644
rect 10968 2592 11020 2644
rect 11704 2592 11756 2644
rect 2688 2456 2740 2508
rect 4988 2524 5040 2576
rect 1676 2388 1728 2440
rect 2596 2388 2648 2440
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4804 2499 4856 2508
rect 4068 2456 4120 2465
rect 4804 2465 4813 2499
rect 4813 2465 4847 2499
rect 4847 2465 4856 2499
rect 4804 2456 4856 2465
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 2044 2320 2096 2372
rect 2780 2252 2832 2304
rect 3608 2320 3660 2372
rect 5080 2388 5132 2440
rect 5724 2456 5776 2508
rect 7472 2524 7524 2576
rect 11336 2524 11388 2576
rect 7656 2456 7708 2508
rect 8116 2456 8168 2508
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 5816 2252 5868 2304
rect 6276 2252 6328 2304
rect 7380 2320 7432 2372
rect 7840 2388 7892 2440
rect 7932 2320 7984 2372
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8668 2431 8720 2440
rect 8392 2388 8444 2397
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 13084 2431 13136 2440
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 9220 2363 9272 2372
rect 9220 2329 9229 2363
rect 9229 2329 9263 2363
rect 9263 2329 9272 2363
rect 9220 2320 9272 2329
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 11060 2320 11112 2372
rect 13268 2320 13320 2372
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 12716 2252 12768 2304
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 2688 2048 2740 2100
rect 3608 2048 3660 2100
rect 4068 2091 4120 2100
rect 4068 2057 4077 2091
rect 4077 2057 4111 2091
rect 4111 2057 4120 2091
rect 4068 2048 4120 2057
rect 7656 2048 7708 2100
rect 9588 2048 9640 2100
rect 10416 2091 10468 2100
rect 4988 1980 5040 2032
rect 5540 2023 5592 2032
rect 5540 1989 5549 2023
rect 5549 1989 5583 2023
rect 5583 1989 5592 2023
rect 5540 1980 5592 1989
rect 6736 2023 6788 2032
rect 1676 1955 1728 1964
rect 1676 1921 1685 1955
rect 1685 1921 1719 1955
rect 1719 1921 1728 1955
rect 1676 1912 1728 1921
rect 1860 1955 1912 1964
rect 1860 1921 1869 1955
rect 1869 1921 1903 1955
rect 1903 1921 1912 1955
rect 1860 1912 1912 1921
rect 2044 1955 2096 1964
rect 2044 1921 2053 1955
rect 2053 1921 2087 1955
rect 2087 1921 2096 1955
rect 2044 1912 2096 1921
rect 5816 1955 5868 1964
rect 5816 1921 5825 1955
rect 5825 1921 5859 1955
rect 5859 1921 5868 1955
rect 5816 1912 5868 1921
rect 3332 1844 3384 1896
rect 2504 1708 2556 1760
rect 6000 1751 6052 1760
rect 6000 1717 6009 1751
rect 6009 1717 6043 1751
rect 6043 1717 6052 1751
rect 6000 1708 6052 1717
rect 6736 1989 6745 2023
rect 6745 1989 6779 2023
rect 6779 1989 6788 2023
rect 6736 1980 6788 1989
rect 7748 1980 7800 2032
rect 9680 1980 9732 2032
rect 8024 1912 8076 1964
rect 10416 2057 10425 2091
rect 10425 2057 10459 2091
rect 10459 2057 10468 2091
rect 10416 2048 10468 2057
rect 11060 2091 11112 2100
rect 11060 2057 11069 2091
rect 11069 2057 11103 2091
rect 11103 2057 11112 2091
rect 11060 2048 11112 2057
rect 11244 2048 11296 2100
rect 11428 2048 11480 2100
rect 13084 2048 13136 2100
rect 13268 2091 13320 2100
rect 13268 2057 13277 2091
rect 13277 2057 13311 2091
rect 13311 2057 13320 2091
rect 13268 2048 13320 2057
rect 11796 1980 11848 2032
rect 11888 1980 11940 2032
rect 11244 1955 11296 1964
rect 7288 1844 7340 1896
rect 7380 1844 7432 1896
rect 8944 1887 8996 1896
rect 8944 1853 8953 1887
rect 8953 1853 8987 1887
rect 8987 1853 8996 1887
rect 8944 1844 8996 1853
rect 11244 1921 11253 1955
rect 11253 1921 11287 1955
rect 11287 1921 11296 1955
rect 11244 1912 11296 1921
rect 11336 1912 11388 1964
rect 7472 1708 7524 1760
rect 7932 1708 7984 1760
rect 11060 1844 11112 1896
rect 11152 1776 11204 1828
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 3332 1547 3384 1556
rect 3332 1513 3341 1547
rect 3341 1513 3375 1547
rect 3375 1513 3384 1547
rect 3332 1504 3384 1513
rect 7472 1504 7524 1556
rect 2872 1479 2924 1488
rect 2872 1445 2881 1479
rect 2881 1445 2915 1479
rect 2915 1445 2924 1479
rect 2872 1436 2924 1445
rect 5080 1436 5132 1488
rect 7748 1479 7800 1488
rect 7748 1445 7757 1479
rect 7757 1445 7791 1479
rect 7791 1445 7800 1479
rect 7748 1436 7800 1445
rect 9220 1504 9272 1556
rect 3608 1368 3660 1420
rect 1400 1343 1452 1352
rect 1400 1309 1409 1343
rect 1409 1309 1443 1343
rect 1443 1309 1452 1343
rect 1400 1300 1452 1309
rect 4068 1232 4120 1284
rect 6000 1368 6052 1420
rect 6368 1368 6420 1420
rect 4712 1343 4764 1352
rect 4712 1309 4721 1343
rect 4721 1309 4755 1343
rect 4755 1309 4764 1343
rect 4712 1300 4764 1309
rect 4804 1343 4856 1352
rect 4804 1309 4813 1343
rect 4813 1309 4847 1343
rect 4847 1309 4856 1343
rect 4988 1343 5040 1352
rect 4804 1300 4856 1309
rect 4988 1309 4997 1343
rect 4997 1309 5031 1343
rect 5031 1309 5040 1343
rect 4988 1300 5040 1309
rect 5632 1300 5684 1352
rect 7104 1300 7156 1352
rect 7564 1368 7616 1420
rect 7472 1343 7524 1352
rect 7472 1309 7481 1343
rect 7481 1309 7515 1343
rect 7515 1309 7524 1343
rect 7472 1300 7524 1309
rect 7840 1368 7892 1420
rect 8668 1368 8720 1420
rect 9680 1411 9732 1420
rect 7932 1343 7984 1352
rect 7380 1275 7432 1284
rect 7380 1241 7389 1275
rect 7389 1241 7423 1275
rect 7423 1241 7432 1275
rect 7380 1232 7432 1241
rect 7932 1309 7941 1343
rect 7941 1309 7975 1343
rect 7975 1309 7984 1343
rect 7932 1300 7984 1309
rect 9036 1300 9088 1352
rect 9220 1343 9272 1352
rect 9220 1309 9229 1343
rect 9229 1309 9263 1343
rect 9263 1309 9272 1343
rect 9220 1300 9272 1309
rect 9404 1343 9456 1352
rect 9404 1309 9413 1343
rect 9413 1309 9447 1343
rect 9447 1309 9456 1343
rect 9404 1300 9456 1309
rect 9680 1377 9689 1411
rect 9689 1377 9723 1411
rect 9723 1377 9732 1411
rect 9680 1368 9732 1377
rect 9956 1300 10008 1352
rect 11244 1368 11296 1420
rect 11060 1300 11112 1352
rect 11520 1343 11572 1352
rect 11520 1309 11529 1343
rect 11529 1309 11563 1343
rect 11563 1309 11572 1343
rect 11520 1300 11572 1309
rect 11796 1368 11848 1420
rect 11888 1343 11940 1352
rect 11888 1309 11897 1343
rect 11897 1309 11931 1343
rect 11931 1309 11940 1343
rect 11888 1300 11940 1309
rect 12624 1343 12676 1352
rect 12624 1309 12633 1343
rect 12633 1309 12667 1343
rect 12667 1309 12676 1343
rect 12624 1300 12676 1309
rect 10968 1232 11020 1284
rect 8576 1164 8628 1216
rect 8944 1164 8996 1216
rect 11152 1164 11204 1216
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
<< metal2 >>
rect 570 14200 626 15000
rect 1674 14362 1730 15000
rect 1674 14334 1992 14362
rect 1674 14200 1730 14334
rect 584 10606 612 14200
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1412 12617 1440 13126
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1398 12608 1454 12617
rect 1398 12543 1454 12552
rect 1780 11762 1808 12718
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1398 11656 1454 11665
rect 1398 11591 1400 11600
rect 1452 11591 1454 11600
rect 1400 11562 1452 11568
rect 1412 11218 1440 11562
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 572 10600 624 10606
rect 572 10542 624 10548
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9654 1716 9862
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1780 9178 1808 9522
rect 1872 9382 1900 13262
rect 1964 12918 1992 14334
rect 2870 14200 2926 15000
rect 3330 14512 3386 14521
rect 3330 14447 3386 14456
rect 2884 13462 2912 14200
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 1952 12912 2004 12918
rect 1952 12854 2004 12860
rect 2056 12238 2084 13194
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2240 11830 2268 12650
rect 2608 12238 2636 12786
rect 2700 12374 2728 13194
rect 2792 12986 2820 13194
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 3068 12850 3096 13194
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11830 2636 12174
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 3068 11762 3096 12786
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2700 11286 2728 11698
rect 2872 11688 2924 11694
rect 2792 11636 2872 11642
rect 2792 11630 2924 11636
rect 2792 11614 2912 11630
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1964 9994 1992 10950
rect 2332 10674 2360 11086
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2700 10538 2728 11222
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1964 9654 1992 9930
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 2700 9518 2728 9998
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8498 1624 8774
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 2700 8430 2728 9114
rect 2792 9042 2820 11614
rect 3160 11014 3188 13126
rect 3344 12102 3372 14447
rect 3974 14200 4030 15000
rect 5170 14200 5226 15000
rect 6274 14200 6330 15000
rect 7470 14200 7526 15000
rect 8574 14200 8630 15000
rect 9770 14362 9826 15000
rect 10874 14362 10930 15000
rect 9770 14334 9904 14362
rect 9770 14200 9826 14334
rect 3514 13560 3570 13569
rect 3514 13495 3516 13504
rect 3568 13495 3570 13504
rect 3516 13466 3568 13472
rect 3528 13326 3556 13466
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3436 12374 3464 12786
rect 3896 12714 3924 13194
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3436 11762 3464 12310
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3528 11694 3556 12650
rect 3988 12322 4016 14200
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4172 12628 4200 13262
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4080 12600 4200 12628
rect 4080 12442 4108 12600
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4172 12322 4200 12378
rect 3988 12294 4200 12322
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11830 3648 12038
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11218 3648 11494
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3804 11082 3832 11698
rect 3988 11150 4016 11698
rect 4632 11626 4660 12786
rect 4816 12238 4844 13194
rect 4908 12374 4936 13262
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 5000 12730 5028 13126
rect 5092 12850 5120 13262
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5000 12702 5120 12730
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 5000 12306 5028 12378
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 5092 12170 5120 12702
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2884 9994 2912 10610
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2884 9654 2912 9930
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2976 9042 3004 9862
rect 3068 9518 3096 10406
rect 3160 10033 3188 10950
rect 3330 10704 3386 10713
rect 3620 10674 3648 11018
rect 3698 10976 3754 10985
rect 3698 10911 3754 10920
rect 3712 10810 3740 10911
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3516 10668 3568 10674
rect 3386 10648 3464 10656
rect 3330 10639 3332 10648
rect 3384 10628 3464 10648
rect 3332 10610 3384 10616
rect 3240 10056 3292 10062
rect 3146 10024 3202 10033
rect 3292 10016 3372 10044
rect 3240 9998 3292 10004
rect 3146 9959 3202 9968
rect 3160 9926 3188 9959
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3252 9761 3280 9862
rect 3238 9752 3294 9761
rect 3238 9687 3294 9696
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3068 8906 3096 9454
rect 3344 9450 3372 10016
rect 3436 9722 3464 10628
rect 3516 10610 3568 10616
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3528 10470 3556 10610
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3606 9752 3662 9761
rect 3424 9716 3476 9722
rect 3606 9687 3662 9696
rect 3424 9658 3476 9664
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3344 8974 3372 9386
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8498 2820 8774
rect 3344 8566 3372 8910
rect 3436 8906 3464 9522
rect 3620 9178 3648 9687
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 1412 1358 1440 8366
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 1676 8016 1728 8022
rect 3252 7993 3280 8230
rect 3712 8090 3740 10746
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 9586 4016 9998
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4724 9353 4752 11698
rect 4816 11694 4844 11766
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4816 10985 4844 11630
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4908 11121 4936 11154
rect 5000 11150 5028 12038
rect 5184 11286 5212 14200
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5276 11762 5304 12854
rect 5460 12850 5488 13126
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5262 11656 5318 11665
rect 5262 11591 5318 11600
rect 5276 11354 5304 11591
rect 5368 11558 5396 12582
rect 5644 12442 5672 13194
rect 6196 12918 6224 13262
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 6090 12200 6146 12209
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 4988 11144 5040 11150
rect 4894 11112 4950 11121
rect 4988 11086 5040 11092
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 4894 11047 4950 11056
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 4802 10976 4858 10985
rect 4802 10911 4858 10920
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4908 10062 4936 10678
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9722 4936 9998
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5092 9654 5120 10134
rect 5184 10130 5212 11018
rect 5276 10985 5304 11018
rect 5262 10976 5318 10985
rect 5262 10911 5318 10920
rect 5368 10810 5396 11086
rect 5460 11014 5488 11698
rect 5552 11354 5580 12174
rect 5724 12164 5776 12170
rect 5908 12164 5960 12170
rect 5776 12124 5856 12152
rect 5724 12106 5776 12112
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5276 10538 5304 10678
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5736 10198 5764 11630
rect 5828 10792 5856 12124
rect 6090 12135 6092 12144
rect 5908 12106 5960 12112
rect 6144 12135 6146 12144
rect 6092 12106 6144 12112
rect 5920 12073 5948 12106
rect 5906 12064 5962 12073
rect 5906 11999 5962 12008
rect 6104 11830 6132 12106
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6196 11898 6224 12038
rect 6288 11898 6316 14200
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7024 13326 7052 13738
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12918 7052 13126
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6380 12238 6408 12786
rect 6918 12336 6974 12345
rect 6552 12300 6604 12306
rect 6918 12271 6974 12280
rect 6552 12242 6604 12248
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6564 11898 6592 12242
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5920 11150 5948 11494
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5828 10764 5948 10792
rect 5814 10704 5870 10713
rect 5814 10639 5816 10648
rect 5868 10639 5870 10648
rect 5816 10610 5868 10616
rect 5920 10577 5948 10764
rect 5906 10568 5962 10577
rect 5906 10503 5962 10512
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5460 9654 5488 9862
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4710 9344 4766 9353
rect 4214 9276 4522 9285
rect 4710 9279 4766 9288
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3790 8800 3846 8809
rect 3790 8735 3846 8744
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 1676 7958 1728 7964
rect 2502 7984 2558 7993
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1504 7002 1532 7482
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1504 6390 1532 6938
rect 1492 6384 1544 6390
rect 1492 6326 1544 6332
rect 1596 6202 1624 7822
rect 1504 6174 1624 6202
rect 1504 6118 1532 6174
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1582 6080 1638 6089
rect 1504 5710 1532 6054
rect 1582 6015 1638 6024
rect 1596 5846 1624 6015
rect 1584 5840 1636 5846
rect 1584 5782 1636 5788
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1596 5556 1624 5782
rect 1688 5642 1716 7958
rect 2502 7919 2558 7928
rect 3238 7984 3294 7993
rect 3238 7919 3294 7928
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 1780 7342 1808 7822
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1780 6458 1808 7278
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1780 6322 1808 6394
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1872 6186 1900 7754
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 1872 5710 1900 6122
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1964 5574 1992 7686
rect 2148 7546 2176 7822
rect 2516 7546 2544 7919
rect 3252 7886 3280 7919
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3804 7818 3832 8735
rect 3988 8498 4016 8978
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4448 8498 4476 8910
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4436 8492 4488 8498
rect 4488 8452 4660 8480
rect 4436 8434 4488 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8090 4660 8452
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3896 7886 3924 7958
rect 4724 7954 4752 9279
rect 4908 8906 4936 9522
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5276 8906 5304 9386
rect 5644 8974 5672 9998
rect 5736 9926 5764 10134
rect 5920 10062 5948 10503
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 6012 9586 6040 11494
rect 6288 11286 6316 11834
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6276 11280 6328 11286
rect 6380 11257 6408 11766
rect 6656 11762 6684 12106
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6276 11222 6328 11228
rect 6366 11248 6422 11257
rect 6092 10668 6144 10674
rect 6196 10656 6224 11222
rect 6472 11218 6500 11698
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6366 11183 6422 11192
rect 6460 11212 6512 11218
rect 6276 10668 6328 10674
rect 6196 10628 6276 10656
rect 6092 10610 6144 10616
rect 6276 10610 6328 10616
rect 6104 9994 6132 10610
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6012 8974 6040 9522
rect 6104 9518 6132 9930
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6196 9178 6224 10134
rect 6288 10062 6316 10202
rect 6380 10130 6408 11183
rect 6460 11154 6512 11160
rect 6472 10810 6500 11154
rect 6564 11132 6592 11630
rect 6644 11144 6696 11150
rect 6564 11104 6644 11132
rect 6644 11086 6696 11092
rect 6748 11082 6776 11630
rect 6932 11354 6960 12271
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7024 11286 7052 12854
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7208 12238 7236 12786
rect 7300 12306 7328 13194
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7392 12170 7420 13262
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7102 12064 7158 12073
rect 7102 11999 7158 12008
rect 7116 11801 7144 11999
rect 7102 11792 7158 11801
rect 7484 11762 7512 14200
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7576 13326 7604 13398
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 12850 7604 13126
rect 7668 12986 7696 13398
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8588 13274 8616 14200
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8772 13326 8800 13806
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 13462 9076 13670
rect 9036 13456 9088 13462
rect 8850 13424 8906 13433
rect 9036 13398 9088 13404
rect 9324 13394 9352 13874
rect 9312 13388 9364 13394
rect 8850 13359 8906 13368
rect 8760 13320 8812 13326
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7668 12374 7696 12650
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7840 12300 7892 12306
rect 7944 12288 7972 13194
rect 8036 12918 8064 13194
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 7892 12260 7972 12288
rect 7840 12242 7892 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7102 11727 7158 11736
rect 7472 11756 7524 11762
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6840 11014 6868 11086
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6472 10470 6500 10746
rect 6564 10606 6592 10950
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6472 10266 6500 10406
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6564 9994 6592 10542
rect 7116 10538 7144 11727
rect 7472 11698 7524 11704
rect 7378 11520 7434 11529
rect 7378 11455 7434 11464
rect 7194 11384 7250 11393
rect 7194 11319 7250 11328
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6564 9722 6592 9930
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6656 9654 6684 9930
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 4908 8362 4936 8842
rect 5000 8634 5028 8842
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5644 8498 5672 8910
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4802 7984 4858 7993
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 4712 7948 4764 7954
rect 4802 7919 4858 7928
rect 4712 7890 4764 7896
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2240 6322 2268 7142
rect 2608 6372 2636 7686
rect 2688 6724 2740 6730
rect 2792 6712 2820 7754
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2870 7032 2926 7041
rect 2870 6967 2926 6976
rect 2740 6684 2820 6712
rect 2688 6666 2740 6672
rect 2608 6344 2728 6372
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 2332 5710 2360 5782
rect 2700 5710 2728 6344
rect 2884 6322 2912 6967
rect 2976 6866 3004 7142
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6458 3004 6666
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2884 5914 2912 6258
rect 3068 6186 3096 7754
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3528 7002 3556 7278
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3804 6798 3832 7754
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3436 6186 3464 6734
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3712 6118 3740 6258
rect 3896 6236 3924 7482
rect 3988 7342 4016 7890
rect 4816 7886 4844 7919
rect 6104 7886 6132 8366
rect 6196 7886 6224 9114
rect 6380 8906 6408 9590
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6472 9178 6500 9522
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6380 8498 6408 8842
rect 6656 8838 6684 9590
rect 6748 9450 6776 10406
rect 6828 10056 6880 10062
rect 6932 10044 6960 10474
rect 6880 10016 6960 10044
rect 6828 9998 6880 10004
rect 6826 9480 6882 9489
rect 6736 9444 6788 9450
rect 6826 9415 6828 9424
rect 6736 9386 6788 9392
rect 6880 9415 6882 9424
rect 6828 9386 6880 9392
rect 6932 9110 6960 10016
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7024 9217 7052 9930
rect 7208 9926 7236 11319
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 7300 11082 7328 11222
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7392 10606 7420 11455
rect 7484 11370 7512 11698
rect 7576 11558 7604 12174
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7484 11354 7604 11370
rect 7484 11348 7616 11354
rect 7484 11342 7564 11348
rect 7564 11290 7616 11296
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7472 11144 7524 11150
rect 7576 11121 7604 11154
rect 7472 11086 7524 11092
rect 7562 11112 7618 11121
rect 7484 10713 7512 11086
rect 7562 11047 7618 11056
rect 7470 10704 7526 10713
rect 7470 10639 7526 10648
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7286 10296 7342 10305
rect 7286 10231 7342 10240
rect 7300 10130 7328 10231
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7300 9654 7328 9930
rect 7288 9648 7340 9654
rect 7392 9625 7420 10542
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7288 9590 7340 9596
rect 7378 9616 7434 9625
rect 7104 9580 7156 9586
rect 7156 9540 7236 9568
rect 7378 9551 7434 9560
rect 7104 9522 7156 9528
rect 7208 9500 7236 9540
rect 7208 9472 7328 9500
rect 7010 9208 7066 9217
rect 7066 9178 7144 9194
rect 7066 9172 7156 9178
rect 7066 9166 7104 9172
rect 7010 9143 7066 9152
rect 7104 9114 7156 9120
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7196 9104 7248 9110
rect 7300 9081 7328 9472
rect 7196 9046 7248 9052
rect 7286 9072 7342 9081
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6840 8498 6868 8910
rect 7208 8906 7236 9046
rect 7286 9007 7342 9016
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7392 8820 7420 9551
rect 7484 9382 7512 10406
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7576 10062 7604 10134
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7576 9110 7604 9862
rect 7668 9178 7696 12038
rect 7944 11898 7972 12260
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11898 8064 12038
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7852 11778 7880 11834
rect 7748 11756 7800 11762
rect 7852 11750 7972 11778
rect 7748 11698 7800 11704
rect 7760 11529 7788 11698
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7746 11520 7802 11529
rect 7746 11455 7802 11464
rect 7746 10704 7802 10713
rect 7746 10639 7802 10648
rect 7760 10062 7788 10639
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7760 9160 7788 9998
rect 7852 9722 7880 11630
rect 7944 11558 7972 11750
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7944 11150 7972 11290
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8022 11112 8078 11121
rect 8022 11047 8078 11056
rect 7932 11008 7984 11014
rect 8036 10996 8064 11047
rect 7984 10968 8064 10996
rect 7932 10950 7984 10956
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7944 10062 7972 10610
rect 8036 10606 8064 10968
rect 8128 10810 8156 13262
rect 8588 13246 8708 13274
rect 8760 13262 8812 13268
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8214 13084 8522 13093
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13019 8522 13028
rect 8588 12306 8616 13126
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8214 11996 8522 12005
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11931 8522 11940
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8220 11218 8248 11766
rect 8484 11756 8536 11762
rect 8536 11716 8616 11744
rect 8484 11698 8536 11704
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8214 10908 8522 10917
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10843 8522 10852
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8024 10600 8076 10606
rect 8392 10600 8444 10606
rect 8024 10542 8076 10548
rect 8220 10560 8392 10588
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7840 9172 7892 9178
rect 7760 9132 7840 9160
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7300 8792 7420 8820
rect 7300 8566 7328 8792
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6380 8294 6408 8434
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7410 4108 7686
rect 5368 7410 5396 7754
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4264 6458 4292 6666
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4632 6390 4660 7142
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 3976 6248 4028 6254
rect 3896 6208 3976 6236
rect 3976 6190 4028 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 1504 5528 1624 5556
rect 1952 5568 2004 5574
rect 1504 5370 1532 5528
rect 1952 5510 2004 5516
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 2044 5160 2096 5166
rect 2042 5128 2044 5137
rect 2096 5128 2098 5137
rect 1952 5092 2004 5098
rect 2240 5098 2268 5510
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2042 5063 2098 5072
rect 2228 5092 2280 5098
rect 1952 5034 2004 5040
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1492 4548 1544 4554
rect 1492 4490 1544 4496
rect 1504 4214 1532 4490
rect 1492 4208 1544 4214
rect 1490 4176 1492 4185
rect 1544 4176 1546 4185
rect 1490 4111 1546 4120
rect 1688 3670 1716 4558
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1780 3466 1808 4082
rect 1964 4078 1992 5034
rect 2056 4486 2084 5063
rect 2228 5034 2280 5040
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1964 3738 1992 4014
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2056 3602 2084 4422
rect 2148 4146 2176 4694
rect 2424 4570 2452 5170
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4622 2820 5102
rect 2884 4622 2912 5578
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 4622 3096 5510
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3514 5128 3570 5137
rect 3514 5063 3570 5072
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 2780 4616 2832 4622
rect 2424 4542 2728 4570
rect 2780 4558 2832 4564
rect 2872 4616 2924 4622
rect 3056 4616 3108 4622
rect 2872 4558 2924 4564
rect 2976 4576 3056 4604
rect 2700 4486 2728 4542
rect 2688 4480 2740 4486
rect 2410 4448 2466 4457
rect 2688 4422 2740 4428
rect 2410 4383 2466 4392
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2148 3534 2176 4082
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 2424 3058 2452 4383
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 3670 2544 4082
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1596 2281 1624 2994
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1582 2272 1638 2281
rect 1582 2207 1638 2216
rect 1688 1970 1716 2382
rect 1872 1970 1900 2926
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 2056 1970 2084 2314
rect 1676 1964 1728 1970
rect 1676 1906 1728 1912
rect 1860 1964 1912 1970
rect 1860 1906 1912 1912
rect 2044 1964 2096 1970
rect 2044 1906 2096 1912
rect 2516 1766 2544 3606
rect 2608 2446 2636 4014
rect 2700 3398 2728 4422
rect 2792 3534 2820 4558
rect 2884 4214 2912 4558
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2884 3738 2912 4014
rect 2976 3942 3004 4576
rect 3056 4558 3108 4564
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3160 4282 3188 4558
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3344 4146 3372 4626
rect 3528 4468 3556 5063
rect 3620 4690 3648 5306
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3608 4480 3660 4486
rect 3528 4440 3608 4468
rect 3608 4422 3660 4428
rect 3620 4214 3648 4422
rect 3608 4208 3660 4214
rect 3514 4176 3570 4185
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3332 4140 3384 4146
rect 3608 4150 3660 4156
rect 3514 4111 3570 4120
rect 3332 4082 3384 4088
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2686 3224 2742 3233
rect 2686 3159 2742 3168
rect 2700 2990 2728 3159
rect 2792 3126 2820 3334
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2976 3058 3004 3402
rect 3068 3398 3096 4082
rect 3160 3602 3188 4082
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3160 3210 3188 3334
rect 3068 3182 3188 3210
rect 3252 3194 3280 3470
rect 3344 3466 3372 4082
rect 3528 3738 3556 4111
rect 3606 4040 3662 4049
rect 3606 3975 3608 3984
rect 3660 3975 3662 3984
rect 3608 3946 3660 3952
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3528 3398 3556 3674
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3240 3188 3292 3194
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3068 2990 3096 3182
rect 3240 3130 3292 3136
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2700 2514 2728 2926
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2700 2106 2728 2450
rect 3528 2446 3556 2858
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3620 2378 3648 2994
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2688 2100 2740 2106
rect 2688 2042 2740 2048
rect 2504 1760 2556 1766
rect 2504 1702 2556 1708
rect 1400 1352 1452 1358
rect 1400 1294 1452 1300
rect 2792 513 2820 2246
rect 3620 2106 3648 2314
rect 3608 2100 3660 2106
rect 3608 2042 3660 2048
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 3344 1562 3372 1838
rect 3332 1556 3384 1562
rect 3332 1498 3384 1504
rect 2872 1488 2924 1494
rect 2872 1430 2924 1436
rect 2884 1329 2912 1430
rect 3620 1426 3648 2042
rect 3608 1420 3660 1426
rect 3608 1362 3660 1368
rect 2870 1320 2926 1329
rect 2870 1255 2926 1264
rect 3712 800 3740 6054
rect 4080 5896 4108 6122
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4160 5908 4212 5914
rect 4080 5868 4160 5896
rect 4160 5850 4212 5856
rect 4632 5778 4660 6326
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 3896 5302 3924 5510
rect 4172 5370 4200 5510
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3804 4622 3832 5102
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3896 4282 3924 4966
rect 3988 4622 4016 5170
rect 4540 5098 4568 5646
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3988 3738 4016 4558
rect 4436 4480 4488 4486
rect 4434 4448 4436 4457
rect 4488 4448 4490 4457
rect 4434 4383 4490 4392
rect 4632 4146 4660 5714
rect 4724 5710 4752 6054
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4724 4690 4752 5646
rect 4816 5302 4844 7210
rect 5276 6866 5304 7278
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4908 5710 4936 6054
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 5000 5114 5028 5850
rect 5276 5692 5304 6802
rect 5368 6118 5396 7346
rect 5460 6322 5488 7822
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5552 7002 5580 7686
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5644 6662 5672 7822
rect 6840 7818 6868 8434
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 8129 6960 8298
rect 7484 8294 7512 8910
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 6918 8120 6974 8129
rect 7484 8090 7512 8230
rect 6918 8055 6974 8064
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7562 7984 7618 7993
rect 7668 7954 7696 8434
rect 7562 7919 7618 7928
rect 7656 7948 7708 7954
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5644 6186 5672 6598
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5448 5704 5500 5710
rect 5276 5664 5448 5692
rect 5448 5646 5500 5652
rect 5460 5370 5488 5646
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 4816 5086 5028 5114
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4632 3618 4660 3878
rect 4724 3754 4752 4626
rect 4816 4146 4844 5086
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4690 4936 4966
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4908 4554 4936 4626
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 4908 4146 4936 4490
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5000 4214 5028 4422
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4724 3726 4936 3754
rect 5092 3738 5120 4014
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4448 3590 4660 3618
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 3398 4292 3470
rect 4356 3466 4384 3538
rect 4448 3534 4476 3590
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4540 3194 4568 3470
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4712 3392 4764 3398
rect 4632 3352 4712 3380
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4632 3097 4660 3352
rect 4712 3334 4764 3340
rect 4618 3088 4674 3097
rect 4816 3058 4844 3402
rect 4618 3023 4620 3032
rect 4672 3023 4674 3032
rect 4804 3052 4856 3058
rect 4620 2994 4672 3000
rect 4804 2994 4856 3000
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4080 2514 4108 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4816 2514 4844 2994
rect 4908 2922 4936 3726
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 5000 2582 5028 3402
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5092 2854 5120 3130
rect 5184 3058 5212 4082
rect 5736 4078 5764 4490
rect 5828 4128 5856 7754
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5920 7410 5948 7686
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6840 7274 6868 7754
rect 7484 7750 7512 7822
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7300 7546 7328 7686
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6380 6322 6408 6734
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6104 5914 6132 6190
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6092 5568 6144 5574
rect 6196 5556 6224 6258
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6144 5528 6224 5556
rect 6092 5510 6144 5516
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5920 4826 5948 5170
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6196 4554 6224 5528
rect 6472 5302 6500 5578
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 5908 4140 5960 4146
rect 5828 4100 5908 4128
rect 5908 4082 5960 4088
rect 5724 4072 5776 4078
rect 5776 4032 5856 4060
rect 5724 4014 5776 4020
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5276 3738 5304 3946
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5368 2990 5396 3334
rect 5460 3058 5488 3538
rect 5644 3534 5672 3674
rect 5828 3534 5856 4032
rect 5632 3528 5684 3534
rect 5816 3528 5868 3534
rect 5684 3488 5764 3516
rect 5632 3470 5684 3476
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4080 2106 4108 2450
rect 5080 2440 5132 2446
rect 4710 2408 4766 2417
rect 5080 2382 5132 2388
rect 4710 2343 4766 2352
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4080 1290 4108 2042
rect 4214 1660 4522 1669
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1595 4522 1604
rect 4724 1358 4752 2343
rect 4988 2032 5040 2038
rect 4988 1974 5040 1980
rect 4802 1456 4858 1465
rect 4802 1391 4858 1400
rect 4816 1358 4844 1391
rect 5000 1358 5028 1974
rect 5092 1494 5120 2382
rect 5552 2038 5580 3130
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5644 2825 5672 2926
rect 5630 2816 5686 2825
rect 5630 2751 5686 2760
rect 5736 2632 5764 3488
rect 5816 3470 5868 3476
rect 5828 3398 5856 3470
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5920 3040 5948 4082
rect 6012 3670 6040 4490
rect 6196 3670 6224 4490
rect 6274 4448 6330 4457
rect 6274 4383 6330 4392
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6000 3052 6052 3058
rect 5920 3012 6000 3040
rect 6000 2994 6052 3000
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 5814 2816 5870 2825
rect 5814 2751 5870 2760
rect 5644 2604 5764 2632
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5080 1488 5132 1494
rect 5080 1430 5132 1436
rect 5644 1358 5672 2604
rect 5724 2508 5776 2514
rect 5828 2496 5856 2751
rect 5776 2468 5856 2496
rect 5724 2450 5776 2456
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 1970 5856 2246
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 6012 1766 6040 2858
rect 6288 2310 6316 4383
rect 6380 4214 6408 4558
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6000 1760 6052 1766
rect 6000 1702 6052 1708
rect 6012 1426 6040 1702
rect 6380 1426 6408 2926
rect 6472 2854 6500 4558
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6564 3466 6592 3946
rect 6656 3942 6684 4558
rect 6840 4298 6868 6938
rect 6932 6458 6960 7414
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7024 6186 7052 6666
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 6322 7144 6598
rect 7300 6458 7328 6666
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6932 5778 6960 6122
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6932 5234 6960 5714
rect 7116 5642 7144 6258
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7208 5710 7236 6054
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 7116 5302 7144 5578
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6932 4826 6960 5170
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7116 4758 7144 5238
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7116 4554 7144 4694
rect 7208 4622 7236 5646
rect 7300 4690 7328 6190
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6840 4270 7052 4298
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6826 4040 6882 4049
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6748 3670 6776 4014
rect 6826 3975 6882 3984
rect 6840 3942 6868 3975
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6656 3097 6684 3130
rect 6642 3088 6698 3097
rect 6748 3058 6776 3606
rect 6932 3602 6960 4150
rect 7024 3738 7052 4270
rect 7300 4078 7328 4626
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7392 4486 7420 4558
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 7024 3534 7052 3674
rect 7576 3602 7604 7919
rect 7656 7890 7708 7896
rect 7760 6322 7788 9132
rect 7840 9114 7892 9120
rect 7838 9072 7894 9081
rect 7838 9007 7894 9016
rect 7852 8974 7880 9007
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7852 8634 7880 8910
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7840 8492 7892 8498
rect 7944 8480 7972 9998
rect 7892 8452 7972 8480
rect 7840 8434 7892 8440
rect 7852 8022 7880 8434
rect 8036 8362 8064 10542
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8128 10266 8156 10474
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8220 10062 8248 10560
rect 8392 10542 8444 10548
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8312 10266 8340 10406
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8404 10062 8432 10406
rect 8496 10198 8524 10746
rect 8588 10724 8616 11716
rect 8680 11354 8708 13246
rect 8864 12442 8892 13359
rect 9232 13348 9312 13376
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8772 11082 8800 11834
rect 8864 11830 8892 12378
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8588 10696 8800 10724
rect 8666 10432 8722 10441
rect 8666 10367 8722 10376
rect 8484 10192 8536 10198
rect 8576 10192 8628 10198
rect 8484 10134 8536 10140
rect 8574 10160 8576 10169
rect 8628 10160 8630 10169
rect 8484 10090 8536 10096
rect 8574 10095 8630 10104
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8392 10056 8444 10062
rect 8536 10038 8616 10044
rect 8484 10032 8616 10038
rect 8496 10016 8616 10032
rect 8392 9998 8444 10004
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8128 9722 8156 9930
rect 8214 9820 8522 9829
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9755 8522 9764
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8312 9654 8524 9674
rect 8300 9648 8524 9654
rect 8220 9608 8300 9636
rect 8220 9353 8248 9608
rect 8352 9646 8524 9648
rect 8300 9590 8352 9596
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8206 9344 8262 9353
rect 8206 9279 8262 9288
rect 8114 9208 8170 9217
rect 8114 9143 8170 9152
rect 8128 8974 8156 9143
rect 8312 9081 8340 9454
rect 8298 9072 8354 9081
rect 8298 9007 8354 9016
rect 8116 8968 8168 8974
rect 8404 8945 8432 9522
rect 8116 8910 8168 8916
rect 8390 8936 8446 8945
rect 8128 8566 8156 8910
rect 8390 8871 8446 8880
rect 8496 8888 8524 9646
rect 8588 9489 8616 10016
rect 8574 9480 8630 9489
rect 8680 9450 8708 10367
rect 8772 9586 8800 10696
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8864 9450 8892 11630
rect 8956 11257 8984 12242
rect 9232 12238 9260 13348
rect 9312 13330 9364 13336
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12714 9352 13126
rect 9600 12986 9628 13262
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9508 12782 9536 12922
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12356 9720 12582
rect 9772 12368 9824 12374
rect 9692 12328 9772 12356
rect 9772 12310 9824 12316
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9496 12232 9548 12238
rect 9772 12232 9824 12238
rect 9496 12174 9548 12180
rect 9600 12192 9772 12220
rect 9128 11824 9180 11830
rect 9128 11766 9180 11772
rect 9036 11552 9088 11558
rect 9140 11529 9168 11766
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9036 11494 9088 11500
rect 9126 11520 9182 11529
rect 9048 11354 9076 11494
rect 9126 11455 9182 11464
rect 9324 11393 9352 11630
rect 9310 11384 9366 11393
rect 9036 11348 9088 11354
rect 9310 11319 9366 11328
rect 9036 11290 9088 11296
rect 8942 11248 8998 11257
rect 8942 11183 8998 11192
rect 8956 11082 8984 11183
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 9048 10674 9076 11290
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 11008 9180 11014
rect 9126 10976 9128 10985
rect 9180 10976 9182 10985
rect 9126 10911 9182 10920
rect 9232 10849 9260 11086
rect 9218 10840 9274 10849
rect 9218 10775 9274 10784
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8944 10600 8996 10606
rect 8942 10568 8944 10577
rect 8996 10568 8998 10577
rect 8942 10503 8998 10512
rect 8956 9976 8984 10503
rect 9048 10441 9076 10610
rect 9126 10568 9182 10577
rect 9126 10503 9182 10512
rect 9140 10470 9168 10503
rect 9128 10464 9180 10470
rect 9034 10432 9090 10441
rect 9128 10406 9180 10412
rect 9416 10418 9444 11698
rect 9508 11558 9536 12174
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9600 11014 9628 12192
rect 9772 12174 9824 12180
rect 9770 11928 9826 11937
rect 9770 11863 9826 11872
rect 9784 11762 9812 11863
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9678 11384 9734 11393
rect 9678 11319 9734 11328
rect 9692 11286 9720 11319
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9876 11200 9904 14334
rect 10520 14334 10930 14362
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 12306 9996 12582
rect 10060 12374 10088 12854
rect 10244 12850 10272 13262
rect 10324 13252 10376 13258
rect 10324 13194 10376 13200
rect 10336 12918 10364 13194
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 10152 11880 10180 12582
rect 10324 12368 10376 12374
rect 10322 12336 10324 12345
rect 10376 12336 10378 12345
rect 10322 12271 10378 12280
rect 10428 12220 10456 13262
rect 10520 12434 10548 14334
rect 10874 14200 10930 14334
rect 12070 14200 12126 15000
rect 13174 14362 13230 15000
rect 13004 14334 13230 14362
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10796 13326 10824 13466
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10704 12918 10732 13126
rect 10796 12986 10824 13126
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10690 12472 10746 12481
rect 10520 12406 10640 12434
rect 10690 12407 10692 12416
rect 10506 12336 10562 12345
rect 10506 12271 10562 12280
rect 10060 11852 10180 11880
rect 10336 12192 10456 12220
rect 10060 11336 10088 11852
rect 10232 11824 10284 11830
rect 10230 11792 10232 11801
rect 10284 11792 10286 11801
rect 10140 11756 10192 11762
rect 10230 11727 10286 11736
rect 10140 11698 10192 11704
rect 9968 11308 10088 11336
rect 9968 11218 9996 11308
rect 10152 11286 10180 11698
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10230 11248 10286 11257
rect 9784 11172 9904 11200
rect 9956 11212 10008 11218
rect 9678 11112 9734 11121
rect 9678 11047 9680 11056
rect 9732 11047 9734 11056
rect 9680 11018 9732 11024
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9678 10976 9734 10985
rect 9494 10840 9550 10849
rect 9494 10775 9550 10784
rect 9508 10742 9536 10775
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9600 10674 9628 10950
rect 9678 10911 9734 10920
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9416 10390 9536 10418
rect 9034 10367 9090 10376
rect 9218 10296 9274 10305
rect 9128 10260 9180 10266
rect 9048 10220 9128 10248
rect 9048 10112 9076 10220
rect 9508 10282 9536 10390
rect 9218 10231 9274 10240
rect 9416 10254 9536 10282
rect 9128 10202 9180 10208
rect 9048 10084 9168 10112
rect 9036 9988 9088 9994
rect 8956 9948 9036 9976
rect 9036 9930 9088 9936
rect 8942 9752 8998 9761
rect 8942 9687 8944 9696
rect 8996 9687 8998 9696
rect 8944 9658 8996 9664
rect 8574 9415 8630 9424
rect 8668 9444 8720 9450
rect 8588 9330 8616 9415
rect 8668 9386 8720 9392
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8944 9376 8996 9382
rect 8588 9302 8800 9330
rect 9048 9353 9076 9930
rect 9140 9926 9168 10084
rect 9128 9920 9180 9926
rect 9232 9908 9260 10231
rect 9416 10112 9444 10254
rect 9600 10169 9628 10610
rect 9692 10470 9720 10911
rect 9680 10464 9732 10470
rect 9784 10441 9812 11172
rect 10230 11183 10286 11192
rect 9956 11154 10008 11160
rect 10244 11150 10272 11183
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10232 11144 10284 11150
rect 10336 11121 10364 12192
rect 10520 11898 10548 12271
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10612 11778 10640 12406
rect 10744 12407 10746 12416
rect 10692 12378 10744 12384
rect 10692 12232 10744 12238
rect 10690 12200 10692 12209
rect 10744 12200 10746 12209
rect 10690 12135 10746 12144
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10428 11750 10640 11778
rect 10232 11086 10284 11092
rect 10322 11112 10378 11121
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9876 10792 9904 11018
rect 10060 10985 10088 11018
rect 10046 10976 10102 10985
rect 10046 10911 10102 10920
rect 10048 10804 10100 10810
rect 9876 10764 10048 10792
rect 9680 10406 9732 10412
rect 9770 10432 9826 10441
rect 9692 10266 9720 10406
rect 9770 10367 9826 10376
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9323 10084 9444 10112
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 9323 10044 9351 10084
rect 9600 10062 9628 10095
rect 9588 10056 9640 10062
rect 9323 10016 9444 10044
rect 9312 9920 9364 9926
rect 9232 9880 9312 9908
rect 9128 9862 9180 9868
rect 9312 9862 9364 9868
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 8944 9318 8996 9324
rect 9034 9344 9090 9353
rect 8772 9178 8800 9302
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8496 8860 8616 8888
rect 8214 8732 8522 8741
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8667 8522 8676
rect 8588 8634 8616 8860
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7944 6866 7972 7754
rect 8036 7426 8064 8298
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7546 8156 7686
rect 8214 7644 8522 7653
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7579 8522 7588
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8220 7426 8248 7482
rect 8036 7398 8248 7426
rect 8300 7336 8352 7342
rect 8036 7296 8300 7324
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 8036 6254 8064 7296
rect 8300 7278 8352 7284
rect 8312 6730 8340 7278
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 6254 8156 6598
rect 8214 6556 8522 6565
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6491 8522 6500
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7300 3466 7604 3482
rect 7300 3460 7616 3466
rect 7300 3454 7564 3460
rect 7300 3398 7328 3454
rect 7564 3402 7616 3408
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7392 3058 7420 3334
rect 6642 3023 6698 3032
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6748 2038 6776 2586
rect 7116 2310 7144 2994
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 6736 2032 6788 2038
rect 6736 1974 6788 1980
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 6368 1420 6420 1426
rect 6368 1362 6420 1368
rect 7116 1358 7144 2246
rect 7300 1902 7328 2926
rect 7392 2378 7420 2994
rect 7484 2582 7512 3334
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7576 2446 7604 3402
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7668 2650 7696 2994
rect 7760 2774 7788 5510
rect 8214 5468 8522 5477
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5403 8522 5412
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7852 4758 7880 5238
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 8128 4128 8156 5306
rect 8214 4380 8522 4389
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4315 8522 4324
rect 8588 4146 8616 8434
rect 8680 8090 8708 9114
rect 8956 9092 8984 9318
rect 9034 9279 9090 9288
rect 8864 9064 8984 9092
rect 8760 9036 8812 9042
rect 8864 9024 8892 9064
rect 9048 9058 9076 9279
rect 9140 9217 9168 9522
rect 9416 9217 9444 10016
rect 9494 10024 9550 10033
rect 9588 9998 9640 10004
rect 9494 9959 9550 9968
rect 9126 9208 9182 9217
rect 9126 9143 9182 9152
rect 9402 9208 9458 9217
rect 9402 9143 9458 9152
rect 9048 9030 9168 9058
rect 8812 8996 8892 9024
rect 8760 8978 8812 8984
rect 9036 8968 9088 8974
rect 8942 8936 8998 8945
rect 9036 8910 9088 8916
rect 8942 8871 8998 8880
rect 8852 8832 8904 8838
rect 8850 8800 8852 8809
rect 8904 8800 8906 8809
rect 8850 8735 8906 8744
rect 8850 8664 8906 8673
rect 8772 8622 8850 8650
rect 8772 8498 8800 8622
rect 8850 8599 8906 8608
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8772 8294 8800 8434
rect 8956 8294 8984 8871
rect 9048 8634 9076 8910
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8498 9168 9030
rect 9220 8946 9272 8952
rect 9220 8888 9272 8894
rect 9310 8936 9366 8945
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 8129 8984 8230
rect 8942 8120 8998 8129
rect 8668 8084 8720 8090
rect 8942 8055 8998 8064
rect 8668 8026 8720 8032
rect 9036 8016 9088 8022
rect 9034 7984 9036 7993
rect 9088 7984 9090 7993
rect 9034 7919 9090 7928
rect 9140 7750 9168 8434
rect 9232 8362 9260 8888
rect 9310 8871 9366 8880
rect 9324 8537 9352 8871
rect 9416 8566 9444 9143
rect 9508 9110 9536 9959
rect 9586 9616 9642 9625
rect 9784 9586 9812 10367
rect 9876 10305 9904 10764
rect 10048 10746 10100 10752
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 10046 10568 10102 10577
rect 9862 10296 9918 10305
rect 9862 10231 9918 10240
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9586 9551 9588 9560
rect 9640 9551 9642 9560
rect 9772 9580 9824 9586
rect 9588 9522 9640 9528
rect 9692 9518 9720 9549
rect 9772 9522 9824 9528
rect 9680 9512 9732 9518
rect 9678 9480 9680 9489
rect 9732 9480 9734 9489
rect 9600 9438 9678 9466
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9494 8800 9550 8809
rect 9494 8735 9550 8744
rect 9508 8634 9536 8735
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9404 8560 9456 8566
rect 9310 8528 9366 8537
rect 9404 8502 9456 8508
rect 9310 8463 9312 8472
rect 9364 8463 9366 8472
rect 9496 8492 9548 8498
rect 9312 8434 9364 8440
rect 9600 8480 9628 9438
rect 9678 9415 9734 9424
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8945 9720 8978
rect 9678 8936 9734 8945
rect 9678 8871 9734 8880
rect 9680 8492 9732 8498
rect 9548 8452 9680 8480
rect 9496 8434 9548 8440
rect 9680 8434 9732 8440
rect 9784 8430 9812 9046
rect 9876 8974 9904 10066
rect 9968 9722 9996 10542
rect 10046 10503 10102 10512
rect 10060 10266 10088 10503
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10060 10130 10088 10202
rect 10152 10130 10180 11086
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10048 9920 10100 9926
rect 10100 9880 10180 9908
rect 10048 9862 10100 9868
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9876 8566 9904 8910
rect 9968 8906 9996 9522
rect 10046 9208 10102 9217
rect 10046 9143 10048 9152
rect 10100 9143 10102 9152
rect 10048 9114 10100 9120
rect 10152 8974 10180 9880
rect 10244 9722 10272 11086
rect 10322 11047 10378 11056
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 9908 10364 10950
rect 10428 10062 10456 11750
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10520 11150 10548 11562
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10520 10418 10548 11086
rect 10612 11014 10640 11630
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10612 10674 10640 10950
rect 10704 10810 10732 12038
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10690 10704 10746 10713
rect 10600 10668 10652 10674
rect 10690 10639 10692 10648
rect 10600 10610 10652 10616
rect 10744 10639 10746 10648
rect 10692 10610 10744 10616
rect 10600 10532 10652 10538
rect 10796 10520 10824 12786
rect 10980 12345 11008 12922
rect 10966 12336 11022 12345
rect 10966 12271 11022 12280
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11286 10916 11494
rect 10980 11354 11008 12174
rect 11072 12170 11100 13262
rect 11164 12986 11192 13330
rect 11532 13258 11560 13806
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13394 11652 13670
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12238 11284 13194
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10876 11280 10928 11286
rect 11072 11234 11100 12106
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11152 11688 11204 11694
rect 11256 11665 11284 11698
rect 11152 11630 11204 11636
rect 11242 11656 11298 11665
rect 10876 11222 10928 11228
rect 10980 11206 11100 11234
rect 10874 11112 10930 11121
rect 10874 11047 10930 11056
rect 10888 10713 10916 11047
rect 10980 10985 11008 11206
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10966 10976 11022 10985
rect 10966 10911 11022 10920
rect 10968 10736 11020 10742
rect 10874 10704 10930 10713
rect 11072 10713 11100 11086
rect 11164 10810 11192 11630
rect 11242 11591 11298 11600
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10968 10678 11020 10684
rect 11058 10704 11114 10713
rect 10874 10639 10930 10648
rect 10652 10492 10824 10520
rect 10600 10474 10652 10480
rect 10520 10390 10916 10418
rect 10690 10296 10746 10305
rect 10690 10231 10746 10240
rect 10704 10062 10732 10231
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10416 9920 10468 9926
rect 10336 9880 10416 9908
rect 10416 9862 10468 9868
rect 10428 9761 10456 9862
rect 10414 9752 10470 9761
rect 10232 9716 10284 9722
rect 10414 9687 10470 9696
rect 10232 9658 10284 9664
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 10060 8838 10088 8910
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 8772 7410 8800 7686
rect 9232 7546 9260 7958
rect 9324 7886 9352 8230
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9140 6798 9168 7346
rect 9324 7290 9352 7822
rect 9416 7410 9444 8026
rect 9876 7886 9904 8502
rect 10048 8424 10100 8430
rect 10152 8412 10180 8910
rect 10244 8634 10272 9658
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10336 8945 10364 9590
rect 10322 8936 10378 8945
rect 10322 8871 10378 8880
rect 10428 8838 10456 9687
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9353 10548 9522
rect 10506 9344 10562 9353
rect 10506 9279 10562 9288
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10100 8384 10180 8412
rect 10324 8424 10376 8430
rect 10230 8392 10286 8401
rect 10048 8366 10100 8372
rect 10324 8366 10376 8372
rect 10230 8327 10286 8336
rect 10244 8294 10272 8327
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9324 7262 9628 7290
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 6458 9168 6734
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6458 9352 6598
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8864 5574 8892 5646
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 9140 4690 9168 6258
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9232 4622 9260 4966
rect 9220 4616 9272 4622
rect 8666 4584 8722 4593
rect 9220 4558 9272 4564
rect 8666 4519 8668 4528
rect 8720 4519 8722 4528
rect 8668 4490 8720 4496
rect 8208 4140 8260 4146
rect 8128 4100 8208 4128
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7944 3534 7972 3674
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7852 3058 7880 3402
rect 8036 3194 8064 3538
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8024 2984 8076 2990
rect 8128 2972 8156 4100
rect 8208 4082 8260 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 9232 3942 9260 4558
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8214 3292 8522 3301
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3227 8522 3236
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8076 2944 8156 2972
rect 8024 2926 8076 2932
rect 7760 2746 7880 2774
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7392 1902 7420 2314
rect 7288 1896 7340 1902
rect 7288 1838 7340 1844
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 4712 1352 4764 1358
rect 4712 1294 4764 1300
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5632 1352 5684 1358
rect 5632 1294 5684 1300
rect 7104 1352 7156 1358
rect 7104 1294 7156 1300
rect 7392 1290 7420 1838
rect 7472 1760 7524 1766
rect 7472 1702 7524 1708
rect 7484 1562 7512 1702
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 7484 1358 7512 1498
rect 7576 1426 7604 2382
rect 7668 2106 7696 2450
rect 7852 2446 7880 2746
rect 8036 2496 8064 2926
rect 8116 2508 8168 2514
rect 8036 2468 8116 2496
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7748 2032 7800 2038
rect 7748 1974 7800 1980
rect 7760 1494 7788 1974
rect 7748 1488 7800 1494
rect 7748 1430 7800 1436
rect 7852 1426 7880 2382
rect 7932 2372 7984 2378
rect 7932 2314 7984 2320
rect 7944 1766 7972 2314
rect 8036 1970 8064 2468
rect 8116 2450 8168 2456
rect 8404 2446 8432 3130
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8392 2440 8444 2446
rect 8390 2408 8392 2417
rect 8444 2408 8446 2417
rect 8390 2343 8446 2352
rect 8214 2204 8522 2213
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2139 8522 2148
rect 8024 1964 8076 1970
rect 8024 1906 8076 1912
rect 7932 1760 7984 1766
rect 7932 1702 7984 1708
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 7840 1420 7892 1426
rect 7840 1362 7892 1368
rect 7944 1358 7972 1702
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7932 1352 7984 1358
rect 7932 1294 7984 1300
rect 4068 1284 4120 1290
rect 4068 1226 4120 1232
rect 7380 1284 7432 1290
rect 7380 1226 7432 1232
rect 8588 1222 8616 3062
rect 8680 2446 8708 3470
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8772 3126 8800 3402
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8680 1465 8708 2382
rect 8944 1896 8996 1902
rect 8944 1838 8996 1844
rect 8666 1456 8722 1465
rect 8666 1391 8668 1400
rect 8720 1391 8722 1400
rect 8668 1362 8720 1368
rect 8680 1331 8708 1362
rect 8956 1222 8984 1838
rect 9048 1358 9076 3606
rect 9324 3534 9352 5034
rect 9416 4622 9444 5034
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9416 4214 9444 4558
rect 9508 4282 9536 5170
rect 9600 4486 9628 7262
rect 9692 6322 9720 7822
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 6798 9904 7278
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 6390 9904 6734
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9680 5908 9732 5914
rect 9784 5896 9812 6054
rect 9732 5868 9812 5896
rect 9680 5850 9732 5856
rect 9876 5370 9904 6122
rect 9968 5710 9996 6938
rect 10060 6118 10088 7890
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7478 10272 7686
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10152 6798 10180 7346
rect 10336 6866 10364 8366
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7546 10456 7686
rect 10520 7546 10548 8230
rect 10612 7818 10640 9930
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10704 9110 10732 9862
rect 10796 9625 10824 9930
rect 10782 9616 10838 9625
rect 10782 9551 10838 9560
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10796 8974 10824 9318
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10692 8492 10744 8498
rect 10796 8480 10824 8910
rect 10744 8452 10824 8480
rect 10692 8434 10744 8440
rect 10796 8090 10824 8452
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10428 7002 10456 7210
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6458 10364 6598
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10428 6390 10456 6666
rect 10416 6384 10468 6390
rect 10414 6352 10416 6361
rect 10468 6352 10470 6361
rect 10140 6316 10192 6322
rect 10192 6276 10272 6304
rect 10414 6287 10470 6296
rect 10140 6258 10192 6264
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 3194 9352 3470
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9232 1562 9260 2314
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9220 1352 9272 1358
rect 9324 1340 9352 2858
rect 9402 2408 9458 2417
rect 9402 2343 9458 2352
rect 9416 1358 9444 2343
rect 9600 2106 9628 4422
rect 9784 4282 9812 4490
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9772 4072 9824 4078
rect 9876 4060 9904 5170
rect 9824 4032 9904 4060
rect 9772 4014 9824 4020
rect 9968 3738 9996 5238
rect 10060 5098 10088 5646
rect 10244 5574 10272 6276
rect 10428 6254 10456 6287
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 6118 10548 6190
rect 10612 6186 10640 7346
rect 10796 6458 10824 7822
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10888 6225 10916 10390
rect 10980 10130 11008 10678
rect 11058 10639 11114 10648
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10441 11100 10474
rect 11164 10470 11192 10746
rect 11152 10464 11204 10470
rect 11058 10432 11114 10441
rect 11152 10406 11204 10412
rect 11058 10367 11114 10376
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 11256 9654 11284 11494
rect 11348 11234 11376 12310
rect 11532 12238 11560 13194
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11520 12232 11572 12238
rect 11426 12200 11482 12209
rect 11520 12174 11572 12180
rect 11426 12135 11482 12144
rect 11440 12050 11468 12135
rect 11440 12022 11560 12050
rect 11532 11898 11560 12022
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11440 11370 11468 11834
rect 11520 11756 11572 11762
rect 11572 11716 11652 11744
rect 11520 11698 11572 11704
rect 11440 11354 11560 11370
rect 11440 11348 11572 11354
rect 11440 11342 11520 11348
rect 11520 11290 11572 11296
rect 11348 11206 11560 11234
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11348 10810 11376 10950
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11440 10577 11468 10746
rect 11426 10568 11482 10577
rect 11336 10532 11388 10538
rect 11426 10503 11482 10512
rect 11336 10474 11388 10480
rect 11348 9874 11376 10474
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11440 10169 11468 10406
rect 11426 10160 11482 10169
rect 11426 10095 11482 10104
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11440 9897 11468 9930
rect 11426 9888 11482 9897
rect 11348 9846 11426 9874
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11072 8974 11100 9590
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11164 9110 11192 9386
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10966 8664 11022 8673
rect 10966 8599 10968 8608
rect 11020 8599 11022 8608
rect 10968 8570 11020 8576
rect 10980 8498 11008 8570
rect 11072 8537 11100 8910
rect 11058 8528 11114 8537
rect 10968 8492 11020 8498
rect 11058 8463 11114 8472
rect 10968 8434 11020 8440
rect 11072 8294 11100 8463
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10980 7002 11008 7890
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10980 6390 11008 6938
rect 11072 6934 11100 7822
rect 11164 7750 11192 9046
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11256 8022 11284 8978
rect 11348 8974 11376 9846
rect 11426 9823 11482 9832
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11440 9489 11468 9522
rect 11426 9480 11482 9489
rect 11426 9415 11482 9424
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11348 7410 11376 7890
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10874 6216 10930 6225
rect 10600 6180 10652 6186
rect 10874 6151 10930 6160
rect 10600 6122 10652 6128
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5302 10272 5510
rect 10336 5370 10364 5714
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10232 5296 10284 5302
rect 10232 5238 10284 5244
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 10060 3890 10088 5034
rect 10336 4826 10364 5102
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10230 4584 10286 4593
rect 10230 4519 10232 4528
rect 10284 4519 10286 4528
rect 10232 4490 10284 4496
rect 10428 4282 10456 5510
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10796 4146 10824 4626
rect 11072 4282 11100 6666
rect 11440 6390 11468 9415
rect 11532 8129 11560 11206
rect 11624 10062 11652 11716
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11518 8120 11574 8129
rect 11518 8055 11574 8064
rect 11520 7880 11572 7886
rect 11624 7868 11652 9590
rect 11716 9586 11744 12242
rect 11900 12238 11928 12854
rect 12084 12434 12112 14200
rect 12214 13628 12522 13637
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13563 12522 13572
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12176 12850 12204 13262
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12636 12918 12664 13194
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12214 12540 12522 12549
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12475 12522 12484
rect 12084 12406 12204 12434
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11978 11928 12034 11937
rect 11978 11863 12034 11872
rect 11992 11762 12020 11863
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11808 11082 11836 11698
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11886 11384 11942 11393
rect 11886 11319 11888 11328
rect 11940 11319 11942 11328
rect 11888 11290 11940 11296
rect 11992 11286 12020 11494
rect 11980 11280 12032 11286
rect 11886 11248 11942 11257
rect 11980 11222 12032 11228
rect 12084 11218 12112 12038
rect 12176 11694 12204 12406
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12360 11626 12388 12106
rect 12820 11762 12848 13262
rect 12912 12646 12940 13262
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12214 11452 12522 11461
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11387 12522 11396
rect 13004 11218 13032 14334
rect 13174 14200 13230 14334
rect 14370 14200 14426 15000
rect 14384 13938 14412 14200
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12238 13216 13126
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13280 11626 13308 13194
rect 13372 12986 13400 13738
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13372 12434 13400 12922
rect 13372 12406 13492 12434
rect 13464 12170 13492 12406
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13464 11762 13492 12106
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 11886 11183 11942 11192
rect 12072 11212 12124 11218
rect 11900 11150 11928 11183
rect 12992 11212 13044 11218
rect 12124 11172 12204 11200
rect 12072 11154 12124 11160
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 11808 10470 11836 11018
rect 11978 10840 12034 10849
rect 11978 10775 12034 10784
rect 11992 10674 12020 10775
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12084 10606 12112 11018
rect 12176 10742 12204 11172
rect 12992 11154 13044 11160
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12636 10674 12664 11086
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11702 8936 11758 8945
rect 11702 8871 11758 8880
rect 11716 8362 11744 8871
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11900 8129 11928 8434
rect 11886 8120 11942 8129
rect 11886 8055 11942 8064
rect 11992 8022 12020 10066
rect 12084 8906 12112 10542
rect 13004 10418 13032 11154
rect 13280 11150 13308 11562
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13096 10538 13124 11018
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10674 13400 10950
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13176 10464 13228 10470
rect 13004 10390 13124 10418
rect 13176 10406 13228 10412
rect 12214 10364 12522 10373
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10299 12522 10308
rect 12716 10056 12768 10062
rect 12452 10004 12716 10010
rect 12452 9998 12768 10004
rect 12452 9982 12756 9998
rect 12900 9988 12952 9994
rect 12452 9926 12480 9982
rect 12900 9930 12952 9936
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12214 9276 12522 9285
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9211 12522 9220
rect 12636 8974 12664 9318
rect 12820 9178 12848 9454
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12084 8480 12112 8842
rect 12544 8498 12572 8842
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12532 8492 12584 8498
rect 12084 8452 12204 8480
rect 12176 8362 12204 8452
rect 12532 8434 12584 8440
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12084 8072 12112 8298
rect 12214 8188 12522 8197
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8123 12522 8132
rect 12084 8044 12204 8072
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11572 7840 11652 7868
rect 11704 7880 11756 7886
rect 11520 7822 11572 7828
rect 11704 7822 11756 7828
rect 11716 7546 11744 7822
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11716 7342 11744 7482
rect 11900 7410 11928 7754
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11886 7304 11942 7313
rect 11886 7239 11942 7248
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11624 7002 11652 7142
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 11256 4826 11284 5238
rect 11532 5234 11560 6258
rect 11716 5302 11744 6258
rect 11808 5302 11836 6598
rect 11900 6458 11928 7239
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11256 4282 11284 4762
rect 11808 4690 11836 5238
rect 11900 5234 11928 6258
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 10060 3862 10180 3890
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10060 3398 10088 3674
rect 10152 3602 10180 3862
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10428 3126 10456 3402
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9588 2100 9640 2106
rect 9588 2042 9640 2048
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9692 1426 9720 1974
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 9968 1358 9996 2790
rect 10428 2106 10456 3062
rect 10796 2938 10824 3402
rect 10980 3058 11008 3674
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 3126 11192 3334
rect 11256 3126 11284 4082
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11348 3602 11376 4014
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10796 2922 10916 2938
rect 10796 2916 10928 2922
rect 10796 2910 10876 2916
rect 10796 2292 10824 2910
rect 10876 2858 10928 2864
rect 10980 2650 11008 2994
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 10968 2304 11020 2310
rect 10796 2264 10968 2292
rect 10968 2246 11020 2252
rect 10416 2100 10468 2106
rect 10416 2042 10468 2048
rect 9272 1312 9352 1340
rect 9404 1352 9456 1358
rect 9220 1294 9272 1300
rect 9404 1294 9456 1300
rect 9956 1352 10008 1358
rect 9956 1294 10008 1300
rect 10980 1290 11008 2246
rect 11072 2106 11100 2314
rect 11256 2106 11284 2926
rect 11348 2582 11376 3538
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 11348 1970 11376 2518
rect 11440 2106 11468 3062
rect 11532 3058 11560 3878
rect 11900 3126 11928 4150
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11532 2666 11560 2994
rect 11532 2650 11744 2666
rect 11532 2644 11756 2650
rect 11532 2638 11704 2644
rect 11428 2100 11480 2106
rect 11428 2042 11480 2048
rect 11244 1964 11296 1970
rect 11244 1906 11296 1912
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11060 1896 11112 1902
rect 11060 1838 11112 1844
rect 11256 1850 11284 1906
rect 11440 1850 11468 2042
rect 11072 1358 11100 1838
rect 11152 1828 11204 1834
rect 11152 1770 11204 1776
rect 11256 1822 11468 1850
rect 11060 1352 11112 1358
rect 11060 1294 11112 1300
rect 10968 1284 11020 1290
rect 10968 1226 11020 1232
rect 11164 1222 11192 1770
rect 11256 1426 11284 1822
rect 11244 1420 11296 1426
rect 11244 1362 11296 1368
rect 11532 1358 11560 2638
rect 11704 2586 11756 2592
rect 11796 2032 11848 2038
rect 11796 1974 11848 1980
rect 11888 2032 11940 2038
rect 11888 1974 11940 1980
rect 11808 1426 11836 1974
rect 11796 1420 11848 1426
rect 11796 1362 11848 1368
rect 11900 1358 11928 1974
rect 11520 1352 11572 1358
rect 11520 1294 11572 1300
rect 11888 1352 11940 1358
rect 11992 1329 12020 7958
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12084 7342 12112 7754
rect 12176 7410 12204 8044
rect 12728 7886 12756 8570
rect 12820 8498 12848 9114
rect 12912 8566 12940 9930
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12624 7744 12676 7750
rect 12820 7732 12848 8298
rect 12624 7686 12676 7692
rect 12728 7704 12848 7732
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12072 7336 12124 7342
rect 12532 7336 12584 7342
rect 12072 7278 12124 7284
rect 12530 7304 12532 7313
rect 12584 7304 12586 7313
rect 12084 6984 12112 7278
rect 12530 7239 12586 7248
rect 12214 7100 12522 7109
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7035 12522 7044
rect 12636 7002 12664 7686
rect 12624 6996 12676 7002
rect 12084 6956 12204 6984
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12084 5778 12112 6802
rect 12176 6662 12204 6956
rect 12624 6938 12676 6944
rect 12728 6798 12756 7704
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12438 6352 12494 6361
rect 12438 6287 12440 6296
rect 12492 6287 12494 6296
rect 12440 6258 12492 6264
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12214 6012 12522 6021
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5947 12522 5956
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12084 5370 12112 5578
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12544 5030 12572 5850
rect 12636 5166 12664 6054
rect 12728 5914 12756 6734
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12820 5710 12848 7210
rect 12912 6458 12940 8366
rect 13096 8022 13124 10390
rect 13188 10266 13216 10406
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 8430 13216 9386
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13004 7342 13032 7822
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13004 6866 13032 7278
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 13188 6866 13216 7210
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13280 6662 13308 9454
rect 13372 8514 13400 10610
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 8634 13492 9318
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13372 8498 13492 8514
rect 13372 8492 13504 8498
rect 13372 8486 13452 8492
rect 13452 8434 13504 8440
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 6730 13400 7686
rect 13464 6798 13492 8434
rect 13556 7206 13584 8842
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12808 5704 12860 5710
rect 12728 5652 12808 5658
rect 12728 5646 12860 5652
rect 12728 5630 12848 5646
rect 12728 5234 12756 5630
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12214 4924 12522 4933
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4859 12522 4868
rect 12214 3836 12522 3845
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3771 12522 3780
rect 12636 3738 12664 4966
rect 12728 4622 12756 5034
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12532 3392 12584 3398
rect 12584 3340 12664 3346
rect 12532 3334 12664 3340
rect 12544 3318 12664 3334
rect 12636 3058 12664 3318
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12214 2748 12522 2757
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2683 12522 2692
rect 12214 1660 12522 1669
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1595 12522 1604
rect 12636 1358 12664 2994
rect 12728 2310 12756 3470
rect 12820 3466 12848 5510
rect 12912 3534 12940 6122
rect 13096 5794 13124 6598
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13004 5778 13124 5794
rect 12992 5772 13124 5778
rect 13044 5766 13124 5772
rect 12992 5714 13044 5720
rect 13004 5234 13032 5714
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13004 3670 13032 5170
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 13096 3534 13124 5102
rect 13188 4010 13216 6258
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13280 5234 13308 5510
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 13188 3398 13216 3946
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13280 3058 13308 4694
rect 13372 4622 13400 6666
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13464 3194 13492 4014
rect 13556 3777 13584 7142
rect 13648 6390 13676 11018
rect 13740 10713 13768 13126
rect 13726 10704 13782 10713
rect 13726 10639 13782 10648
rect 13740 8809 13768 10639
rect 13726 8800 13782 8809
rect 13726 8735 13782 8744
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 6458 13768 8230
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13740 4554 13768 6394
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13542 3768 13598 3777
rect 13542 3703 13598 3712
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 13096 2106 13124 2382
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 13280 2106 13308 2314
rect 13084 2100 13136 2106
rect 13084 2042 13136 2048
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 12624 1352 12676 1358
rect 11888 1294 11940 1300
rect 11978 1320 12034 1329
rect 12624 1294 12676 1300
rect 11978 1255 12034 1264
rect 8576 1216 8628 1222
rect 8576 1158 8628 1164
rect 8944 1216 8996 1222
rect 8944 1158 8996 1164
rect 11152 1216 11204 1222
rect 11152 1158 11204 1164
rect 8214 1116 8522 1125
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1051 8522 1060
rect 11164 800 11192 1158
rect 2778 504 2834 513
rect 2778 439 2834 448
rect 3698 0 3754 800
rect 11150 0 11206 800
<< via2 >>
rect 1398 12552 1454 12608
rect 1398 11620 1454 11656
rect 1398 11600 1400 11620
rect 1400 11600 1452 11620
rect 1452 11600 1454 11620
rect 3330 14456 3386 14512
rect 3514 13524 3570 13560
rect 3514 13504 3516 13524
rect 3516 13504 3568 13524
rect 3568 13504 3570 13524
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 3330 10668 3386 10704
rect 3698 10920 3754 10976
rect 3330 10648 3332 10668
rect 3332 10648 3384 10668
rect 3384 10648 3386 10668
rect 3146 9968 3202 10024
rect 3238 9696 3294 9752
rect 3606 9696 3662 9752
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 5262 11600 5318 11656
rect 4894 11056 4950 11112
rect 4802 10920 4858 10976
rect 5262 10920 5318 10976
rect 6090 12164 6146 12200
rect 6090 12144 6092 12164
rect 6092 12144 6144 12164
rect 6144 12144 6146 12164
rect 5906 12008 5962 12064
rect 6918 12280 6974 12336
rect 5814 10668 5870 10704
rect 5814 10648 5816 10668
rect 5816 10648 5868 10668
rect 5868 10648 5870 10668
rect 5906 10512 5962 10568
rect 4710 9288 4766 9344
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3790 8744 3846 8800
rect 1582 6024 1638 6080
rect 2502 7928 2558 7984
rect 3238 7928 3294 7984
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 6366 11192 6422 11248
rect 7102 12008 7158 12064
rect 7102 11736 7158 11792
rect 8850 13368 8906 13424
rect 7378 11464 7434 11520
rect 7194 11328 7250 11384
rect 4802 7928 4858 7984
rect 2870 6976 2926 7032
rect 6826 9444 6882 9480
rect 6826 9424 6828 9444
rect 6828 9424 6880 9444
rect 6880 9424 6882 9444
rect 7562 11056 7618 11112
rect 7470 10648 7526 10704
rect 7286 10240 7342 10296
rect 7378 9560 7434 9616
rect 7010 9152 7066 9208
rect 7286 9016 7342 9072
rect 7746 11464 7802 11520
rect 7746 10648 7802 10704
rect 8022 11056 8078 11112
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2042 5108 2044 5128
rect 2044 5108 2096 5128
rect 2096 5108 2098 5128
rect 2042 5072 2098 5108
rect 1490 4156 1492 4176
rect 1492 4156 1544 4176
rect 1544 4156 1546 4176
rect 1490 4120 1546 4156
rect 3514 5072 3570 5128
rect 2410 4392 2466 4448
rect 1582 2216 1638 2272
rect 3514 4120 3570 4176
rect 2686 3168 2742 3224
rect 3606 4004 3662 4040
rect 3606 3984 3608 4004
rect 3608 3984 3660 4004
rect 3660 3984 3662 4004
rect 2870 1264 2926 1320
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4434 4428 4436 4448
rect 4436 4428 4488 4448
rect 4488 4428 4490 4448
rect 4434 4392 4490 4428
rect 6918 8064 6974 8120
rect 7562 7928 7618 7984
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4618 3052 4674 3088
rect 4618 3032 4620 3052
rect 4620 3032 4672 3052
rect 4672 3032 4674 3052
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4710 2352 4766 2408
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 4802 1400 4858 1456
rect 5630 2760 5686 2816
rect 6274 4392 6330 4448
rect 5814 2760 5870 2816
rect 6826 3984 6882 4040
rect 6642 3032 6698 3088
rect 7838 9016 7894 9072
rect 8666 10376 8722 10432
rect 8574 10140 8576 10160
rect 8576 10140 8628 10160
rect 8628 10140 8630 10160
rect 8574 10104 8630 10140
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8206 9288 8262 9344
rect 8114 9152 8170 9208
rect 8298 9016 8354 9072
rect 8390 8880 8446 8936
rect 8574 9424 8630 9480
rect 9126 11464 9182 11520
rect 9310 11328 9366 11384
rect 8942 11192 8998 11248
rect 9126 10956 9128 10976
rect 9128 10956 9180 10976
rect 9180 10956 9182 10976
rect 9126 10920 9182 10956
rect 9218 10784 9274 10840
rect 8942 10548 8944 10568
rect 8944 10548 8996 10568
rect 8996 10548 8998 10568
rect 8942 10512 8998 10548
rect 9126 10512 9182 10568
rect 9034 10376 9090 10432
rect 9770 11872 9826 11928
rect 9678 11328 9734 11384
rect 10322 12316 10324 12336
rect 10324 12316 10376 12336
rect 10376 12316 10378 12336
rect 10322 12280 10378 12316
rect 10690 12436 10746 12472
rect 10690 12416 10692 12436
rect 10692 12416 10744 12436
rect 10744 12416 10746 12436
rect 10506 12280 10562 12336
rect 10230 11772 10232 11792
rect 10232 11772 10284 11792
rect 10284 11772 10286 11792
rect 10230 11736 10286 11772
rect 9678 11076 9734 11112
rect 9678 11056 9680 11076
rect 9680 11056 9732 11076
rect 9732 11056 9734 11076
rect 9494 10784 9550 10840
rect 9678 10920 9734 10976
rect 9218 10240 9274 10296
rect 8942 9716 8998 9752
rect 8942 9696 8944 9716
rect 8944 9696 8996 9716
rect 8996 9696 8998 9716
rect 10230 11192 10286 11248
rect 10690 12180 10692 12200
rect 10692 12180 10744 12200
rect 10744 12180 10746 12200
rect 10690 12144 10746 12180
rect 10046 10920 10102 10976
rect 9770 10376 9826 10432
rect 9586 10104 9642 10160
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 9034 9288 9090 9344
rect 9494 9968 9550 10024
rect 9126 9152 9182 9208
rect 9402 9152 9458 9208
rect 8942 8880 8998 8936
rect 8850 8780 8852 8800
rect 8852 8780 8904 8800
rect 8904 8780 8906 8800
rect 8850 8744 8906 8780
rect 8850 8608 8906 8664
rect 8942 8064 8998 8120
rect 9034 7964 9036 7984
rect 9036 7964 9088 7984
rect 9088 7964 9090 7984
rect 9034 7928 9090 7964
rect 9310 8880 9366 8936
rect 9586 9580 9642 9616
rect 9862 10240 9918 10296
rect 9586 9560 9588 9580
rect 9588 9560 9640 9580
rect 9640 9560 9642 9580
rect 9678 9460 9680 9480
rect 9680 9460 9732 9480
rect 9732 9460 9734 9480
rect 9494 8744 9550 8800
rect 9310 8492 9366 8528
rect 9310 8472 9312 8492
rect 9312 8472 9364 8492
rect 9364 8472 9366 8492
rect 9678 9424 9734 9460
rect 9678 8880 9734 8936
rect 10046 10512 10102 10568
rect 10046 9172 10102 9208
rect 10046 9152 10048 9172
rect 10048 9152 10100 9172
rect 10100 9152 10102 9172
rect 10322 11056 10378 11112
rect 10690 10668 10746 10704
rect 10690 10648 10692 10668
rect 10692 10648 10744 10668
rect 10744 10648 10746 10668
rect 10966 12280 11022 12336
rect 10874 11056 10930 11112
rect 10966 10920 11022 10976
rect 10874 10648 10930 10704
rect 11242 11600 11298 11656
rect 10690 10240 10746 10296
rect 10414 9696 10470 9752
rect 10322 8880 10378 8936
rect 10506 9288 10562 9344
rect 10230 8336 10286 8392
rect 8666 4548 8722 4584
rect 8666 4528 8668 4548
rect 8668 4528 8720 4548
rect 8720 4528 8722 4548
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8390 2388 8392 2408
rect 8392 2388 8444 2408
rect 8444 2388 8446 2408
rect 8390 2352 8446 2388
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 8666 1420 8722 1456
rect 8666 1400 8668 1420
rect 8668 1400 8720 1420
rect 8720 1400 8722 1420
rect 10782 9560 10838 9616
rect 10414 6332 10416 6352
rect 10416 6332 10468 6352
rect 10468 6332 10470 6352
rect 10414 6296 10470 6332
rect 9402 2352 9458 2408
rect 11058 10648 11114 10704
rect 11058 10376 11114 10432
rect 11426 12144 11482 12200
rect 11426 10512 11482 10568
rect 11426 10104 11482 10160
rect 10966 8628 11022 8664
rect 10966 8608 10968 8628
rect 10968 8608 11020 8628
rect 11020 8608 11022 8628
rect 11058 8472 11114 8528
rect 11426 9832 11482 9888
rect 11426 9424 11482 9480
rect 10874 6160 10930 6216
rect 10230 4548 10286 4584
rect 10230 4528 10232 4548
rect 10232 4528 10284 4548
rect 10284 4528 10286 4548
rect 11518 8064 11574 8120
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 11978 11872 12034 11928
rect 11886 11348 11942 11384
rect 11886 11328 11888 11348
rect 11888 11328 11940 11348
rect 11940 11328 11942 11348
rect 11886 11192 11942 11248
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 11978 10784 12034 10840
rect 11702 8880 11758 8936
rect 11886 8064 11942 8120
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 11886 7248 11942 7304
rect 12530 7284 12532 7304
rect 12532 7284 12584 7304
rect 12584 7284 12586 7304
rect 12530 7248 12586 7284
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 12438 6316 12494 6352
rect 12438 6296 12440 6316
rect 12440 6296 12492 6316
rect 12492 6296 12494 6316
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 13726 10648 13782 10704
rect 13726 8744 13782 8800
rect 13542 3712 13598 3768
rect 11978 1264 12034 1320
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 2778 448 2834 504
<< metal3 >>
rect 0 14514 800 14544
rect 3325 14514 3391 14517
rect 0 14512 3391 14514
rect 0 14456 3330 14512
rect 3386 14456 3391 14512
rect 0 14454 3391 14456
rect 0 14424 800 14454
rect 3325 14451 3391 14454
rect 14200 13698 15000 13728
rect 12758 13638 15000 13698
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 12210 13632 12526 13633
rect 12210 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12526 13632
rect 12210 13567 12526 13568
rect 3509 13562 3575 13565
rect 0 13560 3575 13562
rect 0 13504 3514 13560
rect 3570 13504 3575 13560
rect 0 13502 3575 13504
rect 0 13472 800 13502
rect 3509 13499 3575 13502
rect 8845 13426 8911 13429
rect 12758 13426 12818 13638
rect 14200 13608 15000 13638
rect 8845 13424 12818 13426
rect 8845 13368 8850 13424
rect 8906 13368 12818 13424
rect 8845 13366 12818 13368
rect 8845 13363 8911 13366
rect 8210 13088 8526 13089
rect 8210 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8526 13088
rect 8210 13023 8526 13024
rect 0 12610 800 12640
rect 1393 12610 1459 12613
rect 0 12608 1459 12610
rect 0 12552 1398 12608
rect 1454 12552 1459 12608
rect 0 12550 1459 12552
rect 0 12520 800 12550
rect 1393 12547 1459 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12210 12544 12526 12545
rect 12210 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12526 12544
rect 12210 12479 12526 12480
rect 9438 12412 9444 12476
rect 9508 12474 9514 12476
rect 10685 12474 10751 12477
rect 9508 12472 10751 12474
rect 9508 12416 10690 12472
rect 10746 12416 10751 12472
rect 9508 12414 10751 12416
rect 9508 12412 9514 12414
rect 10685 12411 10751 12414
rect 6913 12338 6979 12341
rect 10317 12338 10383 12341
rect 6913 12336 10383 12338
rect 6913 12280 6918 12336
rect 6974 12280 10322 12336
rect 10378 12280 10383 12336
rect 6913 12278 10383 12280
rect 6913 12275 6979 12278
rect 10317 12275 10383 12278
rect 10501 12338 10567 12341
rect 10961 12338 11027 12341
rect 10501 12336 11027 12338
rect 10501 12280 10506 12336
rect 10562 12280 10966 12336
rect 11022 12280 11027 12336
rect 10501 12278 11027 12280
rect 10501 12275 10567 12278
rect 10961 12275 11027 12278
rect 6085 12202 6151 12205
rect 8702 12202 8708 12204
rect 6085 12200 8708 12202
rect 6085 12144 6090 12200
rect 6146 12144 8708 12200
rect 6085 12142 8708 12144
rect 6085 12139 6151 12142
rect 8702 12140 8708 12142
rect 8772 12202 8778 12204
rect 10685 12202 10751 12205
rect 11421 12202 11487 12205
rect 8772 12200 11487 12202
rect 8772 12144 10690 12200
rect 10746 12144 11426 12200
rect 11482 12144 11487 12200
rect 8772 12142 11487 12144
rect 8772 12140 8778 12142
rect 10685 12139 10751 12142
rect 11421 12139 11487 12142
rect 5901 12066 5967 12069
rect 7097 12066 7163 12069
rect 5901 12064 7163 12066
rect 5901 12008 5906 12064
rect 5962 12008 7102 12064
rect 7158 12008 7163 12064
rect 5901 12006 7163 12008
rect 5901 12003 5967 12006
rect 7097 12003 7163 12006
rect 8210 12000 8526 12001
rect 8210 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8526 12000
rect 8210 11935 8526 11936
rect 9765 11930 9831 11933
rect 11973 11930 12039 11933
rect 9765 11928 12039 11930
rect 9765 11872 9770 11928
rect 9826 11872 11978 11928
rect 12034 11872 12039 11928
rect 9765 11870 12039 11872
rect 9765 11867 9831 11870
rect 11973 11867 12039 11870
rect 7097 11794 7163 11797
rect 10225 11796 10291 11797
rect 10174 11794 10180 11796
rect 7097 11792 10180 11794
rect 10244 11792 10291 11796
rect 7097 11736 7102 11792
rect 7158 11736 10180 11792
rect 10286 11736 10291 11792
rect 7097 11734 10180 11736
rect 7097 11731 7163 11734
rect 10174 11732 10180 11734
rect 10244 11732 10291 11736
rect 10225 11731 10291 11732
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 5257 11658 5323 11661
rect 11237 11658 11303 11661
rect 5257 11656 11303 11658
rect 5257 11600 5262 11656
rect 5318 11600 11242 11656
rect 11298 11600 11303 11656
rect 5257 11598 11303 11600
rect 5257 11595 5323 11598
rect 11237 11595 11303 11598
rect 7373 11522 7439 11525
rect 7741 11522 7807 11525
rect 9121 11522 9187 11525
rect 7373 11520 9187 11522
rect 7373 11464 7378 11520
rect 7434 11464 7746 11520
rect 7802 11464 9126 11520
rect 9182 11464 9187 11520
rect 7373 11462 9187 11464
rect 7373 11459 7439 11462
rect 7741 11459 7807 11462
rect 9121 11459 9187 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 12210 11456 12526 11457
rect 12210 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12526 11456
rect 12210 11391 12526 11392
rect 7189 11386 7255 11389
rect 9305 11386 9371 11389
rect 7189 11384 9371 11386
rect 7189 11328 7194 11384
rect 7250 11328 9310 11384
rect 9366 11328 9371 11384
rect 7189 11326 9371 11328
rect 7189 11323 7255 11326
rect 9305 11323 9371 11326
rect 9673 11386 9739 11389
rect 11881 11386 11947 11389
rect 9673 11384 11947 11386
rect 9673 11328 9678 11384
rect 9734 11328 11886 11384
rect 11942 11328 11947 11384
rect 9673 11326 11947 11328
rect 9673 11323 9739 11326
rect 11881 11323 11947 11326
rect 6361 11250 6427 11253
rect 8937 11250 9003 11253
rect 6361 11248 9003 11250
rect 6361 11192 6366 11248
rect 6422 11192 8942 11248
rect 8998 11192 9003 11248
rect 6361 11190 9003 11192
rect 6361 11187 6427 11190
rect 8937 11187 9003 11190
rect 10225 11250 10291 11253
rect 11881 11250 11947 11253
rect 14200 11250 15000 11280
rect 10225 11248 11947 11250
rect 10225 11192 10230 11248
rect 10286 11192 11886 11248
rect 11942 11192 11947 11248
rect 10225 11190 11947 11192
rect 10225 11187 10291 11190
rect 11881 11187 11947 11190
rect 12022 11190 15000 11250
rect 4889 11114 4955 11117
rect 7557 11114 7623 11117
rect 4889 11112 7623 11114
rect 4889 11056 4894 11112
rect 4950 11056 7562 11112
rect 7618 11056 7623 11112
rect 4889 11054 7623 11056
rect 4889 11051 4955 11054
rect 7557 11051 7623 11054
rect 8017 11114 8083 11117
rect 9673 11114 9739 11117
rect 8017 11112 9739 11114
rect 8017 11056 8022 11112
rect 8078 11056 9678 11112
rect 9734 11056 9739 11112
rect 8017 11054 9739 11056
rect 8017 11051 8083 11054
rect 9673 11051 9739 11054
rect 10317 11114 10383 11117
rect 10869 11114 10935 11117
rect 12022 11114 12082 11190
rect 14200 11160 15000 11190
rect 10317 11112 12082 11114
rect 10317 11056 10322 11112
rect 10378 11056 10874 11112
rect 10930 11056 12082 11112
rect 10317 11054 12082 11056
rect 10317 11051 10383 11054
rect 10869 11051 10935 11054
rect 3693 10978 3759 10981
rect 4797 10978 4863 10981
rect 5257 10978 5323 10981
rect 3693 10976 5323 10978
rect 3693 10920 3698 10976
rect 3754 10920 4802 10976
rect 4858 10920 5262 10976
rect 5318 10920 5323 10976
rect 3693 10918 5323 10920
rect 3693 10915 3759 10918
rect 4797 10915 4863 10918
rect 5257 10915 5323 10918
rect 9121 10978 9187 10981
rect 9673 10978 9739 10981
rect 9121 10976 9739 10978
rect 9121 10920 9126 10976
rect 9182 10920 9678 10976
rect 9734 10920 9739 10976
rect 9121 10918 9739 10920
rect 9121 10915 9187 10918
rect 9673 10915 9739 10918
rect 10041 10978 10107 10981
rect 10961 10978 11027 10981
rect 10041 10976 11027 10978
rect 10041 10920 10046 10976
rect 10102 10920 10966 10976
rect 11022 10920 11027 10976
rect 10041 10918 11027 10920
rect 10041 10915 10107 10918
rect 10961 10915 11027 10918
rect 8210 10912 8526 10913
rect 8210 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8526 10912
rect 8210 10847 8526 10848
rect 9213 10844 9279 10845
rect 9213 10840 9260 10844
rect 9324 10842 9330 10844
rect 9489 10842 9555 10845
rect 11973 10842 12039 10845
rect 9213 10784 9218 10840
rect 9213 10780 9260 10784
rect 9324 10782 9370 10842
rect 9489 10840 12039 10842
rect 9489 10784 9494 10840
rect 9550 10784 11978 10840
rect 12034 10784 12039 10840
rect 9489 10782 12039 10784
rect 9324 10780 9330 10782
rect 9213 10779 9279 10780
rect 9489 10779 9555 10782
rect 11973 10779 12039 10782
rect 0 10706 800 10736
rect 3325 10706 3391 10709
rect 0 10704 3391 10706
rect 0 10648 3330 10704
rect 3386 10648 3391 10704
rect 0 10646 3391 10648
rect 0 10616 800 10646
rect 3325 10643 3391 10646
rect 5809 10706 5875 10709
rect 7465 10706 7531 10709
rect 5809 10704 7531 10706
rect 5809 10648 5814 10704
rect 5870 10648 7470 10704
rect 7526 10648 7531 10704
rect 5809 10646 7531 10648
rect 5809 10643 5875 10646
rect 7465 10643 7531 10646
rect 7741 10706 7807 10709
rect 9438 10706 9444 10708
rect 7741 10704 9444 10706
rect 7741 10648 7746 10704
rect 7802 10648 9444 10704
rect 7741 10646 9444 10648
rect 7741 10643 7807 10646
rect 9438 10644 9444 10646
rect 9508 10644 9514 10708
rect 10685 10706 10751 10709
rect 10869 10706 10935 10709
rect 10685 10704 10935 10706
rect 10685 10648 10690 10704
rect 10746 10648 10874 10704
rect 10930 10648 10935 10704
rect 10685 10646 10935 10648
rect 10685 10643 10751 10646
rect 10869 10643 10935 10646
rect 11053 10706 11119 10709
rect 13721 10706 13787 10709
rect 11053 10704 13787 10706
rect 11053 10648 11058 10704
rect 11114 10648 13726 10704
rect 13782 10648 13787 10704
rect 11053 10646 13787 10648
rect 11053 10643 11119 10646
rect 13721 10643 13787 10646
rect 5901 10570 5967 10573
rect 8937 10570 9003 10573
rect 9121 10572 9187 10573
rect 5901 10568 9003 10570
rect 5901 10512 5906 10568
rect 5962 10512 8942 10568
rect 8998 10512 9003 10568
rect 5901 10510 9003 10512
rect 5901 10507 5967 10510
rect 8937 10507 9003 10510
rect 9070 10508 9076 10572
rect 9140 10570 9187 10572
rect 10041 10570 10107 10573
rect 11421 10570 11487 10573
rect 9140 10568 9232 10570
rect 9182 10512 9232 10568
rect 9140 10510 9232 10512
rect 10041 10568 11487 10570
rect 10041 10512 10046 10568
rect 10102 10512 11426 10568
rect 11482 10512 11487 10568
rect 10041 10510 11487 10512
rect 9140 10508 9187 10510
rect 9121 10507 9187 10508
rect 10041 10507 10107 10510
rect 11421 10507 11487 10510
rect 8661 10434 8727 10437
rect 9029 10434 9095 10437
rect 8661 10432 9095 10434
rect 8661 10376 8666 10432
rect 8722 10376 9034 10432
rect 9090 10376 9095 10432
rect 8661 10374 9095 10376
rect 8661 10371 8727 10374
rect 9029 10371 9095 10374
rect 9765 10434 9831 10437
rect 11053 10434 11119 10437
rect 9765 10432 11119 10434
rect 9765 10376 9770 10432
rect 9826 10376 11058 10432
rect 11114 10376 11119 10432
rect 9765 10374 11119 10376
rect 9765 10371 9831 10374
rect 11053 10371 11119 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12210 10368 12526 10369
rect 12210 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12526 10368
rect 12210 10303 12526 10304
rect 7281 10298 7347 10301
rect 9213 10298 9279 10301
rect 7281 10296 9279 10298
rect 7281 10240 7286 10296
rect 7342 10240 9218 10296
rect 9274 10240 9279 10296
rect 7281 10238 9279 10240
rect 7281 10235 7347 10238
rect 9213 10235 9279 10238
rect 9857 10298 9923 10301
rect 10685 10298 10751 10301
rect 9857 10296 10751 10298
rect 9857 10240 9862 10296
rect 9918 10240 10690 10296
rect 10746 10240 10751 10296
rect 9857 10238 10751 10240
rect 9857 10235 9923 10238
rect 10685 10235 10751 10238
rect 8569 10162 8635 10165
rect 9581 10162 9647 10165
rect 11421 10162 11487 10165
rect 8569 10160 9092 10162
rect 8569 10104 8574 10160
rect 8630 10128 9092 10160
rect 9581 10160 11487 10162
rect 8630 10104 9138 10128
rect 8569 10102 9138 10104
rect 8569 10099 8635 10102
rect 9032 10068 9138 10102
rect 9581 10104 9586 10160
rect 9642 10104 11426 10160
rect 11482 10104 11487 10160
rect 9581 10102 11487 10104
rect 9581 10099 9647 10102
rect 11421 10099 11487 10102
rect 3141 10026 3207 10029
rect 3141 10024 8954 10026
rect 3141 9968 3146 10024
rect 3202 9968 8954 10024
rect 3141 9966 8954 9968
rect 3141 9963 3207 9966
rect 8894 9890 8954 9966
rect 9078 9890 9138 10068
rect 9254 9964 9260 10028
rect 9324 10026 9330 10028
rect 9489 10026 9555 10029
rect 9324 10024 9555 10026
rect 9324 9968 9494 10024
rect 9550 9968 9555 10024
rect 9324 9966 9555 9968
rect 9324 9964 9330 9966
rect 9489 9963 9555 9966
rect 11421 9890 11487 9893
rect 8894 9830 9000 9890
rect 9078 9888 11487 9890
rect 9078 9832 11426 9888
rect 11482 9832 11487 9888
rect 9078 9830 11487 9832
rect 8210 9824 8526 9825
rect 0 9754 800 9784
rect 8210 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8526 9824
rect 8210 9759 8526 9760
rect 8940 9757 9000 9830
rect 11421 9827 11487 9830
rect 3233 9754 3299 9757
rect 3601 9754 3667 9757
rect 0 9752 3667 9754
rect 0 9696 3238 9752
rect 3294 9696 3606 9752
rect 3662 9696 3667 9752
rect 0 9694 3667 9696
rect 0 9664 800 9694
rect 3233 9691 3299 9694
rect 3601 9691 3667 9694
rect 8937 9754 9003 9757
rect 10409 9754 10475 9757
rect 8937 9752 10475 9754
rect 8937 9696 8942 9752
rect 8998 9696 10414 9752
rect 10470 9696 10475 9752
rect 8937 9694 10475 9696
rect 8937 9691 9003 9694
rect 10409 9691 10475 9694
rect 7373 9618 7439 9621
rect 9581 9618 9647 9621
rect 10777 9618 10843 9621
rect 7373 9616 10843 9618
rect 7373 9560 7378 9616
rect 7434 9560 9586 9616
rect 9642 9560 10782 9616
rect 10838 9560 10843 9616
rect 7373 9558 10843 9560
rect 7373 9555 7439 9558
rect 9581 9555 9647 9558
rect 10777 9555 10843 9558
rect 6821 9482 6887 9485
rect 8569 9482 8635 9485
rect 6821 9480 8635 9482
rect 6821 9424 6826 9480
rect 6882 9424 8574 9480
rect 8630 9424 8635 9480
rect 6821 9422 8635 9424
rect 6821 9419 6887 9422
rect 8569 9419 8635 9422
rect 9673 9482 9739 9485
rect 11421 9482 11487 9485
rect 9673 9480 11487 9482
rect 9673 9424 9678 9480
rect 9734 9424 11426 9480
rect 11482 9424 11487 9480
rect 9673 9422 11487 9424
rect 9673 9419 9739 9422
rect 11421 9419 11487 9422
rect 4705 9346 4771 9349
rect 8201 9346 8267 9349
rect 4705 9344 8267 9346
rect 4705 9288 4710 9344
rect 4766 9288 8206 9344
rect 8262 9288 8267 9344
rect 4705 9286 8267 9288
rect 4705 9283 4771 9286
rect 8201 9283 8267 9286
rect 9029 9346 9095 9349
rect 10501 9346 10567 9349
rect 9029 9344 10567 9346
rect 9029 9288 9034 9344
rect 9090 9288 10506 9344
rect 10562 9288 10567 9344
rect 9029 9286 10567 9288
rect 9029 9283 9095 9286
rect 10501 9283 10567 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12210 9280 12526 9281
rect 12210 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12526 9280
rect 12210 9215 12526 9216
rect 7005 9210 7071 9213
rect 8109 9210 8175 9213
rect 7005 9208 8175 9210
rect 7005 9152 7010 9208
rect 7066 9152 8114 9208
rect 8170 9152 8175 9208
rect 7005 9150 8175 9152
rect 7005 9147 7071 9150
rect 8109 9147 8175 9150
rect 9121 9208 9187 9213
rect 9121 9152 9126 9208
rect 9182 9152 9187 9208
rect 9121 9147 9187 9152
rect 9397 9210 9463 9213
rect 10041 9210 10107 9213
rect 9397 9208 10107 9210
rect 9397 9152 9402 9208
rect 9458 9152 10046 9208
rect 10102 9152 10107 9208
rect 9397 9150 10107 9152
rect 9397 9147 9463 9150
rect 10041 9147 10107 9150
rect 7281 9074 7347 9077
rect 7833 9074 7899 9077
rect 8293 9074 8359 9077
rect 8702 9074 8708 9076
rect 7281 9072 8708 9074
rect 7281 9016 7286 9072
rect 7342 9016 7838 9072
rect 7894 9016 8298 9072
rect 8354 9016 8708 9072
rect 7281 9014 8708 9016
rect 7281 9011 7347 9014
rect 7833 9011 7899 9014
rect 8293 9011 8359 9014
rect 8702 9012 8708 9014
rect 8772 9012 8778 9076
rect 9124 9074 9184 9147
rect 9124 9014 9368 9074
rect 9308 8941 9368 9014
rect 8385 8938 8451 8941
rect 8937 8938 9003 8941
rect 8385 8936 9003 8938
rect 8385 8880 8390 8936
rect 8446 8880 8942 8936
rect 8998 8880 9003 8936
rect 8385 8878 9003 8880
rect 8385 8875 8451 8878
rect 8937 8875 9003 8878
rect 9305 8936 9371 8941
rect 9305 8880 9310 8936
rect 9366 8880 9371 8936
rect 9305 8875 9371 8880
rect 9673 8938 9739 8941
rect 10317 8938 10383 8941
rect 11697 8938 11763 8941
rect 9673 8936 11763 8938
rect 9673 8880 9678 8936
rect 9734 8880 10322 8936
rect 10378 8880 11702 8936
rect 11758 8880 11763 8936
rect 9673 8878 11763 8880
rect 9673 8875 9739 8878
rect 10317 8875 10383 8878
rect 11697 8875 11763 8878
rect 0 8802 800 8832
rect 3785 8802 3851 8805
rect 0 8800 3851 8802
rect 0 8744 3790 8800
rect 3846 8744 3851 8800
rect 0 8742 3851 8744
rect 0 8712 800 8742
rect 3785 8739 3851 8742
rect 8845 8802 8911 8805
rect 9070 8802 9076 8804
rect 8845 8800 9076 8802
rect 8845 8744 8850 8800
rect 8906 8744 9076 8800
rect 8845 8742 9076 8744
rect 8845 8739 8911 8742
rect 9070 8740 9076 8742
rect 9140 8802 9146 8804
rect 9489 8802 9555 8805
rect 9140 8800 9555 8802
rect 9140 8744 9494 8800
rect 9550 8744 9555 8800
rect 9140 8742 9555 8744
rect 9140 8740 9146 8742
rect 9489 8739 9555 8742
rect 13721 8802 13787 8805
rect 14200 8802 15000 8832
rect 13721 8800 15000 8802
rect 13721 8744 13726 8800
rect 13782 8744 15000 8800
rect 13721 8742 15000 8744
rect 13721 8739 13787 8742
rect 8210 8736 8526 8737
rect 8210 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8526 8736
rect 14200 8712 15000 8742
rect 8210 8671 8526 8672
rect 8845 8666 8911 8669
rect 10961 8666 11027 8669
rect 8845 8664 11027 8666
rect 8845 8608 8850 8664
rect 8906 8608 10966 8664
rect 11022 8608 11027 8664
rect 8845 8606 11027 8608
rect 8845 8603 8911 8606
rect 10961 8603 11027 8606
rect 9305 8530 9371 8533
rect 11053 8530 11119 8533
rect 9305 8528 11119 8530
rect 9305 8472 9310 8528
rect 9366 8472 11058 8528
rect 11114 8472 11119 8528
rect 9305 8470 11119 8472
rect 9305 8467 9371 8470
rect 11053 8467 11119 8470
rect 10225 8396 10291 8397
rect 10174 8332 10180 8396
rect 10244 8394 10291 8396
rect 10244 8392 10336 8394
rect 10286 8336 10336 8392
rect 10244 8334 10336 8336
rect 10244 8332 10291 8334
rect 10225 8331 10291 8332
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 12210 8192 12526 8193
rect 12210 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12526 8192
rect 12210 8127 12526 8128
rect 6913 8122 6979 8125
rect 8937 8122 9003 8125
rect 11513 8122 11579 8125
rect 11881 8122 11947 8125
rect 6913 8120 11947 8122
rect 6913 8064 6918 8120
rect 6974 8064 8942 8120
rect 8998 8064 11518 8120
rect 11574 8064 11886 8120
rect 11942 8064 11947 8120
rect 6913 8062 11947 8064
rect 6913 8059 6979 8062
rect 8937 8059 9003 8062
rect 11513 8059 11579 8062
rect 11881 8059 11947 8062
rect 0 7986 800 8016
rect 2497 7986 2563 7989
rect 3233 7986 3299 7989
rect 0 7984 3299 7986
rect 0 7928 2502 7984
rect 2558 7928 3238 7984
rect 3294 7928 3299 7984
rect 0 7926 3299 7928
rect 0 7896 800 7926
rect 2497 7923 2563 7926
rect 3233 7923 3299 7926
rect 4797 7986 4863 7989
rect 7557 7986 7623 7989
rect 9029 7986 9095 7989
rect 4797 7984 9095 7986
rect 4797 7928 4802 7984
rect 4858 7928 7562 7984
rect 7618 7928 9034 7984
rect 9090 7928 9095 7984
rect 4797 7926 9095 7928
rect 4797 7923 4863 7926
rect 7557 7923 7623 7926
rect 9029 7923 9095 7926
rect 8210 7648 8526 7649
rect 8210 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8526 7648
rect 8210 7583 8526 7584
rect 11881 7306 11947 7309
rect 12525 7306 12591 7309
rect 11881 7304 12591 7306
rect 11881 7248 11886 7304
rect 11942 7248 12530 7304
rect 12586 7248 12591 7304
rect 11881 7246 12591 7248
rect 11881 7243 11947 7246
rect 12525 7243 12591 7246
rect 4210 7104 4526 7105
rect 0 7034 800 7064
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12210 7104 12526 7105
rect 12210 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12526 7104
rect 12210 7039 12526 7040
rect 2865 7034 2931 7037
rect 0 7032 2931 7034
rect 0 6976 2870 7032
rect 2926 6976 2931 7032
rect 0 6974 2931 6976
rect 0 6944 800 6974
rect 2865 6971 2931 6974
rect 8210 6560 8526 6561
rect 8210 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8526 6560
rect 8210 6495 8526 6496
rect 10409 6354 10475 6357
rect 12433 6354 12499 6357
rect 10409 6352 12499 6354
rect 10409 6296 10414 6352
rect 10470 6296 12438 6352
rect 12494 6296 12499 6352
rect 10409 6294 12499 6296
rect 10409 6291 10475 6294
rect 12433 6291 12499 6294
rect 10869 6218 10935 6221
rect 14200 6218 15000 6248
rect 10869 6216 15000 6218
rect 10869 6160 10874 6216
rect 10930 6160 15000 6216
rect 10869 6158 15000 6160
rect 10869 6155 10935 6158
rect 14200 6128 15000 6158
rect 0 6082 800 6112
rect 1577 6082 1643 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 800 6022
rect 1577 6019 1643 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12210 6016 12526 6017
rect 12210 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12526 6016
rect 12210 5951 12526 5952
rect 8210 5472 8526 5473
rect 8210 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8526 5472
rect 8210 5407 8526 5408
rect 0 5130 800 5160
rect 2037 5130 2103 5133
rect 3509 5130 3575 5133
rect 0 5128 3575 5130
rect 0 5072 2042 5128
rect 2098 5072 3514 5128
rect 3570 5072 3575 5128
rect 0 5070 3575 5072
rect 0 5040 800 5070
rect 2037 5067 2103 5070
rect 3509 5067 3575 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12210 4928 12526 4929
rect 12210 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12526 4928
rect 12210 4863 12526 4864
rect 8661 4586 8727 4589
rect 10225 4586 10291 4589
rect 8661 4584 10291 4586
rect 8661 4528 8666 4584
rect 8722 4528 10230 4584
rect 10286 4528 10291 4584
rect 8661 4526 10291 4528
rect 8661 4523 8727 4526
rect 10225 4523 10291 4526
rect 2405 4450 2471 4453
rect 4429 4450 4495 4453
rect 6269 4450 6335 4453
rect 2405 4448 6335 4450
rect 2405 4392 2410 4448
rect 2466 4392 4434 4448
rect 4490 4392 6274 4448
rect 6330 4392 6335 4448
rect 2405 4390 6335 4392
rect 2405 4387 2471 4390
rect 4429 4387 4495 4390
rect 6269 4387 6335 4390
rect 8210 4384 8526 4385
rect 8210 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8526 4384
rect 8210 4319 8526 4320
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 3509 4178 3575 4181
rect 0 4176 3575 4178
rect 0 4120 1490 4176
rect 1546 4120 3514 4176
rect 3570 4120 3575 4176
rect 0 4118 3575 4120
rect 0 4088 800 4118
rect 1485 4115 1551 4118
rect 3509 4115 3575 4118
rect 3601 4042 3667 4045
rect 6821 4042 6887 4045
rect 3601 4040 6887 4042
rect 3601 3984 3606 4040
rect 3662 3984 6826 4040
rect 6882 3984 6887 4040
rect 3601 3982 6887 3984
rect 3601 3979 3667 3982
rect 6821 3979 6887 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12210 3840 12526 3841
rect 12210 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12526 3840
rect 12210 3775 12526 3776
rect 13537 3770 13603 3773
rect 14200 3770 15000 3800
rect 13537 3768 15000 3770
rect 13537 3712 13542 3768
rect 13598 3712 15000 3768
rect 13537 3710 15000 3712
rect 13537 3707 13603 3710
rect 14200 3680 15000 3710
rect 8210 3296 8526 3297
rect 0 3226 800 3256
rect 8210 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8526 3296
rect 8210 3231 8526 3232
rect 2681 3226 2747 3229
rect 0 3224 2747 3226
rect 0 3168 2686 3224
rect 2742 3168 2747 3224
rect 0 3166 2747 3168
rect 0 3136 800 3166
rect 2681 3163 2747 3166
rect 4613 3090 4679 3093
rect 6637 3090 6703 3093
rect 4613 3088 6703 3090
rect 4613 3032 4618 3088
rect 4674 3032 6642 3088
rect 6698 3032 6703 3088
rect 4613 3030 6703 3032
rect 4613 3027 4679 3030
rect 6637 3027 6703 3030
rect 5625 2818 5691 2821
rect 5809 2818 5875 2821
rect 5625 2816 5875 2818
rect 5625 2760 5630 2816
rect 5686 2760 5814 2816
rect 5870 2760 5875 2816
rect 5625 2758 5875 2760
rect 5625 2755 5691 2758
rect 5809 2755 5875 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12210 2752 12526 2753
rect 12210 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12526 2752
rect 12210 2687 12526 2688
rect 4705 2410 4771 2413
rect 8385 2410 8451 2413
rect 9397 2410 9463 2413
rect 4705 2408 9463 2410
rect 4705 2352 4710 2408
rect 4766 2352 8390 2408
rect 8446 2352 9402 2408
rect 9458 2352 9463 2408
rect 4705 2350 9463 2352
rect 4705 2347 4771 2350
rect 8385 2347 8451 2350
rect 9397 2347 9463 2350
rect 0 2274 800 2304
rect 1577 2274 1643 2277
rect 0 2272 1643 2274
rect 0 2216 1582 2272
rect 1638 2216 1643 2272
rect 0 2214 1643 2216
rect 0 2184 800 2214
rect 1577 2211 1643 2214
rect 8210 2208 8526 2209
rect 8210 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8526 2208
rect 8210 2143 8526 2144
rect 4210 1664 4526 1665
rect 4210 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4526 1664
rect 4210 1599 4526 1600
rect 12210 1664 12526 1665
rect 12210 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12526 1664
rect 12210 1599 12526 1600
rect 4797 1458 4863 1461
rect 8661 1458 8727 1461
rect 4797 1456 8727 1458
rect 4797 1400 4802 1456
rect 4858 1400 8666 1456
rect 8722 1400 8727 1456
rect 4797 1398 8727 1400
rect 4797 1395 4863 1398
rect 8661 1395 8727 1398
rect 0 1322 800 1352
rect 2865 1322 2931 1325
rect 0 1320 2931 1322
rect 0 1264 2870 1320
rect 2926 1264 2931 1320
rect 0 1262 2931 1264
rect 0 1232 800 1262
rect 2865 1259 2931 1262
rect 11973 1322 12039 1325
rect 14200 1322 15000 1352
rect 11973 1320 15000 1322
rect 11973 1264 11978 1320
rect 12034 1264 15000 1320
rect 11973 1262 15000 1264
rect 11973 1259 12039 1262
rect 14200 1232 15000 1262
rect 8210 1120 8526 1121
rect 8210 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8526 1120
rect 8210 1055 8526 1056
rect 0 506 800 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 800 446
rect 2773 443 2839 446
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 9444 12412 9508 12476
rect 8708 12140 8772 12204
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 10180 11792 10244 11796
rect 10180 11736 10230 11792
rect 10230 11736 10244 11792
rect 10180 11732 10244 11736
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 9260 10840 9324 10844
rect 9260 10784 9274 10840
rect 9274 10784 9324 10840
rect 9260 10780 9324 10784
rect 9444 10644 9508 10708
rect 9076 10568 9140 10572
rect 9076 10512 9126 10568
rect 9126 10512 9140 10568
rect 9076 10508 9140 10512
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 9260 9964 9324 10028
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 8708 9012 8772 9076
rect 9076 8740 9140 8804
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 10180 8392 10244 8396
rect 10180 8336 10230 8392
rect 10230 8336 10244 8392
rect 10180 8332 10244 8336
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12488 4296 12544
rect 4360 12488 4376 12544
rect 4440 12488 4456 12544
rect 4520 12480 4528 12544
rect 4208 12252 4250 12480
rect 4486 12252 4528 12480
rect 4208 11456 4528 12252
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4488 4528 4864
rect 4208 4252 4250 4488
rect 4486 4252 4528 4488
rect 4208 3840 4528 4252
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12488 12296 12544
rect 12360 12488 12376 12544
rect 12440 12488 12456 12544
rect 12520 12480 12528 12544
rect 9443 12476 9509 12477
rect 9443 12412 9444 12476
rect 9508 12412 9509 12476
rect 9443 12411 9509 12412
rect 8707 12204 8773 12205
rect 8707 12140 8708 12204
rect 8772 12140 8773 12204
rect 8707 12139 8773 12140
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8710 9077 8770 12139
rect 9259 10844 9325 10845
rect 9259 10780 9260 10844
rect 9324 10780 9325 10844
rect 9259 10779 9325 10780
rect 9075 10572 9141 10573
rect 9075 10508 9076 10572
rect 9140 10508 9141 10572
rect 9075 10507 9141 10508
rect 8707 9076 8773 9077
rect 8707 9012 8708 9076
rect 8772 9012 8773 9076
rect 8707 9011 8773 9012
rect 9078 8805 9138 10507
rect 9262 10029 9322 10779
rect 9446 10709 9506 12411
rect 12208 12252 12250 12480
rect 12486 12252 12528 12480
rect 10179 11796 10245 11797
rect 10179 11732 10180 11796
rect 10244 11732 10245 11796
rect 10179 11731 10245 11732
rect 9443 10708 9509 10709
rect 9443 10644 9444 10708
rect 9508 10644 9509 10708
rect 9443 10643 9509 10644
rect 9259 10028 9325 10029
rect 9259 9964 9260 10028
rect 9324 9964 9325 10028
rect 9259 9963 9325 9964
rect 9075 8804 9141 8805
rect 9075 8740 9076 8804
rect 9140 8740 9141 8804
rect 9075 8739 9141 8740
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 8488 8528 8672
rect 8208 8252 8250 8488
rect 8486 8252 8528 8488
rect 10182 8397 10242 11731
rect 12208 11456 12528 12252
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 10179 8396 10245 8397
rect 10179 8332 10180 8396
rect 10244 8332 10245 8396
rect 10179 8331 10245 8332
rect 8208 7648 8528 8252
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 4488 12528 4864
rect 12208 4252 12250 4488
rect 12486 4252 12528 4488
rect 12208 3840 12528 4252
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
<< via4 >>
rect 4250 12480 4280 12488
rect 4280 12480 4296 12488
rect 4296 12480 4360 12488
rect 4360 12480 4376 12488
rect 4376 12480 4440 12488
rect 4440 12480 4456 12488
rect 4456 12480 4486 12488
rect 4250 12252 4486 12480
rect 4250 4252 4486 4488
rect 12250 12480 12280 12488
rect 12280 12480 12296 12488
rect 12296 12480 12360 12488
rect 12360 12480 12376 12488
rect 12376 12480 12440 12488
rect 12440 12480 12456 12488
rect 12456 12480 12486 12488
rect 12250 12252 12486 12480
rect 8250 8252 8486 8488
rect 12250 4252 12486 4488
<< metal5 >>
rect 1056 12488 13940 12530
rect 1056 12252 4250 12488
rect 4486 12252 12250 12488
rect 12486 12252 13940 12488
rect 1056 12210 13940 12252
rect 1056 8488 13940 8530
rect 1056 8252 8250 8488
rect 8486 8252 13940 8488
rect 1056 8210 13940 8252
rect 1056 4488 13940 4530
rect 1056 4252 4250 4488
rect 4486 4252 12250 4488
rect 12486 4252 13940 4488
rect 1056 4210 13940 4252
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 1564 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A1
timestamp 1665323087
transform -1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__B2
timestamp 1665323087
transform -1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A1
timestamp 1665323087
transform 1 0 1472 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B1
timestamp 1665323087
transform 1 0 1472 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__B1
timestamp 1665323087
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1665323087
transform -1 0 3680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__B1
timestamp 1665323087
transform -1 0 3680 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__B1
timestamp 1665323087
transform -1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A1
timestamp 1665323087
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1665323087
transform -1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1665323087
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1665323087
transform 1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A1
timestamp 1665323087
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A_N
timestamp 1665323087
transform -1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A2
timestamp 1665323087
transform -1 0 3680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1665323087
transform -1 0 2668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A2
timestamp 1665323087
transform -1 0 4784 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A2
timestamp 1665323087
transform -1 0 1564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A2
timestamp 1665323087
transform -1 0 1564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A2
timestamp 1665323087
transform -1 0 3680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A2
timestamp 1665323087
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A2
timestamp 1665323087
transform -1 0 3956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A2
timestamp 1665323087
transform 1 0 4416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A2
timestamp 1665323087
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1665323087
transform 1 0 3864 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1665323087
transform 1 0 7360 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__B1
timestamp 1665323087
transform 1 0 5704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A2
timestamp 1665323087
transform -1 0 6624 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A2
timestamp 1665323087
transform -1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A2
timestamp 1665323087
transform -1 0 7728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__B
timestamp 1665323087
transform -1 0 11408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__B1
timestamp 1665323087
transform -1 0 11408 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A2
timestamp 1665323087
transform -1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__B1
timestamp 1665323087
transform -1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A2
timestamp 1665323087
transform -1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A2
timestamp 1665323087
transform -1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__B1
timestamp 1665323087
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A2
timestamp 1665323087
transform -1 0 10764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__B1
timestamp 1665323087
transform -1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A2
timestamp 1665323087
transform -1 0 12512 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A2
timestamp 1665323087
transform 1 0 13432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A2
timestamp 1665323087
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1665323087
transform -1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__B
timestamp 1665323087
transform -1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__D
timestamp 1665323087
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1665323087
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8096 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1665323087
transform 1 0 8648 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10120 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118
timestamp 1665323087
transform 1 0 11960 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13248 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1665323087
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_79 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8372 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1665323087
transform 1 0 13432 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_132
timestamp 1665323087
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1665323087
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1665323087
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1665323087
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_118
timestamp 1665323087
transform 1 0 11960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1665323087
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1665323087
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_62
timestamp 1665323087
transform 1 0 6808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_78
timestamp 1665323087
transform 1 0 8280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_94
timestamp 1665323087
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_101
timestamp 1665323087
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp 1665323087
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1665323087
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_48
timestamp 1665323087
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp 1665323087
transform 1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_91
timestamp 1665323087
transform 1 0 9476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_105
timestamp 1665323087
transform 1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1665323087
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_67
timestamp 1665323087
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1665323087
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1665323087
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_112
timestamp 1665323087
transform 1 0 11408 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_122
timestamp 1665323087
transform 1 0 12328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1665323087
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_64
timestamp 1665323087
transform 1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_88
timestamp 1665323087
transform 1 0 9200 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1665323087
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp 1665323087
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1665323087
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_77
timestamp 1665323087
transform 1 0 8188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1665323087
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1665323087
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1665323087
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_84
timestamp 1665323087
transform 1 0 8832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_52
timestamp 1665323087
transform 1 0 5888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1665323087
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1665323087
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_135
timestamp 1665323087
transform 1 0 13524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1665323087
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_14
timestamp 1665323087
transform 1 0 2392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_105
timestamp 1665323087
transform 1 0 10764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1665323087
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_41
timestamp 1665323087
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_135
timestamp 1665323087
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_50
timestamp 1665323087
transform 1 0 5704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1665323087
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_84
timestamp 1665323087
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1665323087
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1665323087
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_26
timestamp 1665323087
transform 1 0 3496 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_51
timestamp 1665323087
transform 1 0 5796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_125
timestamp 1665323087
transform 1 0 12604 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1665323087
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1665323087
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_112
timestamp 1665323087
transform 1 0 11408 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_69
timestamp 1665323087
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_86
timestamp 1665323087
transform 1 0 9016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1665323087
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_80
timestamp 1665323087
transform 1 0 8464 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_20
timestamp 1665323087
transform 1 0 2944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_50
timestamp 1665323087
transform 1 0 5704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1665323087
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_79
timestamp 1665323087
transform 1 0 8372 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1665323087
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1665323087
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_106
timestamp 1665323087
transform 1 0 10856 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_135
timestamp 1665323087
transform 1 0 13524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1665323087
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_17
timestamp 1665323087
transform 1 0 2668 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1665323087
transform 1 0 8004 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1665323087
transform 1 0 13524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1665323087
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1665323087
transform 1 0 4968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1665323087
transform 1 0 5704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1665323087
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_98
timestamp 1665323087
transform 1 0 10120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1665323087
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1665323087
transform -1 0 13892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1665323087
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1665323087
transform -1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1665323087
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1665323087
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1665323087
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1665323087
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1665323087
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1665323087
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1665323087
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1665323087
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1665323087
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1665323087
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1665323087
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1665323087
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1665323087
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1665323087
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1665323087
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1665323087
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1665323087
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1665323087
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1665323087
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1665323087
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1665323087
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1665323087
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1665323087
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1665323087
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1665323087
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1665323087
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1665323087
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1665323087
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1665323087
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1665323087
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1665323087
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1665323087
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1665323087
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1665323087
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1665323087
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1665323087
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1665323087
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1665323087
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1665323087
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1665323087
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1665323087
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1665323087
transform -1 0 13892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1665323087
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1665323087
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1665323087
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1665323087
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1665323087
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1665323087
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1665323087
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1665323087
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1665323087
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1665323087
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1665323087
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1665323087
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1665323087
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1665323087
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1665323087
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1665323087
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1665323087
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1665323087
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1665323087
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1665323087
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1665323087
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1665323087
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1665323087
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1665323087
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1665323087
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1665323087
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1665323087
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1665323087
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1665323087
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1665323087
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1665323087
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1665323087
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1665323087
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1665323087
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1665323087
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1665323087
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1665323087
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1665323087
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1665323087
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1665323087
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1665323087
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1665323087
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1665323087
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1665323087
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1665323087
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1665323087
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1665323087
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1665323087
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1665323087
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_2  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 13248 0 1 1088
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6256 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2392 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _212_
timestamp 1665323087
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _213_
timestamp 1665323087
transform 1 0 3312 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _214_
timestamp 1665323087
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _215_
timestamp 1665323087
transform -1 0 5520 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _216_
timestamp 1665323087
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _217_
timestamp 1665323087
transform 1 0 3772 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _218_
timestamp 1665323087
transform -1 0 3588 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _219_
timestamp 1665323087
transform -1 0 6808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _220_
timestamp 1665323087
transform 1 0 6808 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _221_
timestamp 1665323087
transform -1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _222_
timestamp 1665323087
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _223_
timestamp 1665323087
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 6992 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3772 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _227_
timestamp 1665323087
transform -1 0 4968 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3680 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _229_
timestamp 1665323087
transform -1 0 7912 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 7360 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _231_
timestamp 1665323087
transform -1 0 8004 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2024 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _233_
timestamp 1665323087
transform -1 0 2024 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _234_
timestamp 1665323087
transform -1 0 5980 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _235_
timestamp 1665323087
transform -1 0 5520 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _236_
timestamp 1665323087
transform -1 0 3772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3864 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4968 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _239_
timestamp 1665323087
transform -1 0 4324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _240_
timestamp 1665323087
transform -1 0 2024 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2668 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _243_
timestamp 1665323087
transform -1 0 5244 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _244_
timestamp 1665323087
transform 1 0 4968 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _245_
timestamp 1665323087
transform 1 0 6440 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _246_
timestamp 1665323087
transform -1 0 4508 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_2  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1932 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2668 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _249_
timestamp 1665323087
transform -1 0 3220 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_2  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _251_
timestamp 1665323087
transform -1 0 2300 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _252_
timestamp 1665323087
transform -1 0 1932 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _253_
timestamp 1665323087
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1665323087
transform -1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3312 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _256_
timestamp 1665323087
transform 1 0 2300 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _257_
timestamp 1665323087
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3312 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _259_
timestamp 1665323087
transform 1 0 2208 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _260_
timestamp 1665323087
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _261_
timestamp 1665323087
transform -1 0 1840 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1932 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3496 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _264_
timestamp 1665323087
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1665323087
transform -1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _266_
timestamp 1665323087
transform 1 0 13248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1665323087
transform -1 0 11408 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _268_
timestamp 1665323087
transform -1 0 11132 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _269_
timestamp 1665323087
transform -1 0 8464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _271_
timestamp 1665323087
transform -1 0 8004 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _272_
timestamp 1665323087
transform -1 0 12880 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _273_
timestamp 1665323087
transform -1 0 10580 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _274_
timestamp 1665323087
transform 1 0 7912 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_2  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8556 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_2  _276_
timestamp 1665323087
transform -1 0 13248 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_2  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 10396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1656 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _279_
timestamp 1665323087
transform 1 0 1472 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2852 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _281_
timestamp 1665323087
transform 1 0 2760 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9292 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _283_
timestamp 1665323087
transform 1 0 10028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _284_
timestamp 1665323087
transform 1 0 10120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _285_
timestamp 1665323087
transform 1 0 12328 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _286_
timestamp 1665323087
transform -1 0 13248 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _287_
timestamp 1665323087
transform 1 0 12236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _288_
timestamp 1665323087
transform 1 0 12880 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _289_
timestamp 1665323087
transform -1 0 7912 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1665323087
transform -1 0 9568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _291_
timestamp 1665323087
transform 1 0 7636 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _292_
timestamp 1665323087
transform 1 0 11500 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_2  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9844 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _294_
timestamp 1665323087
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_2  _295_
timestamp 1665323087
transform 1 0 8280 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_2  _296_
timestamp 1665323087
transform 1 0 12420 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _297_
timestamp 1665323087
transform -1 0 13432 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _298_
timestamp 1665323087
transform -1 0 11408 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11500 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _300_
timestamp 1665323087
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _301_
timestamp 1665323087
transform -1 0 13248 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _302_
timestamp 1665323087
transform -1 0 13616 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _303_
timestamp 1665323087
transform -1 0 12328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _304_
timestamp 1665323087
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _305_
timestamp 1665323087
transform -1 0 13616 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _306_
timestamp 1665323087
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _307_
timestamp 1665323087
transform -1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1665323087
transform -1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _309_
timestamp 1665323087
transform 1 0 10580 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _310_
timestamp 1665323087
transform 1 0 10212 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _311_
timestamp 1665323087
transform -1 0 10028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _312_
timestamp 1665323087
transform 1 0 6164 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _313_
timestamp 1665323087
transform 1 0 8924 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o2bb2a_2  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9016 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _315_
timestamp 1665323087
transform -1 0 8832 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _316_
timestamp 1665323087
transform 1 0 9292 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_2  _317_
timestamp 1665323087
transform 1 0 9936 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _318_
timestamp 1665323087
transform -1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _319_
timestamp 1665323087
transform -1 0 9476 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _320_
timestamp 1665323087
transform 1 0 10028 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _321_
timestamp 1665323087
transform -1 0 6624 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _322_
timestamp 1665323087
transform -1 0 6164 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _323_
timestamp 1665323087
transform 1 0 4324 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _324_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 5612 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _325_
timestamp 1665323087
transform 1 0 4692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _326_
timestamp 1665323087
transform 1 0 5336 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _327_
timestamp 1665323087
transform 1 0 5428 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _328_
timestamp 1665323087
transform 1 0 5980 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _329_
timestamp 1665323087
transform 1 0 5612 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _330_
timestamp 1665323087
transform 1 0 5060 0 1 1088
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _331_
timestamp 1665323087
transform 1 0 6348 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _332_
timestamp 1665323087
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _333_
timestamp 1665323087
transform 1 0 9936 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _334_
timestamp 1665323087
transform -1 0 10120 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _335_
timestamp 1665323087
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _336_
timestamp 1665323087
transform -1 0 8648 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _337_
timestamp 1665323087
transform -1 0 11224 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _338_
timestamp 1665323087
transform -1 0 9292 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _339_
timestamp 1665323087
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _340_
timestamp 1665323087
transform -1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _341_
timestamp 1665323087
transform -1 0 8832 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _342_
timestamp 1665323087
transform 1 0 4232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _343_
timestamp 1665323087
transform 1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _344_
timestamp 1665323087
transform -1 0 10212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _345_
timestamp 1665323087
transform -1 0 11040 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _346_
timestamp 1665323087
transform -1 0 10120 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _347_
timestamp 1665323087
transform -1 0 6256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_2  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6992 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _349_
timestamp 1665323087
transform -1 0 6256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _350_
timestamp 1665323087
transform -1 0 6716 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _351_
timestamp 1665323087
transform -1 0 3680 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _352_
timestamp 1665323087
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _353_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _354_
timestamp 1665323087
transform -1 0 3036 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _355_
timestamp 1665323087
transform -1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_2  _356_
timestamp 1665323087
transform 1 0 6532 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _357_
timestamp 1665323087
transform -1 0 2208 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _358_
timestamp 1665323087
transform -1 0 6164 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _359_
timestamp 1665323087
transform 1 0 6624 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _360_
timestamp 1665323087
transform 1 0 2852 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _361_
timestamp 1665323087
transform -1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _362_
timestamp 1665323087
transform -1 0 4968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _363_
timestamp 1665323087
transform -1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _364_
timestamp 1665323087
transform -1 0 5888 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _365_
timestamp 1665323087
transform 1 0 4968 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _366_
timestamp 1665323087
transform -1 0 5704 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _367_
timestamp 1665323087
transform 1 0 11960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _368_
timestamp 1665323087
transform 1 0 8280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _369_
timestamp 1665323087
transform -1 0 8280 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _370_
timestamp 1665323087
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _371_
timestamp 1665323087
transform 1 0 7452 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_2  _372_
timestamp 1665323087
transform 1 0 8464 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _373_
timestamp 1665323087
transform -1 0 9844 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _374_
timestamp 1665323087
transform -1 0 7452 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _375_
timestamp 1665323087
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _376_
timestamp 1665323087
transform -1 0 6256 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _377_
timestamp 1665323087
transform 1 0 5888 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _378_
timestamp 1665323087
transform 1 0 5888 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _379_
timestamp 1665323087
transform 1 0 6624 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _380_
timestamp 1665323087
transform 1 0 8924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _381_
timestamp 1665323087
transform 1 0 8188 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _382_
timestamp 1665323087
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _383_
timestamp 1665323087
transform -1 0 8464 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _384_
timestamp 1665323087
transform -1 0 11224 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _385_
timestamp 1665323087
transform 1 0 10672 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _386_
timestamp 1665323087
transform 1 0 9384 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _387_
timestamp 1665323087
transform -1 0 10304 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _388_
timestamp 1665323087
transform -1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _389_
timestamp 1665323087
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _390_
timestamp 1665323087
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _391_
timestamp 1665323087
transform 1 0 10028 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _392_
timestamp 1665323087
transform 1 0 13156 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _393_
timestamp 1665323087
transform -1 0 11868 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _394_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 9108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _395_
timestamp 1665323087
transform 1 0 9476 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _396_
timestamp 1665323087
transform 1 0 9936 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _397_
timestamp 1665323087
transform 1 0 10304 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _398_
timestamp 1665323087
transform 1 0 11868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _399_
timestamp 1665323087
transform -1 0 9660 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _400_
timestamp 1665323087
transform 1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _401_
timestamp 1665323087
transform 1 0 7544 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _402_
timestamp 1665323087
transform 1 0 7912 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _403_
timestamp 1665323087
transform -1 0 8372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _404_
timestamp 1665323087
transform 1 0 7268 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _405_
timestamp 1665323087
transform 1 0 8740 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _406_
timestamp 1665323087
transform 1 0 10212 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _407_
timestamp 1665323087
transform 1 0 7544 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _408_
timestamp 1665323087
transform 1 0 10304 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _409_
timestamp 1665323087
transform -1 0 11224 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _410_
timestamp 1665323087
transform -1 0 11960 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_2  _411_
timestamp 1665323087
transform 1 0 10580 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _412_
timestamp 1665323087
transform 1 0 9936 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _413_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 11868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _414_
timestamp 1665323087
transform 1 0 12696 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _415_
timestamp 1665323087
transform 1 0 10672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _416_
timestamp 1665323087
transform -1 0 3312 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _417_
timestamp 1665323087
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _418_
timestamp 1665323087
transform 1 0 8372 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _419_
timestamp 1665323087
transform 1 0 8372 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _420_
timestamp 1665323087
transform 1 0 9292 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _421_
timestamp 1665323087
transform -1 0 8280 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _422_
timestamp 1665323087
transform 1 0 4600 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _423_
timestamp 1665323087
transform -1 0 7360 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _424_
timestamp 1665323087
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _425_
timestamp 1665323087
transform -1 0 7268 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _426_
timestamp 1665323087
transform -1 0 6992 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _427_
timestamp 1665323087
transform -1 0 6440 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _428_
timestamp 1665323087
transform 1 0 7728 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _429_
timestamp 1665323087
transform 1 0 8188 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _430_
timestamp 1665323087
transform 1 0 7176 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _431_
timestamp 1665323087
transform 1 0 6716 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _432_
timestamp 1665323087
transform 1 0 7728 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _433_
timestamp 1665323087
transform -1 0 10948 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _434_
timestamp 1665323087
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _435_
timestamp 1665323087
transform 1 0 11500 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _436_
timestamp 1665323087
transform 1 0 10948 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _437_
timestamp 1665323087
transform 1 0 11500 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _438_
timestamp 1665323087
transform 1 0 10948 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _439_
timestamp 1665323087
transform 1 0 12788 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _440_
timestamp 1665323087
transform -1 0 8096 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _441_
timestamp 1665323087
transform -1 0 8372 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _442_
timestamp 1665323087
transform 1 0 4600 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _443_
timestamp 1665323087
transform -1 0 4232 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _444_
timestamp 1665323087
transform -1 0 3220 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _445_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 8924 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _446_
timestamp 1665323087
transform 1 0 8004 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _447_
timestamp 1665323087
transform 1 0 8648 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _448_
timestamp 1665323087
transform 1 0 5336 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _449_
timestamp 1665323087
transform -1 0 5888 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _450_
timestamp 1665323087
transform -1 0 8280 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _451_
timestamp 1665323087
transform 1 0 5428 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _452_
timestamp 1665323087
transform 1 0 3956 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _453_
timestamp 1665323087
transform -1 0 9200 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _454_
timestamp 1665323087
transform 1 0 9476 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _455_
timestamp 1665323087
transform 1 0 6440 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _456_
timestamp 1665323087
transform -1 0 8280 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _457_
timestamp 1665323087
transform 1 0 10488 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _458_
timestamp 1665323087
transform 1 0 11500 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _459_
timestamp 1665323087
transform -1 0 12420 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _460_
timestamp 1665323087
transform 1 0 11500 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _461_
timestamp 1665323087
transform -1 0 12788 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _462_
timestamp 1665323087
transform 1 0 10488 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1665323087
transform 1 0 6440 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _464_
timestamp 1665323087
transform 1 0 2024 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _465_
timestamp 1665323087
transform -1 0 5888 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _466_
timestamp 1665323087
transform 1 0 2668 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _467_
timestamp 1665323087
transform -1 0 3312 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 3220 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_1
timestamp 1665323087
transform 1 0 1380 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 5428 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4416 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1665323087
transform -1 0 5796 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4048 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6072 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1665323087
transform -1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1665323087
transform -1 0 4232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1665323087
transform 1 0 3956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1665323087
transform -1 0 5888 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1665323087
transform 1 0 3772 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1665323087
transform -1 0 5244 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1665323087
transform 1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1665323087
transform -1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1665323087
transform -1 0 3036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1665323087
transform -1 0 3128 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1665323087
transform -1 0 4416 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1665323087
transform 1 0 1840 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1665323087
transform -1 0 3864 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1665323087
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1665323087
transform -1 0 3496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1665323087
transform -1 0 1748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1665323087
transform -1 0 2392 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1665323087
transform -1 0 2484 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1665323087
transform 1 0 1380 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1665323087
transform -1 0 2760 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1665323087
transform -1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1665323087
transform -1 0 2944 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1665323087
transform 1 0 2392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1665323087
transform 1 0 2208 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1665323087
transform 1 0 1748 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1665323087
transform 1 0 1472 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1665323087
transform 1 0 1564 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1665323087
transform -1 0 1748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1665323087
transform 1 0 3128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1665323087
transform 1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1665323087
transform 1 0 3036 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1665323087
transform 1 0 3036 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1665323087
transform 1 0 2760 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1665323087
transform -1 0 4784 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1665323087
transform 1 0 3956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1665323087
transform 1 0 3956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1665323087
transform -1 0 4140 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1665323087
transform 1 0 5060 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1665323087
transform -1 0 4968 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1665323087
transform 1 0 4600 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1665323087
transform 1 0 4140 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1665323087
transform 1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1665323087
transform 1 0 6348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1665323087
transform -1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1665323087
transform 1 0 6348 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1665323087
transform 1 0 8004 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1665323087
transform 1 0 6348 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1665323087
transform -1 0 8004 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1665323087
transform -1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1665323087
transform 1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1665323087
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1665323087
transform 1 0 9660 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1665323087
transform -1 0 10120 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1665323087
transform 1 0 8464 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1665323087
transform -1 0 11132 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1665323087
transform -1 0 9476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1665323087
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1665323087
transform -1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1665323087
transform 1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1665323087
transform -1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1665323087
transform 1 0 11500 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1665323087
transform 1 0 10948 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1665323087
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1665323087
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1665323087
transform -1 0 7268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1665323087
transform 1 0 12788 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1665323087
transform -1 0 11408 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1665323087
transform 1 0 12512 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1665323087
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1665323087
transform 1 0 13248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1665323087
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1665323087
transform 1 0 12604 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1665323087
transform 1 0 12696 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1665323087
transform 1 0 11960 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1665323087
transform 1 0 12604 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1665323087
transform -1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform -1 0 6256 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1665323087
transform -1 0 1840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1665323087
transform 1 0 1380 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1665323087
transform 1 0 12144 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1665323087
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1665323087
transform -1 0 12144 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1665323087
transform -1 0 13156 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1665323087
transform -1 0 12696 0 1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1665323087
transform -1 0 12512 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1665323087
transform -1 0 11408 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 10856 0 1 7616
box -38 -48 498 592
<< labels >>
flabel metal4 s 8208 1040 8528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8210 13940 8530 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 1040 4528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12208 1040 12528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4210 13940 4530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12210 13940 12530 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 416 800 536 0 FreeSans 480 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 1232 800 1352 0 FreeSans 480 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 3974 14200 4030 15000 0 FreeSans 224 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 5170 14200 5226 15000 0 FreeSans 224 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 6274 14200 6330 15000 0 FreeSans 224 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 7470 14200 7526 15000 0 FreeSans 224 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 8574 14200 8630 15000 0 FreeSans 224 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 9770 14200 9826 15000 0 FreeSans 224 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 10874 14200 10930 15000 0 FreeSans 224 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 12070 14200 12126 15000 0 FreeSans 224 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 13174 14200 13230 15000 0 FreeSans 224 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 14370 14200 14426 15000 0 FreeSans 224 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 14200 13608 15000 13728 0 FreeSans 480 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 14200 11160 15000 11280 0 FreeSans 480 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 14200 8712 15000 8832 0 FreeSans 480 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 14200 6128 15000 6248 0 FreeSans 480 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 14200 3680 15000 3800 0 FreeSans 480 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 14200 1232 15000 1352 0 FreeSans 480 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 570 14200 626 15000 0 FreeSans 224 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 1674 14200 1730 15000 0 FreeSans 224 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 2870 14200 2926 15000 0 FreeSans 224 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15000 15000
<< end >>
