magic
tech sky130A
magscale 1 2
timestamp 1677512547
<< viali >>
rect 1869 8585 1903 8619
rect 4445 8585 4479 8619
rect 4997 8517 5031 8551
rect 2421 8449 2455 8483
rect 6469 8449 6503 8483
rect 3249 8381 3283 8415
rect 5825 8381 5859 8415
rect 7297 8381 7331 8415
rect 3985 8313 4019 8347
rect 1961 8041 1995 8075
rect 6745 8041 6779 8075
rect 2421 7837 2455 7871
rect 3985 7837 4019 7871
rect 5365 7837 5399 7871
rect 3249 7769 3283 7803
rect 4813 7769 4847 7803
rect 6193 7769 6227 7803
rect 7297 7701 7331 7735
rect 1685 7497 1719 7531
rect 3065 7429 3099 7463
rect 4997 7429 5031 7463
rect 6469 7429 6503 7463
rect 2237 7361 2271 7395
rect 3617 7361 3651 7395
rect 4445 7361 4479 7395
rect 5733 7293 5767 7327
rect 7297 7293 7331 7327
rect 1501 6953 1535 6987
rect 2053 6953 2087 6987
rect 5457 6749 5491 6783
rect 7297 6749 7331 6783
rect 4721 6681 4755 6715
rect 5917 6681 5951 6715
rect 6653 6681 6687 6715
rect 2789 6613 2823 6647
rect 3249 6613 3283 6647
rect 3985 6613 4019 6647
rect 5825 6409 5859 6443
rect 1777 6341 1811 6375
rect 3249 6341 3283 6375
rect 5273 6341 5307 6375
rect 6469 6341 6503 6375
rect 2605 6273 2639 6307
rect 3985 6273 4019 6307
rect 4445 6273 4479 6307
rect 7205 6205 7239 6239
rect 3249 5729 3283 5763
rect 5457 5729 5491 5763
rect 6469 5661 6503 5695
rect 1961 5593 1995 5627
rect 2421 5593 2455 5627
rect 4721 5593 4755 5627
rect 7205 5593 7239 5627
rect 4169 5525 4203 5559
rect 2697 5253 2731 5287
rect 4077 5253 4111 5287
rect 5457 5253 5491 5287
rect 7389 5253 7423 5287
rect 1961 5185 1995 5219
rect 3341 5185 3375 5219
rect 4721 5185 4755 5219
rect 6561 5117 6595 5151
rect 2513 4641 2547 4675
rect 5733 4641 5767 4675
rect 7389 4573 7423 4607
rect 3341 4505 3375 4539
rect 4905 4505 4939 4539
rect 6561 4505 6595 4539
rect 1869 4437 1903 4471
rect 4353 4437 4387 4471
rect 3709 4165 3743 4199
rect 7389 4165 7423 4199
rect 2973 4097 3007 4131
rect 4261 4097 4295 4131
rect 5089 4097 5123 4131
rect 5917 4097 5951 4131
rect 6561 4029 6595 4063
rect 2237 3961 2271 3995
rect 1777 3893 1811 3927
rect 3893 3689 3927 3723
rect 7389 3689 7423 3723
rect 6837 3621 6871 3655
rect 2605 3553 2639 3587
rect 5273 3553 5307 3587
rect 3341 3417 3375 3451
rect 4445 3417 4479 3451
rect 5917 3417 5951 3451
rect 1961 3349 1995 3383
rect 1685 3145 1719 3179
rect 6469 3145 6503 3179
rect 7389 3145 7423 3179
rect 4169 3077 4203 3111
rect 4997 3077 5031 3111
rect 2881 3009 2915 3043
rect 3617 3009 3651 3043
rect 5549 3009 5583 3043
rect 2237 2805 2271 2839
rect 1961 2601 1995 2635
rect 7205 2533 7239 2567
rect 2513 2465 2547 2499
rect 4721 2465 4755 2499
rect 5457 2465 5491 2499
rect 3341 2329 3375 2363
rect 3893 2329 3927 2363
rect 6193 2329 6227 2363
rect 6745 2261 6779 2295
rect 1593 2057 1627 2091
rect 2145 2057 2179 2091
rect 2789 1989 2823 2023
rect 6561 1989 6595 2023
rect 3525 1921 3559 1955
rect 4077 1921 4111 1955
rect 4905 1921 4939 1955
rect 7389 1921 7423 1955
rect 5457 1717 5491 1751
rect 4077 1377 4111 1411
rect 1961 1309 1995 1343
rect 3341 1309 3375 1343
rect 5917 1309 5951 1343
rect 2513 1241 2547 1275
rect 4813 1241 4847 1275
rect 5365 1241 5399 1275
rect 7389 1173 7423 1207
<< metal1 >>
rect 5626 9392 5632 9444
rect 5684 9432 5690 9444
rect 6362 9432 6368 9444
rect 5684 9404 6368 9432
rect 5684 9392 5690 9404
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 7834 9392 7840 9444
rect 7892 9432 7898 9444
rect 8294 9432 8300 9444
rect 7892 9404 8300 9432
rect 7892 9392 7898 9404
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 5534 8888 5540 8900
rect 4120 8860 5540 8888
rect 4120 8848 4126 8860
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 6638 8820 6644 8832
rect 5224 8792 6644 8820
rect 5224 8780 5230 8792
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 1012 8730 8071 8752
rect 1012 8678 2582 8730
rect 2634 8678 2646 8730
rect 2698 8678 2710 8730
rect 2762 8678 2774 8730
rect 2826 8678 2838 8730
rect 2890 8678 4307 8730
rect 4359 8678 4371 8730
rect 4423 8678 4435 8730
rect 4487 8678 4499 8730
rect 4551 8678 4563 8730
rect 4615 8678 6032 8730
rect 6084 8678 6096 8730
rect 6148 8678 6160 8730
rect 6212 8678 6224 8730
rect 6276 8678 6288 8730
rect 6340 8678 7757 8730
rect 7809 8678 7821 8730
rect 7873 8678 7885 8730
rect 7937 8678 7949 8730
rect 8001 8678 8013 8730
rect 8065 8678 8071 8730
rect 1012 8656 8071 8678
rect 1854 8616 1860 8628
rect 1815 8588 1860 8616
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 3694 8576 3700 8628
rect 3752 8616 3758 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 3752 8588 4445 8616
rect 3752 8576 3758 8588
rect 4433 8585 4445 8588
rect 4479 8616 4491 8619
rect 4706 8616 4712 8628
rect 4479 8588 4712 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 1872 8548 1900 8576
rect 4985 8551 5043 8557
rect 4985 8548 4997 8551
rect 1872 8520 4997 8548
rect 4985 8517 4997 8520
rect 5031 8517 5043 8551
rect 4985 8511 5043 8517
rect 2406 8480 2412 8492
rect 2367 8452 2412 8480
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 6457 8483 6515 8489
rect 6457 8480 6469 8483
rect 3936 8452 6469 8480
rect 3936 8440 3942 8452
rect 6457 8449 6469 8452
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 4246 8412 4252 8424
rect 3283 8384 4252 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8412 5871 8415
rect 5902 8412 5908 8424
rect 5859 8384 5908 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 8110 8412 8116 8424
rect 7331 8384 8116 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 934 8304 940 8356
rect 992 8344 998 8356
rect 1486 8344 1492 8356
rect 992 8316 1492 8344
rect 992 8304 998 8316
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 3973 8347 4031 8353
rect 3973 8344 3985 8347
rect 2372 8316 3985 8344
rect 2372 8304 2378 8316
rect 3973 8313 3985 8316
rect 4019 8344 4031 8347
rect 4062 8344 4068 8356
rect 4019 8316 4068 8344
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 1012 8186 7912 8208
rect 1012 8134 1720 8186
rect 1772 8134 1784 8186
rect 1836 8134 1848 8186
rect 1900 8134 1912 8186
rect 1964 8134 1976 8186
rect 2028 8134 3445 8186
rect 3497 8134 3509 8186
rect 3561 8134 3573 8186
rect 3625 8134 3637 8186
rect 3689 8134 3701 8186
rect 3753 8134 5170 8186
rect 5222 8134 5234 8186
rect 5286 8134 5298 8186
rect 5350 8134 5362 8186
rect 5414 8134 5426 8186
rect 5478 8134 6895 8186
rect 6947 8134 6959 8186
rect 7011 8134 7023 8186
rect 7075 8134 7087 8186
rect 7139 8134 7151 8186
rect 7203 8134 7912 8186
rect 1012 8112 7912 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2958 8072 2964 8084
rect 1995 8044 2964 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2958 8032 2964 8044
rect 3016 8072 3022 8084
rect 3878 8072 3884 8084
rect 3016 8044 3884 8072
rect 3016 8032 3022 8044
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6696 8044 6745 8072
rect 6696 8032 6702 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 4798 7964 4804 8016
rect 4856 8004 4862 8016
rect 5166 8004 5172 8016
rect 4856 7976 5172 8004
rect 4856 7964 4862 7976
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 1486 7828 1492 7880
rect 1544 7868 1550 7880
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 1544 7840 2421 7868
rect 1544 7828 1550 7840
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 2409 7831 2467 7837
rect 2746 7840 3985 7868
rect 1302 7760 1308 7812
rect 1360 7800 1366 7812
rect 2746 7800 2774 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 5353 7871 5411 7877
rect 5353 7868 5365 7871
rect 4120 7840 5365 7868
rect 4120 7828 4126 7840
rect 5353 7837 5365 7840
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 1360 7772 2774 7800
rect 3237 7803 3295 7809
rect 1360 7760 1366 7772
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 4154 7800 4160 7812
rect 3283 7772 4160 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 4154 7760 4160 7772
rect 4212 7760 4218 7812
rect 4798 7800 4804 7812
rect 4759 7772 4804 7800
rect 4798 7760 4804 7772
rect 4856 7760 4862 7812
rect 6181 7803 6239 7809
rect 6181 7769 6193 7803
rect 6227 7800 6239 7803
rect 6362 7800 6368 7812
rect 6227 7772 6368 7800
rect 6227 7769 6239 7772
rect 6181 7763 6239 7769
rect 6362 7760 6368 7772
rect 6420 7760 6426 7812
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7248 7704 7297 7732
rect 7248 7692 7254 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7285 7695 7343 7701
rect 1012 7642 8071 7664
rect 1012 7590 2582 7642
rect 2634 7590 2646 7642
rect 2698 7590 2710 7642
rect 2762 7590 2774 7642
rect 2826 7590 2838 7642
rect 2890 7590 4307 7642
rect 4359 7590 4371 7642
rect 4423 7590 4435 7642
rect 4487 7590 4499 7642
rect 4551 7590 4563 7642
rect 4615 7590 6032 7642
rect 6084 7590 6096 7642
rect 6148 7590 6160 7642
rect 6212 7590 6224 7642
rect 6276 7590 6288 7642
rect 6340 7590 7757 7642
rect 7809 7590 7821 7642
rect 7873 7590 7885 7642
rect 7937 7590 7949 7642
rect 8001 7590 8013 7642
rect 8065 7590 8071 7642
rect 1012 7568 8071 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1673 7531 1731 7537
rect 1673 7528 1685 7531
rect 1360 7500 1685 7528
rect 1360 7488 1366 7500
rect 1673 7497 1685 7500
rect 1719 7497 1731 7531
rect 5350 7528 5356 7540
rect 1673 7491 1731 7497
rect 3068 7500 5356 7528
rect 3068 7469 3096 7500
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7429 3111 7463
rect 3053 7423 3111 7429
rect 4706 7420 4712 7472
rect 4764 7460 4770 7472
rect 4985 7463 5043 7469
rect 4985 7460 4997 7463
rect 4764 7432 4997 7460
rect 4764 7420 4770 7432
rect 4985 7429 4997 7432
rect 5031 7429 5043 7463
rect 4985 7423 5043 7429
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 6457 7463 6515 7469
rect 6457 7460 6469 7463
rect 5592 7432 6469 7460
rect 5592 7420 5598 7432
rect 6457 7429 6469 7432
rect 6503 7460 6515 7463
rect 7190 7460 7196 7472
rect 6503 7432 7196 7460
rect 6503 7429 6515 7432
rect 6457 7423 6515 7429
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 7282 7420 7288 7472
rect 7340 7460 7346 7472
rect 7558 7460 7564 7472
rect 7340 7432 7564 7460
rect 7340 7420 7346 7432
rect 7558 7420 7564 7432
rect 7616 7420 7622 7472
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 3292 7364 3617 7392
rect 3292 7352 3298 7364
rect 3605 7361 3617 7364
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 6546 7392 6552 7404
rect 4479 7364 6552 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5721 7327 5779 7333
rect 5721 7324 5733 7327
rect 5592 7296 5733 7324
rect 5592 7284 5598 7296
rect 5721 7293 5733 7296
rect 5767 7293 5779 7327
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 5721 7287 5779 7293
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5166 7188 5172 7200
rect 5040 7160 5172 7188
rect 5040 7148 5046 7160
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 1012 7098 7912 7120
rect 1012 7046 1720 7098
rect 1772 7046 1784 7098
rect 1836 7046 1848 7098
rect 1900 7046 1912 7098
rect 1964 7046 1976 7098
rect 2028 7046 3445 7098
rect 3497 7046 3509 7098
rect 3561 7046 3573 7098
rect 3625 7046 3637 7098
rect 3689 7046 3701 7098
rect 3753 7046 5170 7098
rect 5222 7046 5234 7098
rect 5286 7046 5298 7098
rect 5350 7046 5362 7098
rect 5414 7046 5426 7098
rect 5478 7046 6895 7098
rect 6947 7046 6959 7098
rect 7011 7046 7023 7098
rect 7075 7046 7087 7098
rect 7139 7046 7151 7098
rect 7203 7046 7912 7098
rect 1012 7024 7912 7046
rect 1486 6984 1492 6996
rect 1447 6956 1492 6984
rect 1486 6944 1492 6956
rect 1544 6944 1550 6996
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 2041 6987 2099 6993
rect 2041 6984 2053 6987
rect 1636 6956 2053 6984
rect 1636 6944 1642 6956
rect 2041 6953 2053 6956
rect 2087 6984 2099 6987
rect 2222 6984 2228 6996
rect 2087 6956 2228 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 5718 6780 5724 6792
rect 5491 6752 5724 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 7285 6783 7343 6789
rect 7285 6780 7297 6783
rect 5920 6752 7297 6780
rect 4709 6715 4767 6721
rect 4709 6681 4721 6715
rect 4755 6681 4767 6715
rect 4709 6675 4767 6681
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 3050 6644 3056 6656
rect 2823 6616 3056 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3234 6644 3240 6656
rect 3195 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3970 6644 3976 6656
rect 3931 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4724 6644 4752 6675
rect 4982 6672 4988 6724
rect 5040 6712 5046 6724
rect 5920 6721 5948 6752
rect 7285 6749 7297 6752
rect 7331 6749 7343 6783
rect 7285 6743 7343 6749
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 5040 6684 5917 6712
rect 5040 6672 5046 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 5905 6675 5963 6681
rect 6546 6672 6552 6724
rect 6604 6712 6610 6724
rect 6641 6715 6699 6721
rect 6641 6712 6653 6715
rect 6604 6684 6653 6712
rect 6604 6672 6610 6684
rect 6641 6681 6653 6684
rect 6687 6681 6699 6715
rect 6641 6675 6699 6681
rect 4798 6644 4804 6656
rect 4724 6616 4804 6644
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 7466 6644 7472 6656
rect 5316 6616 7472 6644
rect 5316 6604 5322 6616
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 1012 6554 8071 6576
rect 1012 6502 2582 6554
rect 2634 6502 2646 6554
rect 2698 6502 2710 6554
rect 2762 6502 2774 6554
rect 2826 6502 2838 6554
rect 2890 6502 4307 6554
rect 4359 6502 4371 6554
rect 4423 6502 4435 6554
rect 4487 6502 4499 6554
rect 4551 6502 4563 6554
rect 4615 6502 6032 6554
rect 6084 6502 6096 6554
rect 6148 6502 6160 6554
rect 6212 6502 6224 6554
rect 6276 6502 6288 6554
rect 6340 6502 7757 6554
rect 7809 6502 7821 6554
rect 7873 6502 7885 6554
rect 7937 6502 7949 6554
rect 8001 6502 8013 6554
rect 8065 6502 8071 6554
rect 1012 6480 8071 6502
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5813 6443 5871 6449
rect 5813 6440 5825 6443
rect 5776 6412 5825 6440
rect 5776 6400 5782 6412
rect 5813 6409 5825 6412
rect 5859 6409 5871 6443
rect 5813 6403 5871 6409
rect 1026 6332 1032 6384
rect 1084 6372 1090 6384
rect 1765 6375 1823 6381
rect 1765 6372 1777 6375
rect 1084 6344 1777 6372
rect 1084 6332 1090 6344
rect 1765 6341 1777 6344
rect 1811 6341 1823 6375
rect 1765 6335 1823 6341
rect 3237 6375 3295 6381
rect 3237 6341 3249 6375
rect 3283 6372 3295 6375
rect 3786 6372 3792 6384
rect 3283 6344 3792 6372
rect 3283 6341 3295 6344
rect 3237 6335 3295 6341
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 5258 6372 5264 6384
rect 5219 6344 5264 6372
rect 5258 6332 5264 6344
rect 5316 6332 5322 6384
rect 6457 6375 6515 6381
rect 6457 6341 6469 6375
rect 6503 6372 6515 6375
rect 6638 6372 6644 6384
rect 6503 6344 6644 6372
rect 6503 6341 6515 6344
rect 6457 6335 6515 6341
rect 6638 6332 6644 6344
rect 6696 6332 6702 6384
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 7374 6372 7380 6384
rect 6788 6344 7380 6372
rect 6788 6332 6794 6344
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 3970 6304 3976 6316
rect 2639 6276 2774 6304
rect 3931 6276 3976 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 2746 6236 2774 6276
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4433 6307 4491 6313
rect 4433 6304 4445 6307
rect 4304 6276 4445 6304
rect 4304 6264 4310 6276
rect 4433 6273 4445 6276
rect 4479 6273 4491 6307
rect 4433 6267 4491 6273
rect 3050 6236 3056 6248
rect 2746 6208 3056 6236
rect 3050 6196 3056 6208
rect 3108 6236 3114 6248
rect 3878 6236 3884 6248
rect 3108 6208 3884 6236
rect 3108 6196 3114 6208
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6788 6208 7205 6236
rect 6788 6196 6794 6208
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 1012 6010 7912 6032
rect 1012 5958 1720 6010
rect 1772 5958 1784 6010
rect 1836 5958 1848 6010
rect 1900 5958 1912 6010
rect 1964 5958 1976 6010
rect 2028 5958 3445 6010
rect 3497 5958 3509 6010
rect 3561 5958 3573 6010
rect 3625 5958 3637 6010
rect 3689 5958 3701 6010
rect 3753 5958 5170 6010
rect 5222 5958 5234 6010
rect 5286 5958 5298 6010
rect 5350 5958 5362 6010
rect 5414 5958 5426 6010
rect 5478 5958 6895 6010
rect 6947 5958 6959 6010
rect 7011 5958 7023 6010
rect 7075 5958 7087 6010
rect 7139 5958 7151 6010
rect 7203 5958 7912 6010
rect 1012 5936 7912 5958
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 4062 5760 4068 5772
rect 3283 5732 4068 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 5442 5760 5448 5772
rect 5403 5732 5448 5760
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 3050 5692 3056 5704
rect 1452 5664 3056 5692
rect 1452 5652 1458 5664
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 5902 5652 5908 5704
rect 5960 5692 5966 5704
rect 6454 5692 6460 5704
rect 5960 5664 6460 5692
rect 5960 5652 5966 5664
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 1949 5627 2007 5633
rect 1949 5593 1961 5627
rect 1995 5624 2007 5627
rect 2409 5627 2467 5633
rect 2409 5624 2421 5627
rect 1995 5596 2421 5624
rect 1995 5593 2007 5596
rect 1949 5587 2007 5593
rect 2409 5593 2421 5596
rect 2455 5624 2467 5627
rect 3786 5624 3792 5636
rect 2455 5596 3792 5624
rect 2455 5593 2467 5596
rect 2409 5587 2467 5593
rect 3786 5584 3792 5596
rect 3844 5584 3850 5636
rect 4706 5624 4712 5636
rect 4667 5596 4712 5624
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 6638 5584 6644 5636
rect 6696 5624 6702 5636
rect 7193 5627 7251 5633
rect 7193 5624 7205 5627
rect 6696 5596 7205 5624
rect 6696 5584 6702 5596
rect 7193 5593 7205 5596
rect 7239 5593 7251 5627
rect 7193 5587 7251 5593
rect 2130 5516 2136 5568
rect 2188 5556 2194 5568
rect 2958 5556 2964 5568
rect 2188 5528 2964 5556
rect 2188 5516 2194 5528
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 4154 5556 4160 5568
rect 4115 5528 4160 5556
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 1012 5466 8071 5488
rect 1012 5414 2582 5466
rect 2634 5414 2646 5466
rect 2698 5414 2710 5466
rect 2762 5414 2774 5466
rect 2826 5414 2838 5466
rect 2890 5414 4307 5466
rect 4359 5414 4371 5466
rect 4423 5414 4435 5466
rect 4487 5414 4499 5466
rect 4551 5414 4563 5466
rect 4615 5414 6032 5466
rect 6084 5414 6096 5466
rect 6148 5414 6160 5466
rect 6212 5414 6224 5466
rect 6276 5414 6288 5466
rect 6340 5414 7757 5466
rect 7809 5414 7821 5466
rect 7873 5414 7885 5466
rect 7937 5414 7949 5466
rect 8001 5414 8013 5466
rect 8065 5414 8071 5466
rect 1012 5392 8071 5414
rect 8294 5352 8300 5364
rect 4080 5324 8300 5352
rect 2685 5287 2743 5293
rect 2685 5253 2697 5287
rect 2731 5284 2743 5287
rect 3142 5284 3148 5296
rect 2731 5256 3148 5284
rect 2731 5253 2743 5256
rect 2685 5247 2743 5253
rect 3142 5244 3148 5256
rect 3200 5244 3206 5296
rect 4080 5293 4108 5324
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 4065 5287 4123 5293
rect 4065 5253 4077 5287
rect 4111 5253 4123 5287
rect 4065 5247 4123 5253
rect 5445 5287 5503 5293
rect 5445 5253 5457 5287
rect 5491 5284 5503 5287
rect 5626 5284 5632 5296
rect 5491 5256 5632 5284
rect 5491 5253 5503 5256
rect 5445 5247 5503 5253
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 7374 5284 7380 5296
rect 7335 5256 7380 5284
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 2038 5216 2044 5228
rect 1995 5188 2044 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 2746 5188 3341 5216
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 2746 5148 2774 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4212 5188 4721 5216
rect 4212 5176 4218 5188
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 1360 5120 2774 5148
rect 1360 5108 1366 5120
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 6549 5151 6607 5157
rect 6549 5148 6561 5151
rect 6420 5120 6561 5148
rect 6420 5108 6426 5120
rect 6549 5117 6561 5120
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 1012 4922 7912 4944
rect 1012 4870 1720 4922
rect 1772 4870 1784 4922
rect 1836 4870 1848 4922
rect 1900 4870 1912 4922
rect 1964 4870 1976 4922
rect 2028 4870 3445 4922
rect 3497 4870 3509 4922
rect 3561 4870 3573 4922
rect 3625 4870 3637 4922
rect 3689 4870 3701 4922
rect 3753 4870 5170 4922
rect 5222 4870 5234 4922
rect 5286 4870 5298 4922
rect 5350 4870 5362 4922
rect 5414 4870 5426 4922
rect 5478 4870 6895 4922
rect 6947 4870 6959 4922
rect 7011 4870 7023 4922
rect 7075 4870 7087 4922
rect 7139 4870 7151 4922
rect 7203 4870 7912 4922
rect 1012 4848 7912 4870
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3878 4808 3884 4820
rect 3752 4780 3884 4808
rect 3752 4768 3758 4780
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 8202 4808 8208 4820
rect 5500 4780 8208 4808
rect 5500 4768 5506 4780
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 2498 4672 2504 4684
rect 2459 4644 2504 4672
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 7558 4672 7564 4684
rect 5767 4644 7564 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 7558 4632 7564 4644
rect 7616 4632 7622 4684
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7466 4604 7472 4616
rect 7423 4576 7472 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 3142 4496 3148 4548
rect 3200 4536 3206 4548
rect 3329 4539 3387 4545
rect 3329 4536 3341 4539
rect 3200 4508 3341 4536
rect 3200 4496 3206 4508
rect 3329 4505 3341 4508
rect 3375 4505 3387 4539
rect 3329 4499 3387 4505
rect 4893 4539 4951 4545
rect 4893 4505 4905 4539
rect 4939 4536 4951 4539
rect 5718 4536 5724 4548
rect 4939 4508 5724 4536
rect 4939 4505 4951 4508
rect 4893 4499 4951 4505
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 6454 4496 6460 4548
rect 6512 4536 6518 4548
rect 6549 4539 6607 4545
rect 6549 4536 6561 4539
rect 6512 4508 6561 4536
rect 6512 4496 6518 4508
rect 6549 4505 6561 4508
rect 6595 4505 6607 4539
rect 6549 4499 6607 4505
rect 750 4428 756 4480
rect 808 4468 814 4480
rect 1302 4468 1308 4480
rect 808 4440 1308 4468
rect 808 4428 814 4440
rect 1302 4428 1308 4440
rect 1360 4468 1366 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1360 4440 1869 4468
rect 1360 4428 1366 4440
rect 1857 4437 1869 4440
rect 1903 4437 1915 4471
rect 1857 4431 1915 4437
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 4341 4471 4399 4477
rect 4341 4468 4353 4471
rect 3292 4440 4353 4468
rect 3292 4428 3298 4440
rect 4341 4437 4353 4440
rect 4387 4468 4399 4471
rect 4706 4468 4712 4480
rect 4387 4440 4712 4468
rect 4387 4437 4399 4440
rect 4341 4431 4399 4437
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 1012 4378 8071 4400
rect 1012 4326 2582 4378
rect 2634 4326 2646 4378
rect 2698 4326 2710 4378
rect 2762 4326 2774 4378
rect 2826 4326 2838 4378
rect 2890 4326 4307 4378
rect 4359 4326 4371 4378
rect 4423 4326 4435 4378
rect 4487 4326 4499 4378
rect 4551 4326 4563 4378
rect 4615 4326 6032 4378
rect 6084 4326 6096 4378
rect 6148 4326 6160 4378
rect 6212 4326 6224 4378
rect 6276 4326 6288 4378
rect 6340 4326 7757 4378
rect 7809 4326 7821 4378
rect 7873 4326 7885 4378
rect 7937 4326 7949 4378
rect 8001 4326 8013 4378
rect 8065 4326 8071 4378
rect 1012 4304 8071 4326
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 5534 4264 5540 4276
rect 3660 4236 5540 4264
rect 3660 4224 3666 4236
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 3697 4199 3755 4205
rect 3697 4165 3709 4199
rect 3743 4196 3755 4199
rect 4798 4196 4804 4208
rect 3743 4168 4804 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 7377 4199 7435 4205
rect 7377 4165 7389 4199
rect 7423 4196 7435 4199
rect 7650 4196 7656 4208
rect 7423 4168 7656 4196
rect 7423 4165 7435 4168
rect 7377 4159 7435 4165
rect 7650 4156 7656 4168
rect 7708 4156 7714 4208
rect 2958 4128 2964 4140
rect 2919 4100 2964 4128
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 3528 4100 4261 4128
rect 3528 4060 3556 4100
rect 4249 4097 4261 4100
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5442 4128 5448 4140
rect 5123 4100 5448 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5902 4128 5908 4140
rect 5863 4100 5908 4128
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 2240 4032 3556 4060
rect 290 3952 296 4004
rect 348 3992 354 4004
rect 2240 4001 2268 4032
rect 3694 4020 3700 4072
rect 3752 4060 3758 4072
rect 5626 4060 5632 4072
rect 3752 4032 5632 4060
rect 3752 4020 3758 4032
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 6546 4060 6552 4072
rect 6507 4032 6552 4060
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 2225 3995 2283 4001
rect 2225 3992 2237 3995
rect 348 3964 2237 3992
rect 348 3952 354 3964
rect 2225 3961 2237 3964
rect 2271 3961 2283 3995
rect 2225 3955 2283 3961
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 2038 3924 2044 3936
rect 1811 3896 2044 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 2038 3884 2044 3896
rect 2096 3924 2102 3936
rect 4154 3924 4160 3936
rect 2096 3896 4160 3924
rect 2096 3884 2102 3896
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 1012 3834 7912 3856
rect 1012 3782 1720 3834
rect 1772 3782 1784 3834
rect 1836 3782 1848 3834
rect 1900 3782 1912 3834
rect 1964 3782 1976 3834
rect 2028 3782 3445 3834
rect 3497 3782 3509 3834
rect 3561 3782 3573 3834
rect 3625 3782 3637 3834
rect 3689 3782 3701 3834
rect 3753 3782 5170 3834
rect 5222 3782 5234 3834
rect 5286 3782 5298 3834
rect 5350 3782 5362 3834
rect 5414 3782 5426 3834
rect 5478 3782 6895 3834
rect 6947 3782 6959 3834
rect 7011 3782 7023 3834
rect 7075 3782 7087 3834
rect 7139 3782 7151 3834
rect 7203 3782 7912 3834
rect 1012 3760 7912 3782
rect 2038 3680 2044 3732
rect 2096 3720 2102 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 2096 3692 3893 3720
rect 2096 3680 2102 3692
rect 3881 3689 3893 3692
rect 3927 3720 3939 3723
rect 4246 3720 4252 3732
rect 3927 3692 4252 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 7374 3720 7380 3732
rect 7335 3692 7380 3720
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 6825 3655 6883 3661
rect 6825 3621 6837 3655
rect 6871 3652 6883 3655
rect 7466 3652 7472 3664
rect 6871 3624 7472 3652
rect 6871 3621 6883 3624
rect 6825 3615 6883 3621
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3584 2651 3587
rect 3050 3584 3056 3596
rect 2639 3556 3056 3584
rect 2639 3553 2651 3556
rect 2593 3547 2651 3553
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 5261 3587 5319 3593
rect 5261 3553 5273 3587
rect 5307 3584 5319 3587
rect 5810 3584 5816 3596
rect 5307 3556 5816 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 2130 3476 2136 3528
rect 2188 3516 2194 3528
rect 2188 3488 4476 3516
rect 2188 3476 2194 3488
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 3329 3451 3387 3457
rect 3329 3448 3341 3451
rect 1728 3420 3341 3448
rect 1728 3408 1734 3420
rect 3329 3417 3341 3420
rect 3375 3417 3387 3451
rect 3329 3411 3387 3417
rect 1949 3383 2007 3389
rect 1949 3349 1961 3383
rect 1995 3380 2007 3383
rect 3142 3380 3148 3392
rect 1995 3352 3148 3380
rect 1995 3349 2007 3352
rect 1949 3343 2007 3349
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 3344 3380 3372 3411
rect 3878 3408 3884 3460
rect 3936 3448 3942 3460
rect 4062 3448 4068 3460
rect 3936 3420 4068 3448
rect 3936 3408 3942 3420
rect 4062 3408 4068 3420
rect 4120 3408 4126 3460
rect 4448 3457 4476 3488
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 4706 3448 4712 3460
rect 4479 3420 4712 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 5905 3451 5963 3457
rect 5905 3448 5917 3451
rect 5776 3420 5917 3448
rect 5776 3408 5782 3420
rect 5905 3417 5917 3420
rect 5951 3417 5963 3451
rect 5905 3411 5963 3417
rect 5810 3380 5816 3392
rect 3344 3352 5816 3380
rect 5810 3340 5816 3352
rect 5868 3340 5874 3392
rect 1012 3290 8071 3312
rect 1012 3238 2582 3290
rect 2634 3238 2646 3290
rect 2698 3238 2710 3290
rect 2762 3238 2774 3290
rect 2826 3238 2838 3290
rect 2890 3238 4307 3290
rect 4359 3238 4371 3290
rect 4423 3238 4435 3290
rect 4487 3238 4499 3290
rect 4551 3238 4563 3290
rect 4615 3238 6032 3290
rect 6084 3238 6096 3290
rect 6148 3238 6160 3290
rect 6212 3238 6224 3290
rect 6276 3238 6288 3290
rect 6340 3238 7757 3290
rect 7809 3238 7821 3290
rect 7873 3238 7885 3290
rect 7937 3238 7949 3290
rect 8001 3238 8013 3290
rect 8065 3238 8071 3290
rect 1012 3216 8071 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3200 3148 4292 3176
rect 3200 3136 3206 3148
rect 4157 3111 4215 3117
rect 4157 3108 4169 3111
rect 2746 3080 4169 3108
rect 2746 2972 2774 3080
rect 4157 3077 4169 3080
rect 4203 3077 4215 3111
rect 4157 3071 4215 3077
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3326 3040 3332 3052
rect 2915 3012 3332 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 2424 2944 2774 2972
rect 2424 2848 2452 2944
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2406 2836 2412 2848
rect 2271 2808 2412 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 2406 2796 2412 2808
rect 2464 2796 2470 2848
rect 3142 2796 3148 2848
rect 3200 2836 3206 2848
rect 3620 2836 3648 3003
rect 4264 2972 4292 3148
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 6457 3179 6515 3185
rect 6457 3176 6469 3179
rect 4764 3148 6469 3176
rect 4764 3136 4770 3148
rect 6457 3145 6469 3148
rect 6503 3145 6515 3179
rect 6457 3139 6515 3145
rect 7377 3179 7435 3185
rect 7377 3145 7389 3179
rect 7423 3176 7435 3179
rect 7650 3176 7656 3188
rect 7423 3148 7656 3176
rect 7423 3145 7435 3148
rect 7377 3139 7435 3145
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 4985 3111 5043 3117
rect 4985 3077 4997 3111
rect 5031 3108 5043 3111
rect 5074 3108 5080 3120
rect 5031 3080 5080 3108
rect 5031 3077 5043 3080
rect 4985 3071 5043 3077
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 5626 3068 5632 3120
rect 5684 3108 5690 3120
rect 6270 3108 6276 3120
rect 5684 3080 6276 3108
rect 5684 3068 5690 3080
rect 6270 3068 6276 3080
rect 6328 3068 6334 3120
rect 4798 3000 4804 3052
rect 4856 3040 4862 3052
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 4856 3012 5549 3040
rect 4856 3000 4862 3012
rect 5092 2984 5120 3012
rect 5537 3009 5549 3012
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 4982 2972 4988 2984
rect 4264 2944 4988 2972
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5074 2932 5080 2984
rect 5132 2932 5138 2984
rect 6638 2836 6644 2848
rect 3200 2808 6644 2836
rect 3200 2796 3206 2808
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 1012 2746 7912 2768
rect 1012 2694 1720 2746
rect 1772 2694 1784 2746
rect 1836 2694 1848 2746
rect 1900 2694 1912 2746
rect 1964 2694 1976 2746
rect 2028 2694 3445 2746
rect 3497 2694 3509 2746
rect 3561 2694 3573 2746
rect 3625 2694 3637 2746
rect 3689 2694 3701 2746
rect 3753 2694 5170 2746
rect 5222 2694 5234 2746
rect 5286 2694 5298 2746
rect 5350 2694 5362 2746
rect 5414 2694 5426 2746
rect 5478 2694 6895 2746
rect 6947 2694 6959 2746
rect 7011 2694 7023 2746
rect 7075 2694 7087 2746
rect 7139 2694 7151 2746
rect 7203 2694 7912 2746
rect 1012 2672 7912 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 3142 2632 3148 2644
rect 1995 2604 3148 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 3786 2524 3792 2576
rect 3844 2564 3850 2576
rect 7193 2567 7251 2573
rect 7193 2564 7205 2567
rect 3844 2536 7205 2564
rect 3844 2524 3850 2536
rect 7193 2533 7205 2536
rect 7239 2533 7251 2567
rect 7193 2527 7251 2533
rect 1210 2456 1216 2508
rect 1268 2496 1274 2508
rect 2501 2499 2559 2505
rect 2501 2496 2513 2499
rect 1268 2468 2513 2496
rect 1268 2456 1274 2468
rect 2501 2465 2513 2468
rect 2547 2465 2559 2499
rect 2501 2459 2559 2465
rect 4709 2499 4767 2505
rect 4709 2465 4721 2499
rect 4755 2496 4767 2499
rect 4890 2496 4896 2508
rect 4755 2468 4896 2496
rect 4755 2465 4767 2468
rect 4709 2459 4767 2465
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 5445 2499 5503 2505
rect 5445 2465 5457 2499
rect 5491 2496 5503 2499
rect 5534 2496 5540 2508
rect 5491 2468 5540 2496
rect 5491 2465 5503 2468
rect 5445 2459 5503 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 7282 2428 7288 2440
rect 3344 2400 7288 2428
rect 1578 2320 1584 2372
rect 1636 2360 1642 2372
rect 3344 2369 3372 2400
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 3329 2363 3387 2369
rect 3329 2360 3341 2363
rect 1636 2332 3341 2360
rect 1636 2320 1642 2332
rect 3329 2329 3341 2332
rect 3375 2329 3387 2363
rect 3329 2323 3387 2329
rect 3881 2363 3939 2369
rect 3881 2329 3893 2363
rect 3927 2329 3939 2363
rect 3881 2323 3939 2329
rect 6181 2363 6239 2369
rect 6181 2329 6193 2363
rect 6227 2360 6239 2363
rect 6227 2332 6776 2360
rect 6227 2329 6239 2332
rect 6181 2323 6239 2329
rect 3050 2252 3056 2304
rect 3108 2292 3114 2304
rect 3786 2292 3792 2304
rect 3108 2264 3792 2292
rect 3108 2252 3114 2264
rect 3786 2252 3792 2264
rect 3844 2292 3850 2304
rect 3896 2292 3924 2323
rect 6748 2304 6776 2332
rect 6730 2292 6736 2304
rect 3844 2264 3924 2292
rect 6691 2264 6736 2292
rect 3844 2252 3850 2264
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 1012 2202 8071 2224
rect 1012 2150 2582 2202
rect 2634 2150 2646 2202
rect 2698 2150 2710 2202
rect 2762 2150 2774 2202
rect 2826 2150 2838 2202
rect 2890 2150 4307 2202
rect 4359 2150 4371 2202
rect 4423 2150 4435 2202
rect 4487 2150 4499 2202
rect 4551 2150 4563 2202
rect 4615 2150 6032 2202
rect 6084 2150 6096 2202
rect 6148 2150 6160 2202
rect 6212 2150 6224 2202
rect 6276 2150 6288 2202
rect 6340 2150 7757 2202
rect 7809 2150 7821 2202
rect 7873 2150 7885 2202
rect 7937 2150 7949 2202
rect 8001 2150 8013 2202
rect 8065 2150 8071 2202
rect 1012 2128 8071 2150
rect 1578 2088 1584 2100
rect 1539 2060 1584 2088
rect 1578 2048 1584 2060
rect 1636 2048 1642 2100
rect 2133 2091 2191 2097
rect 2133 2057 2145 2091
rect 2179 2088 2191 2091
rect 2314 2088 2320 2100
rect 2179 2060 2320 2088
rect 2179 2057 2191 2060
rect 2133 2051 2191 2057
rect 2314 2048 2320 2060
rect 2372 2048 2378 2100
rect 2777 2023 2835 2029
rect 2777 1989 2789 2023
rect 2823 2020 2835 2023
rect 2958 2020 2964 2032
rect 2823 1992 2964 2020
rect 2823 1989 2835 1992
rect 2777 1983 2835 1989
rect 2958 1980 2964 1992
rect 3016 1980 3022 2032
rect 3326 1980 3332 2032
rect 3384 2020 3390 2032
rect 6549 2023 6607 2029
rect 6549 2020 6561 2023
rect 3384 1992 6561 2020
rect 3384 1980 3390 1992
rect 6549 1989 6561 1992
rect 6595 1989 6607 2023
rect 6549 1983 6607 1989
rect 3513 1955 3571 1961
rect 3513 1921 3525 1955
rect 3559 1952 3571 1955
rect 3786 1952 3792 1964
rect 3559 1924 3792 1952
rect 3559 1921 3571 1924
rect 3513 1915 3571 1921
rect 3786 1912 3792 1924
rect 3844 1912 3850 1964
rect 4062 1952 4068 1964
rect 4023 1924 4068 1952
rect 4062 1912 4068 1924
rect 4120 1912 4126 1964
rect 4893 1955 4951 1961
rect 4893 1921 4905 1955
rect 4939 1952 4951 1955
rect 7374 1952 7380 1964
rect 4939 1924 5488 1952
rect 7335 1924 7380 1952
rect 4939 1921 4951 1924
rect 4893 1915 4951 1921
rect 5460 1757 5488 1924
rect 7374 1912 7380 1924
rect 7432 1912 7438 1964
rect 5445 1751 5503 1757
rect 5445 1717 5457 1751
rect 5491 1748 5503 1751
rect 8110 1748 8116 1760
rect 5491 1720 8116 1748
rect 5491 1717 5503 1720
rect 5445 1711 5503 1717
rect 8110 1708 8116 1720
rect 8168 1708 8174 1760
rect 1012 1658 7912 1680
rect 1012 1606 1720 1658
rect 1772 1606 1784 1658
rect 1836 1606 1848 1658
rect 1900 1606 1912 1658
rect 1964 1606 1976 1658
rect 2028 1606 3445 1658
rect 3497 1606 3509 1658
rect 3561 1606 3573 1658
rect 3625 1606 3637 1658
rect 3689 1606 3701 1658
rect 3753 1606 5170 1658
rect 5222 1606 5234 1658
rect 5286 1606 5298 1658
rect 5350 1606 5362 1658
rect 5414 1606 5426 1658
rect 5478 1606 6895 1658
rect 6947 1606 6959 1658
rect 7011 1606 7023 1658
rect 7075 1606 7087 1658
rect 7139 1606 7151 1658
rect 7203 1606 7912 1658
rect 1012 1584 7912 1606
rect 3786 1504 3792 1556
rect 3844 1544 3850 1556
rect 8570 1544 8576 1556
rect 3844 1516 8576 1544
rect 3844 1504 3850 1516
rect 8570 1504 8576 1516
rect 8628 1504 8634 1556
rect 3804 1408 3832 1504
rect 3252 1380 3832 1408
rect 4065 1411 4123 1417
rect 1949 1343 2007 1349
rect 1949 1309 1961 1343
rect 1995 1340 2007 1343
rect 3252 1340 3280 1380
rect 4065 1377 4077 1411
rect 4111 1408 4123 1411
rect 4706 1408 4712 1420
rect 4111 1380 4712 1408
rect 4111 1377 4123 1380
rect 4065 1371 4123 1377
rect 4706 1368 4712 1380
rect 4764 1368 4770 1420
rect 1995 1312 3280 1340
rect 3329 1343 3387 1349
rect 1995 1309 2007 1312
rect 1949 1303 2007 1309
rect 3329 1309 3341 1343
rect 3375 1340 3387 1343
rect 5902 1340 5908 1352
rect 3375 1312 5908 1340
rect 3375 1309 3387 1312
rect 3329 1303 3387 1309
rect 5902 1300 5908 1312
rect 5960 1300 5966 1352
rect 2498 1272 2504 1284
rect 2459 1244 2504 1272
rect 2498 1232 2504 1244
rect 2556 1232 2562 1284
rect 4801 1275 4859 1281
rect 4801 1241 4813 1275
rect 4847 1272 4859 1275
rect 5353 1275 5411 1281
rect 5353 1272 5365 1275
rect 4847 1244 5365 1272
rect 4847 1241 4859 1244
rect 4801 1235 4859 1241
rect 5353 1241 5365 1244
rect 5399 1272 5411 1275
rect 7650 1272 7656 1284
rect 5399 1244 7656 1272
rect 5399 1241 5411 1244
rect 5353 1235 5411 1241
rect 7650 1232 7656 1244
rect 7708 1232 7714 1284
rect 1210 1164 1216 1216
rect 1268 1204 1274 1216
rect 5718 1204 5724 1216
rect 1268 1176 5724 1204
rect 1268 1164 1274 1176
rect 5718 1164 5724 1176
rect 5776 1164 5782 1216
rect 7374 1204 7380 1216
rect 7335 1176 7380 1204
rect 7374 1164 7380 1176
rect 7432 1164 7438 1216
rect 1012 1114 8071 1136
rect 1012 1062 2582 1114
rect 2634 1062 2646 1114
rect 2698 1062 2710 1114
rect 2762 1062 2774 1114
rect 2826 1062 2838 1114
rect 2890 1062 4307 1114
rect 4359 1062 4371 1114
rect 4423 1062 4435 1114
rect 4487 1062 4499 1114
rect 4551 1062 4563 1114
rect 4615 1062 6032 1114
rect 6084 1062 6096 1114
rect 6148 1062 6160 1114
rect 6212 1062 6224 1114
rect 6276 1062 6288 1114
rect 6340 1062 7757 1114
rect 7809 1062 7821 1114
rect 7873 1062 7885 1114
rect 7937 1062 7949 1114
rect 8001 1062 8013 1114
rect 8065 1062 8071 1114
rect 1012 1040 8071 1062
rect 2406 960 2412 1012
rect 2464 1000 2470 1012
rect 2590 1000 2596 1012
rect 2464 972 2596 1000
rect 2464 960 2470 972
rect 2590 960 2596 972
rect 2648 960 2654 1012
<< via1 >>
rect 5632 9392 5684 9444
rect 6368 9392 6420 9444
rect 7840 9392 7892 9444
rect 8300 9392 8352 9444
rect 4068 8848 4120 8900
rect 5540 8848 5592 8900
rect 5172 8780 5224 8832
rect 6644 8780 6696 8832
rect 2582 8678 2634 8730
rect 2646 8678 2698 8730
rect 2710 8678 2762 8730
rect 2774 8678 2826 8730
rect 2838 8678 2890 8730
rect 4307 8678 4359 8730
rect 4371 8678 4423 8730
rect 4435 8678 4487 8730
rect 4499 8678 4551 8730
rect 4563 8678 4615 8730
rect 6032 8678 6084 8730
rect 6096 8678 6148 8730
rect 6160 8678 6212 8730
rect 6224 8678 6276 8730
rect 6288 8678 6340 8730
rect 7757 8678 7809 8730
rect 7821 8678 7873 8730
rect 7885 8678 7937 8730
rect 7949 8678 8001 8730
rect 8013 8678 8065 8730
rect 1860 8619 1912 8628
rect 1860 8585 1869 8619
rect 1869 8585 1903 8619
rect 1903 8585 1912 8619
rect 1860 8576 1912 8585
rect 3700 8576 3752 8628
rect 4712 8576 4764 8628
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 3884 8440 3936 8492
rect 4252 8372 4304 8424
rect 5908 8372 5960 8424
rect 8116 8372 8168 8424
rect 940 8304 992 8356
rect 1492 8304 1544 8356
rect 2320 8304 2372 8356
rect 4068 8304 4120 8356
rect 1720 8134 1772 8186
rect 1784 8134 1836 8186
rect 1848 8134 1900 8186
rect 1912 8134 1964 8186
rect 1976 8134 2028 8186
rect 3445 8134 3497 8186
rect 3509 8134 3561 8186
rect 3573 8134 3625 8186
rect 3637 8134 3689 8186
rect 3701 8134 3753 8186
rect 5170 8134 5222 8186
rect 5234 8134 5286 8186
rect 5298 8134 5350 8186
rect 5362 8134 5414 8186
rect 5426 8134 5478 8186
rect 6895 8134 6947 8186
rect 6959 8134 7011 8186
rect 7023 8134 7075 8186
rect 7087 8134 7139 8186
rect 7151 8134 7203 8186
rect 2964 8032 3016 8084
rect 3884 8032 3936 8084
rect 6644 8032 6696 8084
rect 4804 7964 4856 8016
rect 5172 7964 5224 8016
rect 1492 7828 1544 7880
rect 1308 7760 1360 7812
rect 4068 7828 4120 7880
rect 4160 7760 4212 7812
rect 4804 7803 4856 7812
rect 4804 7769 4813 7803
rect 4813 7769 4847 7803
rect 4847 7769 4856 7803
rect 4804 7760 4856 7769
rect 6368 7760 6420 7812
rect 7196 7692 7248 7744
rect 2582 7590 2634 7642
rect 2646 7590 2698 7642
rect 2710 7590 2762 7642
rect 2774 7590 2826 7642
rect 2838 7590 2890 7642
rect 4307 7590 4359 7642
rect 4371 7590 4423 7642
rect 4435 7590 4487 7642
rect 4499 7590 4551 7642
rect 4563 7590 4615 7642
rect 6032 7590 6084 7642
rect 6096 7590 6148 7642
rect 6160 7590 6212 7642
rect 6224 7590 6276 7642
rect 6288 7590 6340 7642
rect 7757 7590 7809 7642
rect 7821 7590 7873 7642
rect 7885 7590 7937 7642
rect 7949 7590 8001 7642
rect 8013 7590 8065 7642
rect 1308 7488 1360 7540
rect 5356 7488 5408 7540
rect 4712 7420 4764 7472
rect 5540 7420 5592 7472
rect 7196 7420 7248 7472
rect 7288 7420 7340 7472
rect 7564 7420 7616 7472
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 3240 7352 3292 7404
rect 6552 7352 6604 7404
rect 5540 7284 5592 7336
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 4988 7148 5040 7200
rect 5172 7148 5224 7200
rect 1720 7046 1772 7098
rect 1784 7046 1836 7098
rect 1848 7046 1900 7098
rect 1912 7046 1964 7098
rect 1976 7046 2028 7098
rect 3445 7046 3497 7098
rect 3509 7046 3561 7098
rect 3573 7046 3625 7098
rect 3637 7046 3689 7098
rect 3701 7046 3753 7098
rect 5170 7046 5222 7098
rect 5234 7046 5286 7098
rect 5298 7046 5350 7098
rect 5362 7046 5414 7098
rect 5426 7046 5478 7098
rect 6895 7046 6947 7098
rect 6959 7046 7011 7098
rect 7023 7046 7075 7098
rect 7087 7046 7139 7098
rect 7151 7046 7203 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 1584 6944 1636 6996
rect 2228 6944 2280 6996
rect 5724 6740 5776 6792
rect 3056 6604 3108 6656
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 4988 6672 5040 6724
rect 6552 6672 6604 6724
rect 4804 6604 4856 6656
rect 5264 6604 5316 6656
rect 7472 6604 7524 6656
rect 2582 6502 2634 6554
rect 2646 6502 2698 6554
rect 2710 6502 2762 6554
rect 2774 6502 2826 6554
rect 2838 6502 2890 6554
rect 4307 6502 4359 6554
rect 4371 6502 4423 6554
rect 4435 6502 4487 6554
rect 4499 6502 4551 6554
rect 4563 6502 4615 6554
rect 6032 6502 6084 6554
rect 6096 6502 6148 6554
rect 6160 6502 6212 6554
rect 6224 6502 6276 6554
rect 6288 6502 6340 6554
rect 7757 6502 7809 6554
rect 7821 6502 7873 6554
rect 7885 6502 7937 6554
rect 7949 6502 8001 6554
rect 8013 6502 8065 6554
rect 5724 6400 5776 6452
rect 1032 6332 1084 6384
rect 3792 6332 3844 6384
rect 5264 6375 5316 6384
rect 5264 6341 5273 6375
rect 5273 6341 5307 6375
rect 5307 6341 5316 6375
rect 5264 6332 5316 6341
rect 6644 6332 6696 6384
rect 6736 6332 6788 6384
rect 7380 6332 7432 6384
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 4252 6264 4304 6316
rect 3056 6196 3108 6248
rect 3884 6196 3936 6248
rect 6736 6196 6788 6248
rect 1720 5958 1772 6010
rect 1784 5958 1836 6010
rect 1848 5958 1900 6010
rect 1912 5958 1964 6010
rect 1976 5958 2028 6010
rect 3445 5958 3497 6010
rect 3509 5958 3561 6010
rect 3573 5958 3625 6010
rect 3637 5958 3689 6010
rect 3701 5958 3753 6010
rect 5170 5958 5222 6010
rect 5234 5958 5286 6010
rect 5298 5958 5350 6010
rect 5362 5958 5414 6010
rect 5426 5958 5478 6010
rect 6895 5958 6947 6010
rect 6959 5958 7011 6010
rect 7023 5958 7075 6010
rect 7087 5958 7139 6010
rect 7151 5958 7203 6010
rect 4068 5720 4120 5772
rect 5448 5763 5500 5772
rect 5448 5729 5457 5763
rect 5457 5729 5491 5763
rect 5491 5729 5500 5763
rect 5448 5720 5500 5729
rect 1400 5652 1452 5704
rect 3056 5652 3108 5704
rect 5908 5652 5960 5704
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 3792 5584 3844 5636
rect 4712 5627 4764 5636
rect 4712 5593 4721 5627
rect 4721 5593 4755 5627
rect 4755 5593 4764 5627
rect 4712 5584 4764 5593
rect 6644 5584 6696 5636
rect 2136 5516 2188 5568
rect 2964 5516 3016 5568
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 2582 5414 2634 5466
rect 2646 5414 2698 5466
rect 2710 5414 2762 5466
rect 2774 5414 2826 5466
rect 2838 5414 2890 5466
rect 4307 5414 4359 5466
rect 4371 5414 4423 5466
rect 4435 5414 4487 5466
rect 4499 5414 4551 5466
rect 4563 5414 4615 5466
rect 6032 5414 6084 5466
rect 6096 5414 6148 5466
rect 6160 5414 6212 5466
rect 6224 5414 6276 5466
rect 6288 5414 6340 5466
rect 7757 5414 7809 5466
rect 7821 5414 7873 5466
rect 7885 5414 7937 5466
rect 7949 5414 8001 5466
rect 8013 5414 8065 5466
rect 3148 5244 3200 5296
rect 8300 5312 8352 5364
rect 5632 5244 5684 5296
rect 7380 5287 7432 5296
rect 7380 5253 7389 5287
rect 7389 5253 7423 5287
rect 7423 5253 7432 5287
rect 7380 5244 7432 5253
rect 2044 5176 2096 5228
rect 1308 5108 1360 5160
rect 4160 5176 4212 5228
rect 6368 5108 6420 5160
rect 1720 4870 1772 4922
rect 1784 4870 1836 4922
rect 1848 4870 1900 4922
rect 1912 4870 1964 4922
rect 1976 4870 2028 4922
rect 3445 4870 3497 4922
rect 3509 4870 3561 4922
rect 3573 4870 3625 4922
rect 3637 4870 3689 4922
rect 3701 4870 3753 4922
rect 5170 4870 5222 4922
rect 5234 4870 5286 4922
rect 5298 4870 5350 4922
rect 5362 4870 5414 4922
rect 5426 4870 5478 4922
rect 6895 4870 6947 4922
rect 6959 4870 7011 4922
rect 7023 4870 7075 4922
rect 7087 4870 7139 4922
rect 7151 4870 7203 4922
rect 3700 4768 3752 4820
rect 3884 4768 3936 4820
rect 5448 4768 5500 4820
rect 8208 4768 8260 4820
rect 2504 4675 2556 4684
rect 2504 4641 2513 4675
rect 2513 4641 2547 4675
rect 2547 4641 2556 4675
rect 2504 4632 2556 4641
rect 7564 4632 7616 4684
rect 7472 4564 7524 4616
rect 3148 4496 3200 4548
rect 5724 4496 5776 4548
rect 6460 4496 6512 4548
rect 756 4428 808 4480
rect 1308 4428 1360 4480
rect 3240 4428 3292 4480
rect 4712 4428 4764 4480
rect 2582 4326 2634 4378
rect 2646 4326 2698 4378
rect 2710 4326 2762 4378
rect 2774 4326 2826 4378
rect 2838 4326 2890 4378
rect 4307 4326 4359 4378
rect 4371 4326 4423 4378
rect 4435 4326 4487 4378
rect 4499 4326 4551 4378
rect 4563 4326 4615 4378
rect 6032 4326 6084 4378
rect 6096 4326 6148 4378
rect 6160 4326 6212 4378
rect 6224 4326 6276 4378
rect 6288 4326 6340 4378
rect 7757 4326 7809 4378
rect 7821 4326 7873 4378
rect 7885 4326 7937 4378
rect 7949 4326 8001 4378
rect 8013 4326 8065 4378
rect 3608 4224 3660 4276
rect 5540 4224 5592 4276
rect 4804 4156 4856 4208
rect 7656 4156 7708 4208
rect 2964 4131 3016 4140
rect 2964 4097 2973 4131
rect 2973 4097 3007 4131
rect 3007 4097 3016 4131
rect 2964 4088 3016 4097
rect 5448 4088 5500 4140
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 296 3952 348 4004
rect 3700 4020 3752 4072
rect 5632 4020 5684 4072
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 2044 3884 2096 3936
rect 4160 3884 4212 3936
rect 1720 3782 1772 3834
rect 1784 3782 1836 3834
rect 1848 3782 1900 3834
rect 1912 3782 1964 3834
rect 1976 3782 2028 3834
rect 3445 3782 3497 3834
rect 3509 3782 3561 3834
rect 3573 3782 3625 3834
rect 3637 3782 3689 3834
rect 3701 3782 3753 3834
rect 5170 3782 5222 3834
rect 5234 3782 5286 3834
rect 5298 3782 5350 3834
rect 5362 3782 5414 3834
rect 5426 3782 5478 3834
rect 6895 3782 6947 3834
rect 6959 3782 7011 3834
rect 7023 3782 7075 3834
rect 7087 3782 7139 3834
rect 7151 3782 7203 3834
rect 2044 3680 2096 3732
rect 4252 3680 4304 3732
rect 7380 3723 7432 3732
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 7472 3612 7524 3664
rect 3056 3544 3108 3596
rect 5816 3544 5868 3596
rect 2136 3476 2188 3528
rect 1676 3408 1728 3460
rect 3148 3340 3200 3392
rect 3884 3408 3936 3460
rect 4068 3408 4120 3460
rect 4712 3408 4764 3460
rect 5724 3408 5776 3460
rect 5816 3340 5868 3392
rect 2582 3238 2634 3290
rect 2646 3238 2698 3290
rect 2710 3238 2762 3290
rect 2774 3238 2826 3290
rect 2838 3238 2890 3290
rect 4307 3238 4359 3290
rect 4371 3238 4423 3290
rect 4435 3238 4487 3290
rect 4499 3238 4551 3290
rect 4563 3238 4615 3290
rect 6032 3238 6084 3290
rect 6096 3238 6148 3290
rect 6160 3238 6212 3290
rect 6224 3238 6276 3290
rect 6288 3238 6340 3290
rect 7757 3238 7809 3290
rect 7821 3238 7873 3290
rect 7885 3238 7937 3290
rect 7949 3238 8001 3290
rect 8013 3238 8065 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 3148 3136 3200 3188
rect 3332 3000 3384 3052
rect 2412 2796 2464 2848
rect 3148 2796 3200 2848
rect 4712 3136 4764 3188
rect 7656 3136 7708 3188
rect 5080 3068 5132 3120
rect 5632 3068 5684 3120
rect 6276 3068 6328 3120
rect 4804 3000 4856 3052
rect 4988 2932 5040 2984
rect 5080 2932 5132 2984
rect 6644 2796 6696 2848
rect 1720 2694 1772 2746
rect 1784 2694 1836 2746
rect 1848 2694 1900 2746
rect 1912 2694 1964 2746
rect 1976 2694 2028 2746
rect 3445 2694 3497 2746
rect 3509 2694 3561 2746
rect 3573 2694 3625 2746
rect 3637 2694 3689 2746
rect 3701 2694 3753 2746
rect 5170 2694 5222 2746
rect 5234 2694 5286 2746
rect 5298 2694 5350 2746
rect 5362 2694 5414 2746
rect 5426 2694 5478 2746
rect 6895 2694 6947 2746
rect 6959 2694 7011 2746
rect 7023 2694 7075 2746
rect 7087 2694 7139 2746
rect 7151 2694 7203 2746
rect 3148 2592 3200 2644
rect 3792 2524 3844 2576
rect 1216 2456 1268 2508
rect 4896 2456 4948 2508
rect 5540 2456 5592 2508
rect 1584 2320 1636 2372
rect 7288 2388 7340 2440
rect 3056 2252 3108 2304
rect 3792 2252 3844 2304
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 2582 2150 2634 2202
rect 2646 2150 2698 2202
rect 2710 2150 2762 2202
rect 2774 2150 2826 2202
rect 2838 2150 2890 2202
rect 4307 2150 4359 2202
rect 4371 2150 4423 2202
rect 4435 2150 4487 2202
rect 4499 2150 4551 2202
rect 4563 2150 4615 2202
rect 6032 2150 6084 2202
rect 6096 2150 6148 2202
rect 6160 2150 6212 2202
rect 6224 2150 6276 2202
rect 6288 2150 6340 2202
rect 7757 2150 7809 2202
rect 7821 2150 7873 2202
rect 7885 2150 7937 2202
rect 7949 2150 8001 2202
rect 8013 2150 8065 2202
rect 1584 2091 1636 2100
rect 1584 2057 1593 2091
rect 1593 2057 1627 2091
rect 1627 2057 1636 2091
rect 1584 2048 1636 2057
rect 2320 2048 2372 2100
rect 2964 1980 3016 2032
rect 3332 1980 3384 2032
rect 3792 1912 3844 1964
rect 4068 1955 4120 1964
rect 4068 1921 4077 1955
rect 4077 1921 4111 1955
rect 4111 1921 4120 1955
rect 4068 1912 4120 1921
rect 7380 1955 7432 1964
rect 7380 1921 7389 1955
rect 7389 1921 7423 1955
rect 7423 1921 7432 1955
rect 7380 1912 7432 1921
rect 8116 1708 8168 1760
rect 1720 1606 1772 1658
rect 1784 1606 1836 1658
rect 1848 1606 1900 1658
rect 1912 1606 1964 1658
rect 1976 1606 2028 1658
rect 3445 1606 3497 1658
rect 3509 1606 3561 1658
rect 3573 1606 3625 1658
rect 3637 1606 3689 1658
rect 3701 1606 3753 1658
rect 5170 1606 5222 1658
rect 5234 1606 5286 1658
rect 5298 1606 5350 1658
rect 5362 1606 5414 1658
rect 5426 1606 5478 1658
rect 6895 1606 6947 1658
rect 6959 1606 7011 1658
rect 7023 1606 7075 1658
rect 7087 1606 7139 1658
rect 7151 1606 7203 1658
rect 3792 1504 3844 1556
rect 8576 1504 8628 1556
rect 4712 1368 4764 1420
rect 5908 1343 5960 1352
rect 5908 1309 5917 1343
rect 5917 1309 5951 1343
rect 5951 1309 5960 1343
rect 5908 1300 5960 1309
rect 2504 1275 2556 1284
rect 2504 1241 2513 1275
rect 2513 1241 2547 1275
rect 2547 1241 2556 1275
rect 2504 1232 2556 1241
rect 7656 1232 7708 1284
rect 1216 1164 1268 1216
rect 5724 1164 5776 1216
rect 7380 1207 7432 1216
rect 7380 1173 7389 1207
rect 7389 1173 7423 1207
rect 7423 1173 7432 1207
rect 7380 1164 7432 1173
rect 2582 1062 2634 1114
rect 2646 1062 2698 1114
rect 2710 1062 2762 1114
rect 2774 1062 2826 1114
rect 2838 1062 2890 1114
rect 4307 1062 4359 1114
rect 4371 1062 4423 1114
rect 4435 1062 4487 1114
rect 4499 1062 4551 1114
rect 4563 1062 4615 1114
rect 6032 1062 6084 1114
rect 6096 1062 6148 1114
rect 6160 1062 6212 1114
rect 6224 1062 6276 1114
rect 6288 1062 6340 1114
rect 7757 1062 7809 1114
rect 7821 1062 7873 1114
rect 7885 1062 7937 1114
rect 7949 1062 8001 1114
rect 8013 1062 8065 1114
rect 2412 960 2464 1012
rect 2596 960 2648 1012
<< metal2 >>
rect 754 9330 810 10000
rect 754 9302 980 9330
rect 754 9200 810 9302
rect 952 8362 980 9302
rect 1030 9200 1086 10000
rect 1306 9200 1362 10000
rect 1582 9330 1638 10000
rect 1412 9302 1638 9330
rect 940 8356 992 8362
rect 940 8298 992 8304
rect 1044 6390 1072 9200
rect 1320 7818 1348 9200
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 1214 7712 1270 7721
rect 1214 7647 1270 7656
rect 1032 6384 1084 6390
rect 1032 6326 1084 6332
rect 756 4480 808 4486
rect 756 4422 808 4428
rect 296 4004 348 4010
rect 296 3946 348 3952
rect 308 800 336 3946
rect 768 800 796 4422
rect 1228 2514 1256 7647
rect 1320 7546 1348 7754
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1412 5710 1440 9302
rect 1582 9200 1638 9302
rect 1858 9200 1914 10000
rect 2134 9200 2190 10000
rect 2410 9200 2466 10000
rect 2686 9330 2742 10000
rect 2516 9302 2742 9330
rect 1872 8634 1900 9200
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 7886 1532 8298
rect 1720 8188 2028 8197
rect 1720 8186 1726 8188
rect 1782 8186 1806 8188
rect 1862 8186 1886 8188
rect 1942 8186 1966 8188
rect 2022 8186 2028 8188
rect 1782 8134 1784 8186
rect 1964 8134 1966 8186
rect 1720 8132 1726 8134
rect 1782 8132 1806 8134
rect 1862 8132 1886 8134
rect 1942 8132 1966 8134
rect 2022 8132 2028 8134
rect 1720 8123 2028 8132
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1504 7002 1532 7822
rect 1720 7100 2028 7109
rect 1720 7098 1726 7100
rect 1782 7098 1806 7100
rect 1862 7098 1886 7100
rect 1942 7098 1966 7100
rect 2022 7098 2028 7100
rect 1782 7046 1784 7098
rect 1964 7046 1966 7098
rect 1720 7044 1726 7046
rect 1782 7044 1806 7046
rect 1862 7044 1886 7046
rect 1942 7044 1966 7046
rect 2022 7044 2028 7046
rect 1582 7032 1638 7041
rect 1720 7035 2028 7044
rect 1492 6996 1544 7002
rect 1582 6967 1584 6976
rect 1492 6938 1544 6944
rect 1636 6967 1638 6976
rect 1584 6938 1636 6944
rect 1720 6012 2028 6021
rect 1720 6010 1726 6012
rect 1782 6010 1806 6012
rect 1862 6010 1886 6012
rect 1942 6010 1966 6012
rect 2022 6010 2028 6012
rect 1782 5958 1784 6010
rect 1964 5958 1966 6010
rect 1720 5956 1726 5958
rect 1782 5956 1806 5958
rect 1862 5956 1886 5958
rect 1942 5956 1966 5958
rect 2022 5956 2028 5958
rect 1720 5947 2028 5956
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 2148 5574 2176 9200
rect 2424 8650 2452 9200
rect 2332 8622 2452 8650
rect 2332 8362 2360 8622
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2424 8401 2452 8434
rect 2410 8392 2466 8401
rect 2320 8356 2372 8362
rect 2410 8327 2466 8336
rect 2320 8298 2372 8304
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 7002 2268 7346
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2424 6914 2452 8327
rect 2332 6886 2452 6914
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4486 1348 5102
rect 1720 4924 2028 4933
rect 1720 4922 1726 4924
rect 1782 4922 1806 4924
rect 1862 4922 1886 4924
rect 1942 4922 1966 4924
rect 2022 4922 2028 4924
rect 1782 4870 1784 4922
rect 1964 4870 1966 4922
rect 1720 4868 1726 4870
rect 1782 4868 1806 4870
rect 1862 4868 1886 4870
rect 1942 4868 1966 4870
rect 2022 4868 2028 4870
rect 1720 4859 2028 4868
rect 1308 4480 1360 4486
rect 1308 4422 1360 4428
rect 2056 3942 2084 5170
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1720 3836 2028 3845
rect 1720 3834 1726 3836
rect 1782 3834 1806 3836
rect 1862 3834 1886 3836
rect 1942 3834 1966 3836
rect 2022 3834 2028 3836
rect 1782 3782 1784 3834
rect 1964 3782 1966 3834
rect 1720 3780 1726 3782
rect 1782 3780 1806 3782
rect 1862 3780 1886 3782
rect 1942 3780 1966 3782
rect 2022 3780 2028 3782
rect 1720 3771 2028 3780
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 3194 1716 3402
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1720 2748 2028 2757
rect 1720 2746 1726 2748
rect 1782 2746 1806 2748
rect 1862 2746 1886 2748
rect 1942 2746 1966 2748
rect 2022 2746 2028 2748
rect 1782 2694 1784 2746
rect 1964 2694 1966 2746
rect 1720 2692 1726 2694
rect 1782 2692 1806 2694
rect 1862 2692 1886 2694
rect 1942 2692 1966 2694
rect 2022 2692 2028 2694
rect 1720 2683 2028 2692
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 1596 2106 1624 2314
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1720 1660 2028 1669
rect 1720 1658 1726 1660
rect 1782 1658 1806 1660
rect 1862 1658 1886 1660
rect 1942 1658 1966 1660
rect 2022 1658 2028 1660
rect 1782 1606 1784 1658
rect 1964 1606 1966 1658
rect 1720 1604 1726 1606
rect 1782 1604 1806 1606
rect 1862 1604 1886 1606
rect 1942 1604 1966 1606
rect 2022 1604 2028 1606
rect 1720 1595 2028 1604
rect 1216 1216 1268 1222
rect 1216 1158 1268 1164
rect 1228 800 1256 1158
rect 1688 870 1808 898
rect 1688 800 1716 870
rect 294 0 350 800
rect 754 0 810 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 1780 762 1808 870
rect 2056 762 2084 3674
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2148 800 2176 3470
rect 2332 2106 2360 6886
rect 2516 4690 2544 9302
rect 2686 9200 2742 9302
rect 2962 9200 3018 10000
rect 3238 9330 3294 10000
rect 3160 9302 3294 9330
rect 2582 8732 2890 8741
rect 2582 8730 2588 8732
rect 2644 8730 2668 8732
rect 2724 8730 2748 8732
rect 2804 8730 2828 8732
rect 2884 8730 2890 8732
rect 2644 8678 2646 8730
rect 2826 8678 2828 8730
rect 2582 8676 2588 8678
rect 2644 8676 2668 8678
rect 2724 8676 2748 8678
rect 2804 8676 2828 8678
rect 2884 8676 2890 8678
rect 2582 8667 2890 8676
rect 2976 8090 3004 9200
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2582 7644 2890 7653
rect 2582 7642 2588 7644
rect 2644 7642 2668 7644
rect 2724 7642 2748 7644
rect 2804 7642 2828 7644
rect 2884 7642 2890 7644
rect 2644 7590 2646 7642
rect 2826 7590 2828 7642
rect 2582 7588 2588 7590
rect 2644 7588 2668 7590
rect 2724 7588 2748 7590
rect 2804 7588 2828 7590
rect 2884 7588 2890 7590
rect 2582 7579 2890 7588
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2582 6556 2890 6565
rect 2582 6554 2588 6556
rect 2644 6554 2668 6556
rect 2724 6554 2748 6556
rect 2804 6554 2828 6556
rect 2884 6554 2890 6556
rect 2644 6502 2646 6554
rect 2826 6502 2828 6554
rect 2582 6500 2588 6502
rect 2644 6500 2668 6502
rect 2724 6500 2748 6502
rect 2804 6500 2828 6502
rect 2884 6500 2890 6502
rect 2582 6491 2890 6500
rect 3068 6254 3096 6598
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2582 5468 2890 5477
rect 2582 5466 2588 5468
rect 2644 5466 2668 5468
rect 2724 5466 2748 5468
rect 2804 5466 2828 5468
rect 2884 5466 2890 5468
rect 2644 5414 2646 5466
rect 2826 5414 2828 5466
rect 2582 5412 2588 5414
rect 2644 5412 2668 5414
rect 2724 5412 2748 5414
rect 2804 5412 2828 5414
rect 2884 5412 2890 5414
rect 2582 5403 2890 5412
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2582 4380 2890 4389
rect 2582 4378 2588 4380
rect 2644 4378 2668 4380
rect 2724 4378 2748 4380
rect 2804 4378 2828 4380
rect 2884 4378 2890 4380
rect 2644 4326 2646 4378
rect 2826 4326 2828 4378
rect 2582 4324 2588 4326
rect 2644 4324 2668 4326
rect 2724 4324 2748 4326
rect 2804 4324 2828 4326
rect 2884 4324 2890 4326
rect 2582 4315 2890 4324
rect 2976 4146 3004 5510
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3068 3602 3096 5646
rect 3160 5302 3188 9302
rect 3238 9200 3294 9302
rect 3514 9330 3570 10000
rect 3514 9302 3740 9330
rect 3514 9200 3570 9302
rect 3330 9072 3386 9081
rect 3330 9007 3386 9016
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3252 6662 3280 7346
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 5681 3280 6598
rect 3238 5672 3294 5681
rect 3238 5607 3294 5616
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3160 3398 3188 4490
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 2582 3292 2890 3301
rect 2582 3290 2588 3292
rect 2644 3290 2668 3292
rect 2724 3290 2748 3292
rect 2804 3290 2828 3292
rect 2884 3290 2890 3292
rect 2644 3238 2646 3290
rect 2826 3238 2828 3290
rect 2582 3236 2588 3238
rect 2644 3236 2668 3238
rect 2724 3236 2748 3238
rect 2804 3236 2828 3238
rect 2884 3236 2890 3238
rect 2582 3227 2890 3236
rect 3160 3194 3188 3334
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 2962 2952 3018 2961
rect 2962 2887 3018 2896
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 2424 1018 2452 2790
rect 2582 2204 2890 2213
rect 2582 2202 2588 2204
rect 2644 2202 2668 2204
rect 2724 2202 2748 2204
rect 2804 2202 2828 2204
rect 2884 2202 2890 2204
rect 2644 2150 2646 2202
rect 2826 2150 2828 2202
rect 2582 2148 2588 2150
rect 2644 2148 2668 2150
rect 2724 2148 2748 2150
rect 2804 2148 2828 2150
rect 2884 2148 2890 2150
rect 2582 2139 2890 2148
rect 2976 2038 3004 2887
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3160 2650 3188 2790
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 2964 2032 3016 2038
rect 2964 1974 3016 1980
rect 2504 1284 2556 1290
rect 2504 1226 2556 1232
rect 2412 1012 2464 1018
rect 2412 954 2464 960
rect 2516 921 2544 1226
rect 2582 1116 2890 1125
rect 2582 1114 2588 1116
rect 2644 1114 2668 1116
rect 2724 1114 2748 1116
rect 2804 1114 2828 1116
rect 2884 1114 2890 1116
rect 2644 1062 2646 1114
rect 2826 1062 2828 1114
rect 2582 1060 2588 1062
rect 2644 1060 2668 1062
rect 2724 1060 2748 1062
rect 2804 1060 2828 1062
rect 2884 1060 2890 1062
rect 2582 1051 2890 1060
rect 2596 1012 2648 1018
rect 2596 954 2648 960
rect 2502 912 2558 921
rect 2502 847 2558 856
rect 2608 800 2636 954
rect 3068 800 3096 2246
rect 3252 1873 3280 4422
rect 3344 3058 3372 9007
rect 3712 8634 3740 9302
rect 3790 9200 3846 10000
rect 4066 9200 4122 10000
rect 4342 9330 4398 10000
rect 4172 9302 4398 9330
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3445 8188 3753 8197
rect 3445 8186 3451 8188
rect 3507 8186 3531 8188
rect 3587 8186 3611 8188
rect 3667 8186 3691 8188
rect 3747 8186 3753 8188
rect 3507 8134 3509 8186
rect 3689 8134 3691 8186
rect 3445 8132 3451 8134
rect 3507 8132 3531 8134
rect 3587 8132 3611 8134
rect 3667 8132 3691 8134
rect 3747 8132 3753 8134
rect 3445 8123 3753 8132
rect 3445 7100 3753 7109
rect 3445 7098 3451 7100
rect 3507 7098 3531 7100
rect 3587 7098 3611 7100
rect 3667 7098 3691 7100
rect 3747 7098 3753 7100
rect 3507 7046 3509 7098
rect 3689 7046 3691 7098
rect 3445 7044 3451 7046
rect 3507 7044 3531 7046
rect 3587 7044 3611 7046
rect 3667 7044 3691 7046
rect 3747 7044 3753 7046
rect 3445 7035 3753 7044
rect 3804 6390 3832 9200
rect 4080 8906 4108 9200
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3884 8492 3936 8498
rect 4172 8480 4200 9302
rect 4342 9200 4398 9302
rect 4618 9330 4674 10000
rect 4618 9302 4844 9330
rect 4618 9200 4674 9302
rect 4307 8732 4615 8741
rect 4307 8730 4313 8732
rect 4369 8730 4393 8732
rect 4449 8730 4473 8732
rect 4529 8730 4553 8732
rect 4609 8730 4615 8732
rect 4369 8678 4371 8730
rect 4551 8678 4553 8730
rect 4307 8676 4313 8678
rect 4369 8676 4393 8678
rect 4449 8676 4473 8678
rect 4529 8676 4553 8678
rect 4609 8676 4615 8678
rect 4307 8667 4615 8676
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 3884 8434 3936 8440
rect 3988 8452 4200 8480
rect 3896 8090 3924 8434
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 6746 4016 8452
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 7886 4108 8298
rect 4068 7880 4120 7886
rect 4264 7857 4292 8366
rect 4068 7822 4120 7828
rect 4250 7848 4306 7857
rect 4160 7812 4212 7818
rect 4250 7783 4306 7792
rect 4160 7754 4212 7760
rect 4172 7313 4200 7754
rect 4307 7644 4615 7653
rect 4307 7642 4313 7644
rect 4369 7642 4393 7644
rect 4449 7642 4473 7644
rect 4529 7642 4553 7644
rect 4609 7642 4615 7644
rect 4369 7590 4371 7642
rect 4551 7590 4553 7642
rect 4307 7588 4313 7590
rect 4369 7588 4393 7590
rect 4449 7588 4473 7590
rect 4529 7588 4553 7590
rect 4609 7588 4615 7590
rect 4307 7579 4615 7588
rect 4724 7478 4752 8570
rect 4816 8022 4844 9302
rect 4894 9200 4950 10000
rect 5170 9200 5226 10000
rect 5446 9200 5502 10000
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4158 7304 4214 7313
rect 4158 7239 4214 7248
rect 4816 6769 4844 7754
rect 4802 6760 4858 6769
rect 3988 6718 4108 6746
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3988 6322 4016 6598
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3445 6012 3753 6021
rect 3445 6010 3451 6012
rect 3507 6010 3531 6012
rect 3587 6010 3611 6012
rect 3667 6010 3691 6012
rect 3747 6010 3753 6012
rect 3507 5958 3509 6010
rect 3689 5958 3691 6010
rect 3445 5956 3451 5958
rect 3507 5956 3531 5958
rect 3587 5956 3611 5958
rect 3667 5956 3691 5958
rect 3747 5956 3753 5958
rect 3445 5947 3753 5956
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3445 4924 3753 4933
rect 3445 4922 3451 4924
rect 3507 4922 3531 4924
rect 3587 4922 3611 4924
rect 3667 4922 3691 4924
rect 3747 4922 3753 4924
rect 3507 4870 3509 4922
rect 3689 4870 3691 4922
rect 3445 4868 3451 4870
rect 3507 4868 3531 4870
rect 3587 4868 3611 4870
rect 3667 4868 3691 4870
rect 3747 4868 3753 4870
rect 3445 4859 3753 4868
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3620 4185 3648 4218
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3712 4078 3740 4762
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3445 3836 3753 3845
rect 3445 3834 3451 3836
rect 3507 3834 3531 3836
rect 3587 3834 3611 3836
rect 3667 3834 3691 3836
rect 3747 3834 3753 3836
rect 3507 3782 3509 3834
rect 3689 3782 3691 3834
rect 3445 3780 3451 3782
rect 3507 3780 3531 3782
rect 3587 3780 3611 3782
rect 3667 3780 3691 3782
rect 3747 3780 3753 3782
rect 3445 3771 3753 3780
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3804 2774 3832 5578
rect 3896 4826 3924 6190
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3882 4720 3938 4729
rect 3882 4655 3938 4664
rect 3896 3466 3924 4655
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 3445 2748 3753 2757
rect 3445 2746 3451 2748
rect 3507 2746 3531 2748
rect 3587 2746 3611 2748
rect 3667 2746 3691 2748
rect 3747 2746 3753 2748
rect 3804 2746 3924 2774
rect 3507 2694 3509 2746
rect 3689 2694 3691 2746
rect 3445 2692 3451 2694
rect 3507 2692 3531 2694
rect 3587 2692 3611 2694
rect 3667 2692 3691 2694
rect 3747 2692 3753 2694
rect 3445 2683 3753 2692
rect 3792 2576 3844 2582
rect 3792 2518 3844 2524
rect 3330 2408 3386 2417
rect 3330 2343 3386 2352
rect 3344 2038 3372 2343
rect 3804 2310 3832 2518
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3332 2032 3384 2038
rect 3332 1974 3384 1980
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3238 1864 3294 1873
rect 3238 1799 3294 1808
rect 3445 1660 3753 1669
rect 3445 1658 3451 1660
rect 3507 1658 3531 1660
rect 3587 1658 3611 1660
rect 3667 1658 3691 1660
rect 3747 1658 3753 1660
rect 3507 1606 3509 1658
rect 3689 1606 3691 1658
rect 3445 1604 3451 1606
rect 3507 1604 3531 1606
rect 3587 1604 3611 1606
rect 3667 1604 3691 1606
rect 3747 1604 3753 1606
rect 3445 1595 3753 1604
rect 3804 1562 3832 1906
rect 3792 1556 3844 1562
rect 3792 1498 3844 1504
rect 3528 870 3648 898
rect 3528 800 3556 870
rect 1780 734 2084 762
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3620 762 3648 870
rect 3896 762 3924 2746
rect 3988 800 4016 6258
rect 4080 5778 4108 6718
rect 4802 6695 4858 6704
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4307 6556 4615 6565
rect 4307 6554 4313 6556
rect 4369 6554 4393 6556
rect 4449 6554 4473 6556
rect 4529 6554 4553 6556
rect 4609 6554 4615 6556
rect 4369 6502 4371 6554
rect 4551 6502 4553 6554
rect 4307 6500 4313 6502
rect 4369 6500 4393 6502
rect 4449 6500 4473 6502
rect 4529 6500 4553 6502
rect 4609 6500 4615 6502
rect 4307 6491 4615 6500
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4264 5658 4292 6258
rect 4172 5630 4292 5658
rect 4712 5636 4764 5642
rect 4172 5574 4200 5630
rect 4712 5578 4764 5584
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5386 4200 5510
rect 4307 5468 4615 5477
rect 4307 5466 4313 5468
rect 4369 5466 4393 5468
rect 4449 5466 4473 5468
rect 4529 5466 4553 5468
rect 4609 5466 4615 5468
rect 4369 5414 4371 5466
rect 4551 5414 4553 5466
rect 4307 5412 4313 5414
rect 4369 5412 4393 5414
rect 4449 5412 4473 5414
rect 4529 5412 4553 5414
rect 4609 5412 4615 5414
rect 4307 5403 4615 5412
rect 4080 5358 4200 5386
rect 4080 3641 4108 5358
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4172 4264 4200 5170
rect 4724 4486 4752 5578
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4307 4380 4615 4389
rect 4307 4378 4313 4380
rect 4369 4378 4393 4380
rect 4449 4378 4473 4380
rect 4529 4378 4553 4380
rect 4609 4378 4615 4380
rect 4369 4326 4371 4378
rect 4551 4326 4553 4378
rect 4307 4324 4313 4326
rect 4369 4324 4393 4326
rect 4449 4324 4473 4326
rect 4529 4324 4553 4326
rect 4609 4324 4615 4326
rect 4307 4315 4615 4324
rect 4816 4298 4844 6598
rect 4724 4270 4844 4298
rect 4172 4236 4292 4264
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4066 3632 4122 3641
rect 4066 3567 4122 3576
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 1970 4108 3402
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 3620 734 3924 762
rect 3974 0 4030 800
rect 4172 762 4200 3878
rect 4264 3738 4292 4236
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4724 3641 4752 4270
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4710 3632 4766 3641
rect 4710 3567 4766 3576
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4307 3292 4615 3301
rect 4307 3290 4313 3292
rect 4369 3290 4393 3292
rect 4449 3290 4473 3292
rect 4529 3290 4553 3292
rect 4609 3290 4615 3292
rect 4369 3238 4371 3290
rect 4551 3238 4553 3290
rect 4307 3236 4313 3238
rect 4369 3236 4393 3238
rect 4449 3236 4473 3238
rect 4529 3236 4553 3238
rect 4609 3236 4615 3238
rect 4307 3227 4615 3236
rect 4724 3194 4752 3402
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4710 3088 4766 3097
rect 4816 3058 4844 4150
rect 4710 3023 4766 3032
rect 4804 3052 4856 3058
rect 4307 2204 4615 2213
rect 4307 2202 4313 2204
rect 4369 2202 4393 2204
rect 4449 2202 4473 2204
rect 4529 2202 4553 2204
rect 4609 2202 4615 2204
rect 4369 2150 4371 2202
rect 4551 2150 4553 2202
rect 4307 2148 4313 2150
rect 4369 2148 4393 2150
rect 4449 2148 4473 2150
rect 4529 2148 4553 2150
rect 4609 2148 4615 2150
rect 4307 2139 4615 2148
rect 4724 1426 4752 3023
rect 4804 2994 4856 3000
rect 4908 2514 4936 9200
rect 5184 8838 5212 9200
rect 5460 8922 5488 9200
rect 5276 8894 5488 8922
rect 5540 8900 5592 8906
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5276 8344 5304 8894
rect 5540 8842 5592 8848
rect 5092 8316 5304 8344
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6730 5028 7142
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 5092 3126 5120 8316
rect 5170 8188 5478 8197
rect 5170 8186 5176 8188
rect 5232 8186 5256 8188
rect 5312 8186 5336 8188
rect 5392 8186 5416 8188
rect 5472 8186 5478 8188
rect 5232 8134 5234 8186
rect 5414 8134 5416 8186
rect 5170 8132 5176 8134
rect 5232 8132 5256 8134
rect 5312 8132 5336 8134
rect 5392 8132 5416 8134
rect 5472 8132 5478 8134
rect 5170 8123 5478 8132
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5354 7984 5410 7993
rect 5184 7206 5212 7958
rect 5354 7919 5410 7928
rect 5368 7546 5396 7919
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5552 7478 5580 8842
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5170 7100 5478 7109
rect 5170 7098 5176 7100
rect 5232 7098 5256 7100
rect 5312 7098 5336 7100
rect 5392 7098 5416 7100
rect 5472 7098 5478 7100
rect 5232 7046 5234 7098
rect 5414 7046 5416 7098
rect 5170 7044 5176 7046
rect 5232 7044 5256 7046
rect 5312 7044 5336 7046
rect 5392 7044 5416 7046
rect 5472 7044 5478 7046
rect 5170 7035 5478 7044
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 6390 5304 6598
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5170 6012 5478 6021
rect 5170 6010 5176 6012
rect 5232 6010 5256 6012
rect 5312 6010 5336 6012
rect 5392 6010 5416 6012
rect 5472 6010 5478 6012
rect 5232 5958 5234 6010
rect 5414 5958 5416 6010
rect 5170 5956 5176 5958
rect 5232 5956 5256 5958
rect 5312 5956 5336 5958
rect 5392 5956 5416 5958
rect 5472 5956 5478 5958
rect 5170 5947 5478 5956
rect 5446 5808 5502 5817
rect 5446 5743 5448 5752
rect 5500 5743 5502 5752
rect 5448 5714 5500 5720
rect 5552 5137 5580 7278
rect 5644 5302 5672 9386
rect 5722 9200 5778 10000
rect 5998 9330 6054 10000
rect 5828 9302 6054 9330
rect 5736 6798 5764 9200
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6458 5764 6734
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5538 5128 5594 5137
rect 5538 5063 5594 5072
rect 5170 4924 5478 4933
rect 5170 4922 5176 4924
rect 5232 4922 5256 4924
rect 5312 4922 5336 4924
rect 5392 4922 5416 4924
rect 5472 4922 5478 4924
rect 5232 4870 5234 4922
rect 5414 4870 5416 4922
rect 5170 4868 5176 4870
rect 5232 4868 5256 4870
rect 5312 4868 5336 4870
rect 5392 4868 5416 4870
rect 5472 4868 5478 4870
rect 5170 4859 5478 4868
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5460 4146 5488 4762
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5170 3836 5478 3845
rect 5170 3834 5176 3836
rect 5232 3834 5256 3836
rect 5312 3834 5336 3836
rect 5392 3834 5416 3836
rect 5472 3834 5478 3836
rect 5232 3782 5234 3834
rect 5414 3782 5416 3834
rect 5170 3780 5176 3782
rect 5232 3780 5256 3782
rect 5312 3780 5336 3782
rect 5392 3780 5416 3782
rect 5472 3780 5478 3782
rect 5170 3771 5478 3780
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 5000 2394 5028 2926
rect 4908 2366 5028 2394
rect 4712 1420 4764 1426
rect 4712 1362 4764 1368
rect 4307 1116 4615 1125
rect 4307 1114 4313 1116
rect 4369 1114 4393 1116
rect 4449 1114 4473 1116
rect 4529 1114 4553 1116
rect 4609 1114 4615 1116
rect 4369 1062 4371 1114
rect 4551 1062 4553 1114
rect 4307 1060 4313 1062
rect 4369 1060 4393 1062
rect 4449 1060 4473 1062
rect 4529 1060 4553 1062
rect 4609 1060 4615 1062
rect 4307 1051 4615 1060
rect 4356 870 4476 898
rect 4356 762 4384 870
rect 4448 800 4476 870
rect 4908 800 4936 2366
rect 4172 734 4384 762
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5092 762 5120 2926
rect 5170 2748 5478 2757
rect 5170 2746 5176 2748
rect 5232 2746 5256 2748
rect 5312 2746 5336 2748
rect 5392 2746 5416 2748
rect 5472 2746 5478 2748
rect 5232 2694 5234 2746
rect 5414 2694 5416 2746
rect 5170 2692 5176 2694
rect 5232 2692 5256 2694
rect 5312 2692 5336 2694
rect 5392 2692 5416 2694
rect 5472 2692 5478 2694
rect 5170 2683 5478 2692
rect 5552 2514 5580 4218
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5644 3126 5672 4014
rect 5736 3466 5764 4490
rect 5828 3602 5856 9302
rect 5998 9200 6054 9302
rect 6274 9330 6330 10000
rect 6550 9466 6606 10000
rect 6380 9450 6606 9466
rect 6368 9444 6606 9450
rect 6420 9438 6606 9444
rect 6368 9386 6420 9392
rect 6274 9302 6500 9330
rect 6274 9200 6330 9302
rect 6032 8732 6340 8741
rect 6032 8730 6038 8732
rect 6094 8730 6118 8732
rect 6174 8730 6198 8732
rect 6254 8730 6278 8732
rect 6334 8730 6340 8732
rect 6094 8678 6096 8730
rect 6276 8678 6278 8730
rect 6032 8676 6038 8678
rect 6094 8676 6118 8678
rect 6174 8676 6198 8678
rect 6254 8676 6278 8678
rect 6334 8676 6340 8678
rect 6032 8667 6340 8676
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5920 6361 5948 8366
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6032 7644 6340 7653
rect 6032 7642 6038 7644
rect 6094 7642 6118 7644
rect 6174 7642 6198 7644
rect 6254 7642 6278 7644
rect 6334 7642 6340 7644
rect 6094 7590 6096 7642
rect 6276 7590 6278 7642
rect 6032 7588 6038 7590
rect 6094 7588 6118 7590
rect 6174 7588 6198 7590
rect 6254 7588 6278 7590
rect 6334 7588 6340 7590
rect 6032 7579 6340 7588
rect 6032 6556 6340 6565
rect 6032 6554 6038 6556
rect 6094 6554 6118 6556
rect 6174 6554 6198 6556
rect 6254 6554 6278 6556
rect 6334 6554 6340 6556
rect 6094 6502 6096 6554
rect 6276 6502 6278 6554
rect 6032 6500 6038 6502
rect 6094 6500 6118 6502
rect 6174 6500 6198 6502
rect 6254 6500 6278 6502
rect 6334 6500 6340 6502
rect 6032 6491 6340 6500
rect 5906 6352 5962 6361
rect 5906 6287 5962 6296
rect 6380 6225 6408 7754
rect 6366 6216 6422 6225
rect 6366 6151 6422 6160
rect 6472 5710 6500 9302
rect 6550 9200 6606 9438
rect 6826 9330 6882 10000
rect 6748 9302 6882 9330
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6550 8392 6606 8401
rect 6550 8327 6606 8336
rect 6564 7410 6592 8327
rect 6656 8090 6684 8774
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 5920 4146 5948 5646
rect 6032 5468 6340 5477
rect 6032 5466 6038 5468
rect 6094 5466 6118 5468
rect 6174 5466 6198 5468
rect 6254 5466 6278 5468
rect 6334 5466 6340 5468
rect 6094 5414 6096 5466
rect 6276 5414 6278 5466
rect 6032 5412 6038 5414
rect 6094 5412 6118 5414
rect 6174 5412 6198 5414
rect 6254 5412 6278 5414
rect 6334 5412 6340 5414
rect 6032 5403 6340 5412
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6032 4380 6340 4389
rect 6032 4378 6038 4380
rect 6094 4378 6118 4380
rect 6174 4378 6198 4380
rect 6254 4378 6278 4380
rect 6334 4378 6340 4380
rect 6094 4326 6096 4378
rect 6276 4326 6278 4378
rect 6032 4324 6038 4326
rect 6094 4324 6118 4326
rect 6174 4324 6198 4326
rect 6254 4324 6278 4326
rect 6334 4324 6340 4326
rect 6032 4315 6340 4324
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5170 1660 5478 1669
rect 5170 1658 5176 1660
rect 5232 1658 5256 1660
rect 5312 1658 5336 1660
rect 5392 1658 5416 1660
rect 5472 1658 5478 1660
rect 5232 1606 5234 1658
rect 5414 1606 5416 1658
rect 5170 1604 5176 1606
rect 5232 1604 5256 1606
rect 5312 1604 5336 1606
rect 5392 1604 5416 1606
rect 5472 1604 5478 1606
rect 5170 1595 5478 1604
rect 5736 1222 5764 3402
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5724 1216 5776 1222
rect 5724 1158 5776 1164
rect 5276 870 5396 898
rect 5276 762 5304 870
rect 5368 800 5396 870
rect 5828 800 5856 3334
rect 6032 3292 6340 3301
rect 6032 3290 6038 3292
rect 6094 3290 6118 3292
rect 6174 3290 6198 3292
rect 6254 3290 6278 3292
rect 6334 3290 6340 3292
rect 6094 3238 6096 3290
rect 6276 3238 6278 3290
rect 6032 3236 6038 3238
rect 6094 3236 6118 3238
rect 6174 3236 6198 3238
rect 6254 3236 6278 3238
rect 6334 3236 6340 3238
rect 6032 3227 6340 3236
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6288 2394 6316 3062
rect 6380 2553 6408 5102
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6366 2544 6422 2553
rect 6366 2479 6422 2488
rect 6472 2417 6500 4490
rect 6564 4185 6592 6666
rect 6656 6390 6684 8026
rect 6748 6390 6776 9302
rect 6826 9200 6882 9302
rect 7102 9330 7158 10000
rect 7102 9302 7328 9330
rect 7102 9200 7158 9302
rect 6895 8188 7203 8197
rect 6895 8186 6901 8188
rect 6957 8186 6981 8188
rect 7037 8186 7061 8188
rect 7117 8186 7141 8188
rect 7197 8186 7203 8188
rect 6957 8134 6959 8186
rect 7139 8134 7141 8186
rect 6895 8132 6901 8134
rect 6957 8132 6981 8134
rect 7037 8132 7061 8134
rect 7117 8132 7141 8134
rect 7197 8132 7203 8134
rect 6895 8123 7203 8132
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 7478 7236 7686
rect 7300 7478 7328 9302
rect 7378 9200 7434 10000
rect 7654 9466 7710 10000
rect 7654 9450 7880 9466
rect 7654 9444 7892 9450
rect 7654 9438 7840 9444
rect 7654 9200 7710 9438
rect 7840 9386 7892 9392
rect 7930 9330 7986 10000
rect 7760 9302 7986 9330
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 6895 7100 7203 7109
rect 6895 7098 6901 7100
rect 6957 7098 6981 7100
rect 7037 7098 7061 7100
rect 7117 7098 7141 7100
rect 7197 7098 7203 7100
rect 6957 7046 6959 7098
rect 7139 7046 7141 7098
rect 6895 7044 6901 7046
rect 6957 7044 6981 7046
rect 7037 7044 7061 7046
rect 7117 7044 7141 7046
rect 7197 7044 7203 7046
rect 6895 7035 7203 7044
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6550 4176 6606 4185
rect 6550 4111 6606 4120
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6458 2408 6514 2417
rect 6288 2366 6408 2394
rect 6032 2204 6340 2213
rect 6032 2202 6038 2204
rect 6094 2202 6118 2204
rect 6174 2202 6198 2204
rect 6254 2202 6278 2204
rect 6334 2202 6340 2204
rect 6094 2150 6096 2202
rect 6276 2150 6278 2202
rect 6032 2148 6038 2150
rect 6094 2148 6118 2150
rect 6174 2148 6198 2150
rect 6254 2148 6278 2150
rect 6334 2148 6340 2150
rect 6032 2139 6340 2148
rect 5906 1456 5962 1465
rect 5906 1391 5962 1400
rect 5920 1358 5948 1391
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 6032 1116 6340 1125
rect 6032 1114 6038 1116
rect 6094 1114 6118 1116
rect 6174 1114 6198 1116
rect 6254 1114 6278 1116
rect 6334 1114 6340 1116
rect 6094 1062 6096 1114
rect 6276 1062 6278 1114
rect 6032 1060 6038 1062
rect 6094 1060 6118 1062
rect 6174 1060 6198 1062
rect 6254 1060 6278 1062
rect 6334 1060 6340 1062
rect 6032 1051 6340 1060
rect 6380 898 6408 2366
rect 6458 2343 6514 2352
rect 6564 1873 6592 4014
rect 6656 3097 6684 5578
rect 6748 4049 6776 6190
rect 6895 6012 7203 6021
rect 6895 6010 6901 6012
rect 6957 6010 6981 6012
rect 7037 6010 7061 6012
rect 7117 6010 7141 6012
rect 7197 6010 7203 6012
rect 6957 5958 6959 6010
rect 7139 5958 7141 6010
rect 6895 5956 6901 5958
rect 6957 5956 6981 5958
rect 7037 5956 7061 5958
rect 7117 5956 7141 5958
rect 7197 5956 7203 5958
rect 6895 5947 7203 5956
rect 6895 4924 7203 4933
rect 6895 4922 6901 4924
rect 6957 4922 6981 4924
rect 7037 4922 7061 4924
rect 7117 4922 7141 4924
rect 7197 4922 7203 4924
rect 6957 4870 6959 4922
rect 7139 4870 7141 4922
rect 6895 4868 6901 4870
rect 6957 4868 6981 4870
rect 7037 4868 7061 4870
rect 7117 4868 7141 4870
rect 7197 4868 7203 4870
rect 6895 4859 7203 4868
rect 7300 4729 7328 7278
rect 7392 6474 7420 9200
rect 7470 8936 7526 8945
rect 7760 8922 7788 9302
rect 7930 9200 7986 9302
rect 8206 9200 8262 10000
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 7470 8871 7526 8880
rect 7668 8894 7788 8922
rect 7484 6662 7512 8871
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7392 6446 7512 6474
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7392 5302 7420 6326
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7286 4720 7342 4729
rect 7286 4655 7342 4664
rect 6734 4040 6790 4049
rect 6734 3975 6790 3984
rect 6895 3836 7203 3845
rect 6895 3834 6901 3836
rect 6957 3834 6981 3836
rect 7037 3834 7061 3836
rect 7117 3834 7141 3836
rect 7197 3834 7203 3836
rect 6957 3782 6959 3834
rect 7139 3782 7141 3834
rect 6895 3780 6901 3782
rect 6957 3780 6981 3782
rect 7037 3780 7061 3782
rect 7117 3780 7141 3782
rect 7197 3780 7203 3782
rect 6895 3771 7203 3780
rect 7392 3738 7420 5238
rect 7484 4622 7512 6446
rect 7576 4690 7604 7414
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7484 3670 7512 4558
rect 7668 4214 7696 8894
rect 7757 8732 8065 8741
rect 7757 8730 7763 8732
rect 7819 8730 7843 8732
rect 7899 8730 7923 8732
rect 7979 8730 8003 8732
rect 8059 8730 8065 8732
rect 7819 8678 7821 8730
rect 8001 8678 8003 8730
rect 7757 8676 7763 8678
rect 7819 8676 7843 8678
rect 7899 8676 7923 8678
rect 7979 8676 8003 8678
rect 8059 8676 8065 8678
rect 7757 8667 8065 8676
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7757 7644 8065 7653
rect 7757 7642 7763 7644
rect 7819 7642 7843 7644
rect 7899 7642 7923 7644
rect 7979 7642 8003 7644
rect 8059 7642 8065 7644
rect 7819 7590 7821 7642
rect 8001 7590 8003 7642
rect 7757 7588 7763 7590
rect 7819 7588 7843 7590
rect 7899 7588 7923 7590
rect 7979 7588 8003 7590
rect 8059 7588 8065 7590
rect 7757 7579 8065 7588
rect 7757 6556 8065 6565
rect 7757 6554 7763 6556
rect 7819 6554 7843 6556
rect 7899 6554 7923 6556
rect 7979 6554 8003 6556
rect 8059 6554 8065 6556
rect 7819 6502 7821 6554
rect 8001 6502 8003 6554
rect 7757 6500 7763 6502
rect 7819 6500 7843 6502
rect 7899 6500 7923 6502
rect 7979 6500 8003 6502
rect 8059 6500 8065 6502
rect 7757 6491 8065 6500
rect 8022 5672 8078 5681
rect 8128 5658 8156 8366
rect 8078 5630 8156 5658
rect 8022 5607 8078 5616
rect 7757 5468 8065 5477
rect 7757 5466 7763 5468
rect 7819 5466 7843 5468
rect 7899 5466 7923 5468
rect 7979 5466 8003 5468
rect 8059 5466 8065 5468
rect 7819 5414 7821 5466
rect 8001 5414 8003 5466
rect 7757 5412 7763 5414
rect 7819 5412 7843 5414
rect 7899 5412 7923 5414
rect 7979 5412 8003 5414
rect 8059 5412 8065 5414
rect 7757 5403 8065 5412
rect 8220 4826 8248 9200
rect 8312 5370 8340 9386
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 7757 4380 8065 4389
rect 7757 4378 7763 4380
rect 7819 4378 7843 4380
rect 7899 4378 7923 4380
rect 7979 4378 8003 4380
rect 8059 4378 8065 4380
rect 7819 4326 7821 4378
rect 8001 4326 8003 4378
rect 7757 4324 7763 4326
rect 7819 4324 7843 4326
rect 7899 4324 7923 4326
rect 7979 4324 8003 4326
rect 8059 4324 8065 4326
rect 7757 4315 8065 4324
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7668 3194 7696 4150
rect 7757 3292 8065 3301
rect 7757 3290 7763 3292
rect 7819 3290 7843 3292
rect 7899 3290 7923 3292
rect 7979 3290 8003 3292
rect 8059 3290 8065 3292
rect 7819 3238 7821 3290
rect 8001 3238 8003 3290
rect 7757 3236 7763 3238
rect 7819 3236 7843 3238
rect 7899 3236 7923 3238
rect 7979 3236 8003 3238
rect 8059 3236 8065 3238
rect 7757 3227 8065 3236
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 6642 3088 6698 3097
rect 6642 3023 6698 3032
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6550 1864 6606 1873
rect 6550 1799 6606 1808
rect 6656 1442 6684 2790
rect 6895 2748 7203 2757
rect 6895 2746 6901 2748
rect 6957 2746 6981 2748
rect 7037 2746 7061 2748
rect 7117 2746 7141 2748
rect 7197 2746 7203 2748
rect 6957 2694 6959 2746
rect 7139 2694 7141 2746
rect 6895 2692 6901 2694
rect 6957 2692 6981 2694
rect 7037 2692 7061 2694
rect 7117 2692 7141 2694
rect 7197 2692 7203 2694
rect 6895 2683 7203 2692
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6748 1578 6776 2246
rect 6895 1660 7203 1669
rect 6895 1658 6901 1660
rect 6957 1658 6981 1660
rect 7037 1658 7061 1660
rect 7117 1658 7141 1660
rect 7197 1658 7203 1660
rect 6957 1606 6959 1658
rect 7139 1606 7141 1658
rect 6895 1604 6901 1606
rect 6957 1604 6981 1606
rect 7037 1604 7061 1606
rect 7117 1604 7141 1606
rect 7197 1604 7203 1606
rect 6895 1595 7203 1604
rect 6748 1550 6868 1578
rect 6656 1414 6776 1442
rect 6288 870 6408 898
rect 6288 800 6316 870
rect 6748 800 6776 1414
rect 5092 734 5304 762
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 6840 649 6868 1550
rect 7300 1306 7328 2382
rect 7757 2204 8065 2213
rect 7757 2202 7763 2204
rect 7819 2202 7843 2204
rect 7899 2202 7923 2204
rect 7979 2202 8003 2204
rect 8059 2202 8065 2204
rect 7819 2150 7821 2202
rect 8001 2150 8003 2202
rect 7757 2148 7763 2150
rect 7819 2148 7843 2150
rect 7899 2148 7923 2150
rect 7979 2148 8003 2150
rect 8059 2148 8065 2150
rect 7757 2139 8065 2148
rect 7380 1964 7432 1970
rect 7380 1906 7432 1912
rect 7208 1278 7328 1306
rect 7208 800 7236 1278
rect 7392 1222 7420 1906
rect 8116 1760 8168 1766
rect 8116 1702 8168 1708
rect 7656 1284 7708 1290
rect 7656 1226 7708 1232
rect 7380 1216 7432 1222
rect 7380 1158 7432 1164
rect 7392 921 7420 1158
rect 7378 912 7434 921
rect 7378 847 7434 856
rect 7668 800 7696 1226
rect 7757 1116 8065 1125
rect 7757 1114 7763 1116
rect 7819 1114 7843 1116
rect 7899 1114 7923 1116
rect 7979 1114 8003 1116
rect 8059 1114 8065 1116
rect 7819 1062 7821 1114
rect 8001 1062 8003 1114
rect 7757 1060 7763 1062
rect 7819 1060 7843 1062
rect 7899 1060 7923 1062
rect 7979 1060 8003 1062
rect 8059 1060 8065 1062
rect 7757 1051 8065 1060
rect 8128 800 8156 1702
rect 8576 1556 8628 1562
rect 8576 1498 8628 1504
rect 8588 800 8616 1498
rect 6826 640 6882 649
rect 6826 575 6882 584
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
<< via2 >>
rect 1214 7656 1270 7712
rect 1726 8186 1782 8188
rect 1806 8186 1862 8188
rect 1886 8186 1942 8188
rect 1966 8186 2022 8188
rect 1726 8134 1772 8186
rect 1772 8134 1782 8186
rect 1806 8134 1836 8186
rect 1836 8134 1848 8186
rect 1848 8134 1862 8186
rect 1886 8134 1900 8186
rect 1900 8134 1912 8186
rect 1912 8134 1942 8186
rect 1966 8134 1976 8186
rect 1976 8134 2022 8186
rect 1726 8132 1782 8134
rect 1806 8132 1862 8134
rect 1886 8132 1942 8134
rect 1966 8132 2022 8134
rect 1726 7098 1782 7100
rect 1806 7098 1862 7100
rect 1886 7098 1942 7100
rect 1966 7098 2022 7100
rect 1726 7046 1772 7098
rect 1772 7046 1782 7098
rect 1806 7046 1836 7098
rect 1836 7046 1848 7098
rect 1848 7046 1862 7098
rect 1886 7046 1900 7098
rect 1900 7046 1912 7098
rect 1912 7046 1942 7098
rect 1966 7046 1976 7098
rect 1976 7046 2022 7098
rect 1726 7044 1782 7046
rect 1806 7044 1862 7046
rect 1886 7044 1942 7046
rect 1966 7044 2022 7046
rect 1582 6996 1638 7032
rect 1582 6976 1584 6996
rect 1584 6976 1636 6996
rect 1636 6976 1638 6996
rect 1726 6010 1782 6012
rect 1806 6010 1862 6012
rect 1886 6010 1942 6012
rect 1966 6010 2022 6012
rect 1726 5958 1772 6010
rect 1772 5958 1782 6010
rect 1806 5958 1836 6010
rect 1836 5958 1848 6010
rect 1848 5958 1862 6010
rect 1886 5958 1900 6010
rect 1900 5958 1912 6010
rect 1912 5958 1942 6010
rect 1966 5958 1976 6010
rect 1976 5958 2022 6010
rect 1726 5956 1782 5958
rect 1806 5956 1862 5958
rect 1886 5956 1942 5958
rect 1966 5956 2022 5958
rect 2410 8336 2466 8392
rect 1726 4922 1782 4924
rect 1806 4922 1862 4924
rect 1886 4922 1942 4924
rect 1966 4922 2022 4924
rect 1726 4870 1772 4922
rect 1772 4870 1782 4922
rect 1806 4870 1836 4922
rect 1836 4870 1848 4922
rect 1848 4870 1862 4922
rect 1886 4870 1900 4922
rect 1900 4870 1912 4922
rect 1912 4870 1942 4922
rect 1966 4870 1976 4922
rect 1976 4870 2022 4922
rect 1726 4868 1782 4870
rect 1806 4868 1862 4870
rect 1886 4868 1942 4870
rect 1966 4868 2022 4870
rect 1726 3834 1782 3836
rect 1806 3834 1862 3836
rect 1886 3834 1942 3836
rect 1966 3834 2022 3836
rect 1726 3782 1772 3834
rect 1772 3782 1782 3834
rect 1806 3782 1836 3834
rect 1836 3782 1848 3834
rect 1848 3782 1862 3834
rect 1886 3782 1900 3834
rect 1900 3782 1912 3834
rect 1912 3782 1942 3834
rect 1966 3782 1976 3834
rect 1976 3782 2022 3834
rect 1726 3780 1782 3782
rect 1806 3780 1862 3782
rect 1886 3780 1942 3782
rect 1966 3780 2022 3782
rect 1726 2746 1782 2748
rect 1806 2746 1862 2748
rect 1886 2746 1942 2748
rect 1966 2746 2022 2748
rect 1726 2694 1772 2746
rect 1772 2694 1782 2746
rect 1806 2694 1836 2746
rect 1836 2694 1848 2746
rect 1848 2694 1862 2746
rect 1886 2694 1900 2746
rect 1900 2694 1912 2746
rect 1912 2694 1942 2746
rect 1966 2694 1976 2746
rect 1976 2694 2022 2746
rect 1726 2692 1782 2694
rect 1806 2692 1862 2694
rect 1886 2692 1942 2694
rect 1966 2692 2022 2694
rect 1726 1658 1782 1660
rect 1806 1658 1862 1660
rect 1886 1658 1942 1660
rect 1966 1658 2022 1660
rect 1726 1606 1772 1658
rect 1772 1606 1782 1658
rect 1806 1606 1836 1658
rect 1836 1606 1848 1658
rect 1848 1606 1862 1658
rect 1886 1606 1900 1658
rect 1900 1606 1912 1658
rect 1912 1606 1942 1658
rect 1966 1606 1976 1658
rect 1976 1606 2022 1658
rect 1726 1604 1782 1606
rect 1806 1604 1862 1606
rect 1886 1604 1942 1606
rect 1966 1604 2022 1606
rect 2588 8730 2644 8732
rect 2668 8730 2724 8732
rect 2748 8730 2804 8732
rect 2828 8730 2884 8732
rect 2588 8678 2634 8730
rect 2634 8678 2644 8730
rect 2668 8678 2698 8730
rect 2698 8678 2710 8730
rect 2710 8678 2724 8730
rect 2748 8678 2762 8730
rect 2762 8678 2774 8730
rect 2774 8678 2804 8730
rect 2828 8678 2838 8730
rect 2838 8678 2884 8730
rect 2588 8676 2644 8678
rect 2668 8676 2724 8678
rect 2748 8676 2804 8678
rect 2828 8676 2884 8678
rect 2588 7642 2644 7644
rect 2668 7642 2724 7644
rect 2748 7642 2804 7644
rect 2828 7642 2884 7644
rect 2588 7590 2634 7642
rect 2634 7590 2644 7642
rect 2668 7590 2698 7642
rect 2698 7590 2710 7642
rect 2710 7590 2724 7642
rect 2748 7590 2762 7642
rect 2762 7590 2774 7642
rect 2774 7590 2804 7642
rect 2828 7590 2838 7642
rect 2838 7590 2884 7642
rect 2588 7588 2644 7590
rect 2668 7588 2724 7590
rect 2748 7588 2804 7590
rect 2828 7588 2884 7590
rect 2588 6554 2644 6556
rect 2668 6554 2724 6556
rect 2748 6554 2804 6556
rect 2828 6554 2884 6556
rect 2588 6502 2634 6554
rect 2634 6502 2644 6554
rect 2668 6502 2698 6554
rect 2698 6502 2710 6554
rect 2710 6502 2724 6554
rect 2748 6502 2762 6554
rect 2762 6502 2774 6554
rect 2774 6502 2804 6554
rect 2828 6502 2838 6554
rect 2838 6502 2884 6554
rect 2588 6500 2644 6502
rect 2668 6500 2724 6502
rect 2748 6500 2804 6502
rect 2828 6500 2884 6502
rect 2588 5466 2644 5468
rect 2668 5466 2724 5468
rect 2748 5466 2804 5468
rect 2828 5466 2884 5468
rect 2588 5414 2634 5466
rect 2634 5414 2644 5466
rect 2668 5414 2698 5466
rect 2698 5414 2710 5466
rect 2710 5414 2724 5466
rect 2748 5414 2762 5466
rect 2762 5414 2774 5466
rect 2774 5414 2804 5466
rect 2828 5414 2838 5466
rect 2838 5414 2884 5466
rect 2588 5412 2644 5414
rect 2668 5412 2724 5414
rect 2748 5412 2804 5414
rect 2828 5412 2884 5414
rect 2588 4378 2644 4380
rect 2668 4378 2724 4380
rect 2748 4378 2804 4380
rect 2828 4378 2884 4380
rect 2588 4326 2634 4378
rect 2634 4326 2644 4378
rect 2668 4326 2698 4378
rect 2698 4326 2710 4378
rect 2710 4326 2724 4378
rect 2748 4326 2762 4378
rect 2762 4326 2774 4378
rect 2774 4326 2804 4378
rect 2828 4326 2838 4378
rect 2838 4326 2884 4378
rect 2588 4324 2644 4326
rect 2668 4324 2724 4326
rect 2748 4324 2804 4326
rect 2828 4324 2884 4326
rect 3330 9016 3386 9072
rect 3238 5616 3294 5672
rect 2588 3290 2644 3292
rect 2668 3290 2724 3292
rect 2748 3290 2804 3292
rect 2828 3290 2884 3292
rect 2588 3238 2634 3290
rect 2634 3238 2644 3290
rect 2668 3238 2698 3290
rect 2698 3238 2710 3290
rect 2710 3238 2724 3290
rect 2748 3238 2762 3290
rect 2762 3238 2774 3290
rect 2774 3238 2804 3290
rect 2828 3238 2838 3290
rect 2838 3238 2884 3290
rect 2588 3236 2644 3238
rect 2668 3236 2724 3238
rect 2748 3236 2804 3238
rect 2828 3236 2884 3238
rect 2962 2896 3018 2952
rect 2588 2202 2644 2204
rect 2668 2202 2724 2204
rect 2748 2202 2804 2204
rect 2828 2202 2884 2204
rect 2588 2150 2634 2202
rect 2634 2150 2644 2202
rect 2668 2150 2698 2202
rect 2698 2150 2710 2202
rect 2710 2150 2724 2202
rect 2748 2150 2762 2202
rect 2762 2150 2774 2202
rect 2774 2150 2804 2202
rect 2828 2150 2838 2202
rect 2838 2150 2884 2202
rect 2588 2148 2644 2150
rect 2668 2148 2724 2150
rect 2748 2148 2804 2150
rect 2828 2148 2884 2150
rect 2588 1114 2644 1116
rect 2668 1114 2724 1116
rect 2748 1114 2804 1116
rect 2828 1114 2884 1116
rect 2588 1062 2634 1114
rect 2634 1062 2644 1114
rect 2668 1062 2698 1114
rect 2698 1062 2710 1114
rect 2710 1062 2724 1114
rect 2748 1062 2762 1114
rect 2762 1062 2774 1114
rect 2774 1062 2804 1114
rect 2828 1062 2838 1114
rect 2838 1062 2884 1114
rect 2588 1060 2644 1062
rect 2668 1060 2724 1062
rect 2748 1060 2804 1062
rect 2828 1060 2884 1062
rect 2502 856 2558 912
rect 3451 8186 3507 8188
rect 3531 8186 3587 8188
rect 3611 8186 3667 8188
rect 3691 8186 3747 8188
rect 3451 8134 3497 8186
rect 3497 8134 3507 8186
rect 3531 8134 3561 8186
rect 3561 8134 3573 8186
rect 3573 8134 3587 8186
rect 3611 8134 3625 8186
rect 3625 8134 3637 8186
rect 3637 8134 3667 8186
rect 3691 8134 3701 8186
rect 3701 8134 3747 8186
rect 3451 8132 3507 8134
rect 3531 8132 3587 8134
rect 3611 8132 3667 8134
rect 3691 8132 3747 8134
rect 3451 7098 3507 7100
rect 3531 7098 3587 7100
rect 3611 7098 3667 7100
rect 3691 7098 3747 7100
rect 3451 7046 3497 7098
rect 3497 7046 3507 7098
rect 3531 7046 3561 7098
rect 3561 7046 3573 7098
rect 3573 7046 3587 7098
rect 3611 7046 3625 7098
rect 3625 7046 3637 7098
rect 3637 7046 3667 7098
rect 3691 7046 3701 7098
rect 3701 7046 3747 7098
rect 3451 7044 3507 7046
rect 3531 7044 3587 7046
rect 3611 7044 3667 7046
rect 3691 7044 3747 7046
rect 4313 8730 4369 8732
rect 4393 8730 4449 8732
rect 4473 8730 4529 8732
rect 4553 8730 4609 8732
rect 4313 8678 4359 8730
rect 4359 8678 4369 8730
rect 4393 8678 4423 8730
rect 4423 8678 4435 8730
rect 4435 8678 4449 8730
rect 4473 8678 4487 8730
rect 4487 8678 4499 8730
rect 4499 8678 4529 8730
rect 4553 8678 4563 8730
rect 4563 8678 4609 8730
rect 4313 8676 4369 8678
rect 4393 8676 4449 8678
rect 4473 8676 4529 8678
rect 4553 8676 4609 8678
rect 4250 7792 4306 7848
rect 4313 7642 4369 7644
rect 4393 7642 4449 7644
rect 4473 7642 4529 7644
rect 4553 7642 4609 7644
rect 4313 7590 4359 7642
rect 4359 7590 4369 7642
rect 4393 7590 4423 7642
rect 4423 7590 4435 7642
rect 4435 7590 4449 7642
rect 4473 7590 4487 7642
rect 4487 7590 4499 7642
rect 4499 7590 4529 7642
rect 4553 7590 4563 7642
rect 4563 7590 4609 7642
rect 4313 7588 4369 7590
rect 4393 7588 4449 7590
rect 4473 7588 4529 7590
rect 4553 7588 4609 7590
rect 4158 7248 4214 7304
rect 3451 6010 3507 6012
rect 3531 6010 3587 6012
rect 3611 6010 3667 6012
rect 3691 6010 3747 6012
rect 3451 5958 3497 6010
rect 3497 5958 3507 6010
rect 3531 5958 3561 6010
rect 3561 5958 3573 6010
rect 3573 5958 3587 6010
rect 3611 5958 3625 6010
rect 3625 5958 3637 6010
rect 3637 5958 3667 6010
rect 3691 5958 3701 6010
rect 3701 5958 3747 6010
rect 3451 5956 3507 5958
rect 3531 5956 3587 5958
rect 3611 5956 3667 5958
rect 3691 5956 3747 5958
rect 3451 4922 3507 4924
rect 3531 4922 3587 4924
rect 3611 4922 3667 4924
rect 3691 4922 3747 4924
rect 3451 4870 3497 4922
rect 3497 4870 3507 4922
rect 3531 4870 3561 4922
rect 3561 4870 3573 4922
rect 3573 4870 3587 4922
rect 3611 4870 3625 4922
rect 3625 4870 3637 4922
rect 3637 4870 3667 4922
rect 3691 4870 3701 4922
rect 3701 4870 3747 4922
rect 3451 4868 3507 4870
rect 3531 4868 3587 4870
rect 3611 4868 3667 4870
rect 3691 4868 3747 4870
rect 3606 4120 3662 4176
rect 3451 3834 3507 3836
rect 3531 3834 3587 3836
rect 3611 3834 3667 3836
rect 3691 3834 3747 3836
rect 3451 3782 3497 3834
rect 3497 3782 3507 3834
rect 3531 3782 3561 3834
rect 3561 3782 3573 3834
rect 3573 3782 3587 3834
rect 3611 3782 3625 3834
rect 3625 3782 3637 3834
rect 3637 3782 3667 3834
rect 3691 3782 3701 3834
rect 3701 3782 3747 3834
rect 3451 3780 3507 3782
rect 3531 3780 3587 3782
rect 3611 3780 3667 3782
rect 3691 3780 3747 3782
rect 3882 4664 3938 4720
rect 3451 2746 3507 2748
rect 3531 2746 3587 2748
rect 3611 2746 3667 2748
rect 3691 2746 3747 2748
rect 3451 2694 3497 2746
rect 3497 2694 3507 2746
rect 3531 2694 3561 2746
rect 3561 2694 3573 2746
rect 3573 2694 3587 2746
rect 3611 2694 3625 2746
rect 3625 2694 3637 2746
rect 3637 2694 3667 2746
rect 3691 2694 3701 2746
rect 3701 2694 3747 2746
rect 3451 2692 3507 2694
rect 3531 2692 3587 2694
rect 3611 2692 3667 2694
rect 3691 2692 3747 2694
rect 3330 2352 3386 2408
rect 3238 1808 3294 1864
rect 3451 1658 3507 1660
rect 3531 1658 3587 1660
rect 3611 1658 3667 1660
rect 3691 1658 3747 1660
rect 3451 1606 3497 1658
rect 3497 1606 3507 1658
rect 3531 1606 3561 1658
rect 3561 1606 3573 1658
rect 3573 1606 3587 1658
rect 3611 1606 3625 1658
rect 3625 1606 3637 1658
rect 3637 1606 3667 1658
rect 3691 1606 3701 1658
rect 3701 1606 3747 1658
rect 3451 1604 3507 1606
rect 3531 1604 3587 1606
rect 3611 1604 3667 1606
rect 3691 1604 3747 1606
rect 4802 6704 4858 6760
rect 4313 6554 4369 6556
rect 4393 6554 4449 6556
rect 4473 6554 4529 6556
rect 4553 6554 4609 6556
rect 4313 6502 4359 6554
rect 4359 6502 4369 6554
rect 4393 6502 4423 6554
rect 4423 6502 4435 6554
rect 4435 6502 4449 6554
rect 4473 6502 4487 6554
rect 4487 6502 4499 6554
rect 4499 6502 4529 6554
rect 4553 6502 4563 6554
rect 4563 6502 4609 6554
rect 4313 6500 4369 6502
rect 4393 6500 4449 6502
rect 4473 6500 4529 6502
rect 4553 6500 4609 6502
rect 4313 5466 4369 5468
rect 4393 5466 4449 5468
rect 4473 5466 4529 5468
rect 4553 5466 4609 5468
rect 4313 5414 4359 5466
rect 4359 5414 4369 5466
rect 4393 5414 4423 5466
rect 4423 5414 4435 5466
rect 4435 5414 4449 5466
rect 4473 5414 4487 5466
rect 4487 5414 4499 5466
rect 4499 5414 4529 5466
rect 4553 5414 4563 5466
rect 4563 5414 4609 5466
rect 4313 5412 4369 5414
rect 4393 5412 4449 5414
rect 4473 5412 4529 5414
rect 4553 5412 4609 5414
rect 4313 4378 4369 4380
rect 4393 4378 4449 4380
rect 4473 4378 4529 4380
rect 4553 4378 4609 4380
rect 4313 4326 4359 4378
rect 4359 4326 4369 4378
rect 4393 4326 4423 4378
rect 4423 4326 4435 4378
rect 4435 4326 4449 4378
rect 4473 4326 4487 4378
rect 4487 4326 4499 4378
rect 4499 4326 4529 4378
rect 4553 4326 4563 4378
rect 4563 4326 4609 4378
rect 4313 4324 4369 4326
rect 4393 4324 4449 4326
rect 4473 4324 4529 4326
rect 4553 4324 4609 4326
rect 4066 3576 4122 3632
rect 4710 3576 4766 3632
rect 4313 3290 4369 3292
rect 4393 3290 4449 3292
rect 4473 3290 4529 3292
rect 4553 3290 4609 3292
rect 4313 3238 4359 3290
rect 4359 3238 4369 3290
rect 4393 3238 4423 3290
rect 4423 3238 4435 3290
rect 4435 3238 4449 3290
rect 4473 3238 4487 3290
rect 4487 3238 4499 3290
rect 4499 3238 4529 3290
rect 4553 3238 4563 3290
rect 4563 3238 4609 3290
rect 4313 3236 4369 3238
rect 4393 3236 4449 3238
rect 4473 3236 4529 3238
rect 4553 3236 4609 3238
rect 4710 3032 4766 3088
rect 4313 2202 4369 2204
rect 4393 2202 4449 2204
rect 4473 2202 4529 2204
rect 4553 2202 4609 2204
rect 4313 2150 4359 2202
rect 4359 2150 4369 2202
rect 4393 2150 4423 2202
rect 4423 2150 4435 2202
rect 4435 2150 4449 2202
rect 4473 2150 4487 2202
rect 4487 2150 4499 2202
rect 4499 2150 4529 2202
rect 4553 2150 4563 2202
rect 4563 2150 4609 2202
rect 4313 2148 4369 2150
rect 4393 2148 4449 2150
rect 4473 2148 4529 2150
rect 4553 2148 4609 2150
rect 5176 8186 5232 8188
rect 5256 8186 5312 8188
rect 5336 8186 5392 8188
rect 5416 8186 5472 8188
rect 5176 8134 5222 8186
rect 5222 8134 5232 8186
rect 5256 8134 5286 8186
rect 5286 8134 5298 8186
rect 5298 8134 5312 8186
rect 5336 8134 5350 8186
rect 5350 8134 5362 8186
rect 5362 8134 5392 8186
rect 5416 8134 5426 8186
rect 5426 8134 5472 8186
rect 5176 8132 5232 8134
rect 5256 8132 5312 8134
rect 5336 8132 5392 8134
rect 5416 8132 5472 8134
rect 5354 7928 5410 7984
rect 5176 7098 5232 7100
rect 5256 7098 5312 7100
rect 5336 7098 5392 7100
rect 5416 7098 5472 7100
rect 5176 7046 5222 7098
rect 5222 7046 5232 7098
rect 5256 7046 5286 7098
rect 5286 7046 5298 7098
rect 5298 7046 5312 7098
rect 5336 7046 5350 7098
rect 5350 7046 5362 7098
rect 5362 7046 5392 7098
rect 5416 7046 5426 7098
rect 5426 7046 5472 7098
rect 5176 7044 5232 7046
rect 5256 7044 5312 7046
rect 5336 7044 5392 7046
rect 5416 7044 5472 7046
rect 5176 6010 5232 6012
rect 5256 6010 5312 6012
rect 5336 6010 5392 6012
rect 5416 6010 5472 6012
rect 5176 5958 5222 6010
rect 5222 5958 5232 6010
rect 5256 5958 5286 6010
rect 5286 5958 5298 6010
rect 5298 5958 5312 6010
rect 5336 5958 5350 6010
rect 5350 5958 5362 6010
rect 5362 5958 5392 6010
rect 5416 5958 5426 6010
rect 5426 5958 5472 6010
rect 5176 5956 5232 5958
rect 5256 5956 5312 5958
rect 5336 5956 5392 5958
rect 5416 5956 5472 5958
rect 5446 5772 5502 5808
rect 5446 5752 5448 5772
rect 5448 5752 5500 5772
rect 5500 5752 5502 5772
rect 5538 5072 5594 5128
rect 5176 4922 5232 4924
rect 5256 4922 5312 4924
rect 5336 4922 5392 4924
rect 5416 4922 5472 4924
rect 5176 4870 5222 4922
rect 5222 4870 5232 4922
rect 5256 4870 5286 4922
rect 5286 4870 5298 4922
rect 5298 4870 5312 4922
rect 5336 4870 5350 4922
rect 5350 4870 5362 4922
rect 5362 4870 5392 4922
rect 5416 4870 5426 4922
rect 5426 4870 5472 4922
rect 5176 4868 5232 4870
rect 5256 4868 5312 4870
rect 5336 4868 5392 4870
rect 5416 4868 5472 4870
rect 5176 3834 5232 3836
rect 5256 3834 5312 3836
rect 5336 3834 5392 3836
rect 5416 3834 5472 3836
rect 5176 3782 5222 3834
rect 5222 3782 5232 3834
rect 5256 3782 5286 3834
rect 5286 3782 5298 3834
rect 5298 3782 5312 3834
rect 5336 3782 5350 3834
rect 5350 3782 5362 3834
rect 5362 3782 5392 3834
rect 5416 3782 5426 3834
rect 5426 3782 5472 3834
rect 5176 3780 5232 3782
rect 5256 3780 5312 3782
rect 5336 3780 5392 3782
rect 5416 3780 5472 3782
rect 4313 1114 4369 1116
rect 4393 1114 4449 1116
rect 4473 1114 4529 1116
rect 4553 1114 4609 1116
rect 4313 1062 4359 1114
rect 4359 1062 4369 1114
rect 4393 1062 4423 1114
rect 4423 1062 4435 1114
rect 4435 1062 4449 1114
rect 4473 1062 4487 1114
rect 4487 1062 4499 1114
rect 4499 1062 4529 1114
rect 4553 1062 4563 1114
rect 4563 1062 4609 1114
rect 4313 1060 4369 1062
rect 4393 1060 4449 1062
rect 4473 1060 4529 1062
rect 4553 1060 4609 1062
rect 5176 2746 5232 2748
rect 5256 2746 5312 2748
rect 5336 2746 5392 2748
rect 5416 2746 5472 2748
rect 5176 2694 5222 2746
rect 5222 2694 5232 2746
rect 5256 2694 5286 2746
rect 5286 2694 5298 2746
rect 5298 2694 5312 2746
rect 5336 2694 5350 2746
rect 5350 2694 5362 2746
rect 5362 2694 5392 2746
rect 5416 2694 5426 2746
rect 5426 2694 5472 2746
rect 5176 2692 5232 2694
rect 5256 2692 5312 2694
rect 5336 2692 5392 2694
rect 5416 2692 5472 2694
rect 6038 8730 6094 8732
rect 6118 8730 6174 8732
rect 6198 8730 6254 8732
rect 6278 8730 6334 8732
rect 6038 8678 6084 8730
rect 6084 8678 6094 8730
rect 6118 8678 6148 8730
rect 6148 8678 6160 8730
rect 6160 8678 6174 8730
rect 6198 8678 6212 8730
rect 6212 8678 6224 8730
rect 6224 8678 6254 8730
rect 6278 8678 6288 8730
rect 6288 8678 6334 8730
rect 6038 8676 6094 8678
rect 6118 8676 6174 8678
rect 6198 8676 6254 8678
rect 6278 8676 6334 8678
rect 6038 7642 6094 7644
rect 6118 7642 6174 7644
rect 6198 7642 6254 7644
rect 6278 7642 6334 7644
rect 6038 7590 6084 7642
rect 6084 7590 6094 7642
rect 6118 7590 6148 7642
rect 6148 7590 6160 7642
rect 6160 7590 6174 7642
rect 6198 7590 6212 7642
rect 6212 7590 6224 7642
rect 6224 7590 6254 7642
rect 6278 7590 6288 7642
rect 6288 7590 6334 7642
rect 6038 7588 6094 7590
rect 6118 7588 6174 7590
rect 6198 7588 6254 7590
rect 6278 7588 6334 7590
rect 6038 6554 6094 6556
rect 6118 6554 6174 6556
rect 6198 6554 6254 6556
rect 6278 6554 6334 6556
rect 6038 6502 6084 6554
rect 6084 6502 6094 6554
rect 6118 6502 6148 6554
rect 6148 6502 6160 6554
rect 6160 6502 6174 6554
rect 6198 6502 6212 6554
rect 6212 6502 6224 6554
rect 6224 6502 6254 6554
rect 6278 6502 6288 6554
rect 6288 6502 6334 6554
rect 6038 6500 6094 6502
rect 6118 6500 6174 6502
rect 6198 6500 6254 6502
rect 6278 6500 6334 6502
rect 5906 6296 5962 6352
rect 6366 6160 6422 6216
rect 6550 8336 6606 8392
rect 6038 5466 6094 5468
rect 6118 5466 6174 5468
rect 6198 5466 6254 5468
rect 6278 5466 6334 5468
rect 6038 5414 6084 5466
rect 6084 5414 6094 5466
rect 6118 5414 6148 5466
rect 6148 5414 6160 5466
rect 6160 5414 6174 5466
rect 6198 5414 6212 5466
rect 6212 5414 6224 5466
rect 6224 5414 6254 5466
rect 6278 5414 6288 5466
rect 6288 5414 6334 5466
rect 6038 5412 6094 5414
rect 6118 5412 6174 5414
rect 6198 5412 6254 5414
rect 6278 5412 6334 5414
rect 6038 4378 6094 4380
rect 6118 4378 6174 4380
rect 6198 4378 6254 4380
rect 6278 4378 6334 4380
rect 6038 4326 6084 4378
rect 6084 4326 6094 4378
rect 6118 4326 6148 4378
rect 6148 4326 6160 4378
rect 6160 4326 6174 4378
rect 6198 4326 6212 4378
rect 6212 4326 6224 4378
rect 6224 4326 6254 4378
rect 6278 4326 6288 4378
rect 6288 4326 6334 4378
rect 6038 4324 6094 4326
rect 6118 4324 6174 4326
rect 6198 4324 6254 4326
rect 6278 4324 6334 4326
rect 5176 1658 5232 1660
rect 5256 1658 5312 1660
rect 5336 1658 5392 1660
rect 5416 1658 5472 1660
rect 5176 1606 5222 1658
rect 5222 1606 5232 1658
rect 5256 1606 5286 1658
rect 5286 1606 5298 1658
rect 5298 1606 5312 1658
rect 5336 1606 5350 1658
rect 5350 1606 5362 1658
rect 5362 1606 5392 1658
rect 5416 1606 5426 1658
rect 5426 1606 5472 1658
rect 5176 1604 5232 1606
rect 5256 1604 5312 1606
rect 5336 1604 5392 1606
rect 5416 1604 5472 1606
rect 6038 3290 6094 3292
rect 6118 3290 6174 3292
rect 6198 3290 6254 3292
rect 6278 3290 6334 3292
rect 6038 3238 6084 3290
rect 6084 3238 6094 3290
rect 6118 3238 6148 3290
rect 6148 3238 6160 3290
rect 6160 3238 6174 3290
rect 6198 3238 6212 3290
rect 6212 3238 6224 3290
rect 6224 3238 6254 3290
rect 6278 3238 6288 3290
rect 6288 3238 6334 3290
rect 6038 3236 6094 3238
rect 6118 3236 6174 3238
rect 6198 3236 6254 3238
rect 6278 3236 6334 3238
rect 6366 2488 6422 2544
rect 6901 8186 6957 8188
rect 6981 8186 7037 8188
rect 7061 8186 7117 8188
rect 7141 8186 7197 8188
rect 6901 8134 6947 8186
rect 6947 8134 6957 8186
rect 6981 8134 7011 8186
rect 7011 8134 7023 8186
rect 7023 8134 7037 8186
rect 7061 8134 7075 8186
rect 7075 8134 7087 8186
rect 7087 8134 7117 8186
rect 7141 8134 7151 8186
rect 7151 8134 7197 8186
rect 6901 8132 6957 8134
rect 6981 8132 7037 8134
rect 7061 8132 7117 8134
rect 7141 8132 7197 8134
rect 6901 7098 6957 7100
rect 6981 7098 7037 7100
rect 7061 7098 7117 7100
rect 7141 7098 7197 7100
rect 6901 7046 6947 7098
rect 6947 7046 6957 7098
rect 6981 7046 7011 7098
rect 7011 7046 7023 7098
rect 7023 7046 7037 7098
rect 7061 7046 7075 7098
rect 7075 7046 7087 7098
rect 7087 7046 7117 7098
rect 7141 7046 7151 7098
rect 7151 7046 7197 7098
rect 6901 7044 6957 7046
rect 6981 7044 7037 7046
rect 7061 7044 7117 7046
rect 7141 7044 7197 7046
rect 6550 4120 6606 4176
rect 6038 2202 6094 2204
rect 6118 2202 6174 2204
rect 6198 2202 6254 2204
rect 6278 2202 6334 2204
rect 6038 2150 6084 2202
rect 6084 2150 6094 2202
rect 6118 2150 6148 2202
rect 6148 2150 6160 2202
rect 6160 2150 6174 2202
rect 6198 2150 6212 2202
rect 6212 2150 6224 2202
rect 6224 2150 6254 2202
rect 6278 2150 6288 2202
rect 6288 2150 6334 2202
rect 6038 2148 6094 2150
rect 6118 2148 6174 2150
rect 6198 2148 6254 2150
rect 6278 2148 6334 2150
rect 5906 1400 5962 1456
rect 6038 1114 6094 1116
rect 6118 1114 6174 1116
rect 6198 1114 6254 1116
rect 6278 1114 6334 1116
rect 6038 1062 6084 1114
rect 6084 1062 6094 1114
rect 6118 1062 6148 1114
rect 6148 1062 6160 1114
rect 6160 1062 6174 1114
rect 6198 1062 6212 1114
rect 6212 1062 6224 1114
rect 6224 1062 6254 1114
rect 6278 1062 6288 1114
rect 6288 1062 6334 1114
rect 6038 1060 6094 1062
rect 6118 1060 6174 1062
rect 6198 1060 6254 1062
rect 6278 1060 6334 1062
rect 6458 2352 6514 2408
rect 6901 6010 6957 6012
rect 6981 6010 7037 6012
rect 7061 6010 7117 6012
rect 7141 6010 7197 6012
rect 6901 5958 6947 6010
rect 6947 5958 6957 6010
rect 6981 5958 7011 6010
rect 7011 5958 7023 6010
rect 7023 5958 7037 6010
rect 7061 5958 7075 6010
rect 7075 5958 7087 6010
rect 7087 5958 7117 6010
rect 7141 5958 7151 6010
rect 7151 5958 7197 6010
rect 6901 5956 6957 5958
rect 6981 5956 7037 5958
rect 7061 5956 7117 5958
rect 7141 5956 7197 5958
rect 6901 4922 6957 4924
rect 6981 4922 7037 4924
rect 7061 4922 7117 4924
rect 7141 4922 7197 4924
rect 6901 4870 6947 4922
rect 6947 4870 6957 4922
rect 6981 4870 7011 4922
rect 7011 4870 7023 4922
rect 7023 4870 7037 4922
rect 7061 4870 7075 4922
rect 7075 4870 7087 4922
rect 7087 4870 7117 4922
rect 7141 4870 7151 4922
rect 7151 4870 7197 4922
rect 6901 4868 6957 4870
rect 6981 4868 7037 4870
rect 7061 4868 7117 4870
rect 7141 4868 7197 4870
rect 7470 8880 7526 8936
rect 7286 4664 7342 4720
rect 6734 3984 6790 4040
rect 6901 3834 6957 3836
rect 6981 3834 7037 3836
rect 7061 3834 7117 3836
rect 7141 3834 7197 3836
rect 6901 3782 6947 3834
rect 6947 3782 6957 3834
rect 6981 3782 7011 3834
rect 7011 3782 7023 3834
rect 7023 3782 7037 3834
rect 7061 3782 7075 3834
rect 7075 3782 7087 3834
rect 7087 3782 7117 3834
rect 7141 3782 7151 3834
rect 7151 3782 7197 3834
rect 6901 3780 6957 3782
rect 6981 3780 7037 3782
rect 7061 3780 7117 3782
rect 7141 3780 7197 3782
rect 7763 8730 7819 8732
rect 7843 8730 7899 8732
rect 7923 8730 7979 8732
rect 8003 8730 8059 8732
rect 7763 8678 7809 8730
rect 7809 8678 7819 8730
rect 7843 8678 7873 8730
rect 7873 8678 7885 8730
rect 7885 8678 7899 8730
rect 7923 8678 7937 8730
rect 7937 8678 7949 8730
rect 7949 8678 7979 8730
rect 8003 8678 8013 8730
rect 8013 8678 8059 8730
rect 7763 8676 7819 8678
rect 7843 8676 7899 8678
rect 7923 8676 7979 8678
rect 8003 8676 8059 8678
rect 7763 7642 7819 7644
rect 7843 7642 7899 7644
rect 7923 7642 7979 7644
rect 8003 7642 8059 7644
rect 7763 7590 7809 7642
rect 7809 7590 7819 7642
rect 7843 7590 7873 7642
rect 7873 7590 7885 7642
rect 7885 7590 7899 7642
rect 7923 7590 7937 7642
rect 7937 7590 7949 7642
rect 7949 7590 7979 7642
rect 8003 7590 8013 7642
rect 8013 7590 8059 7642
rect 7763 7588 7819 7590
rect 7843 7588 7899 7590
rect 7923 7588 7979 7590
rect 8003 7588 8059 7590
rect 7763 6554 7819 6556
rect 7843 6554 7899 6556
rect 7923 6554 7979 6556
rect 8003 6554 8059 6556
rect 7763 6502 7809 6554
rect 7809 6502 7819 6554
rect 7843 6502 7873 6554
rect 7873 6502 7885 6554
rect 7885 6502 7899 6554
rect 7923 6502 7937 6554
rect 7937 6502 7949 6554
rect 7949 6502 7979 6554
rect 8003 6502 8013 6554
rect 8013 6502 8059 6554
rect 7763 6500 7819 6502
rect 7843 6500 7899 6502
rect 7923 6500 7979 6502
rect 8003 6500 8059 6502
rect 8022 5616 8078 5672
rect 7763 5466 7819 5468
rect 7843 5466 7899 5468
rect 7923 5466 7979 5468
rect 8003 5466 8059 5468
rect 7763 5414 7809 5466
rect 7809 5414 7819 5466
rect 7843 5414 7873 5466
rect 7873 5414 7885 5466
rect 7885 5414 7899 5466
rect 7923 5414 7937 5466
rect 7937 5414 7949 5466
rect 7949 5414 7979 5466
rect 8003 5414 8013 5466
rect 8013 5414 8059 5466
rect 7763 5412 7819 5414
rect 7843 5412 7899 5414
rect 7923 5412 7979 5414
rect 8003 5412 8059 5414
rect 7763 4378 7819 4380
rect 7843 4378 7899 4380
rect 7923 4378 7979 4380
rect 8003 4378 8059 4380
rect 7763 4326 7809 4378
rect 7809 4326 7819 4378
rect 7843 4326 7873 4378
rect 7873 4326 7885 4378
rect 7885 4326 7899 4378
rect 7923 4326 7937 4378
rect 7937 4326 7949 4378
rect 7949 4326 7979 4378
rect 8003 4326 8013 4378
rect 8013 4326 8059 4378
rect 7763 4324 7819 4326
rect 7843 4324 7899 4326
rect 7923 4324 7979 4326
rect 8003 4324 8059 4326
rect 7763 3290 7819 3292
rect 7843 3290 7899 3292
rect 7923 3290 7979 3292
rect 8003 3290 8059 3292
rect 7763 3238 7809 3290
rect 7809 3238 7819 3290
rect 7843 3238 7873 3290
rect 7873 3238 7885 3290
rect 7885 3238 7899 3290
rect 7923 3238 7937 3290
rect 7937 3238 7949 3290
rect 7949 3238 7979 3290
rect 8003 3238 8013 3290
rect 8013 3238 8059 3290
rect 7763 3236 7819 3238
rect 7843 3236 7899 3238
rect 7923 3236 7979 3238
rect 8003 3236 8059 3238
rect 6642 3032 6698 3088
rect 6550 1808 6606 1864
rect 6901 2746 6957 2748
rect 6981 2746 7037 2748
rect 7061 2746 7117 2748
rect 7141 2746 7197 2748
rect 6901 2694 6947 2746
rect 6947 2694 6957 2746
rect 6981 2694 7011 2746
rect 7011 2694 7023 2746
rect 7023 2694 7037 2746
rect 7061 2694 7075 2746
rect 7075 2694 7087 2746
rect 7087 2694 7117 2746
rect 7141 2694 7151 2746
rect 7151 2694 7197 2746
rect 6901 2692 6957 2694
rect 6981 2692 7037 2694
rect 7061 2692 7117 2694
rect 7141 2692 7197 2694
rect 6901 1658 6957 1660
rect 6981 1658 7037 1660
rect 7061 1658 7117 1660
rect 7141 1658 7197 1660
rect 6901 1606 6947 1658
rect 6947 1606 6957 1658
rect 6981 1606 7011 1658
rect 7011 1606 7023 1658
rect 7023 1606 7037 1658
rect 7061 1606 7075 1658
rect 7075 1606 7087 1658
rect 7087 1606 7117 1658
rect 7141 1606 7151 1658
rect 7151 1606 7197 1658
rect 6901 1604 6957 1606
rect 6981 1604 7037 1606
rect 7061 1604 7117 1606
rect 7141 1604 7197 1606
rect 7763 2202 7819 2204
rect 7843 2202 7899 2204
rect 7923 2202 7979 2204
rect 8003 2202 8059 2204
rect 7763 2150 7809 2202
rect 7809 2150 7819 2202
rect 7843 2150 7873 2202
rect 7873 2150 7885 2202
rect 7885 2150 7899 2202
rect 7923 2150 7937 2202
rect 7937 2150 7949 2202
rect 7949 2150 7979 2202
rect 8003 2150 8013 2202
rect 8013 2150 8059 2202
rect 7763 2148 7819 2150
rect 7843 2148 7899 2150
rect 7923 2148 7979 2150
rect 8003 2148 8059 2150
rect 7378 856 7434 912
rect 7763 1114 7819 1116
rect 7843 1114 7899 1116
rect 7923 1114 7979 1116
rect 8003 1114 8059 1116
rect 7763 1062 7809 1114
rect 7809 1062 7819 1114
rect 7843 1062 7873 1114
rect 7873 1062 7885 1114
rect 7885 1062 7899 1114
rect 7923 1062 7937 1114
rect 7937 1062 7949 1114
rect 7949 1062 7979 1114
rect 8003 1062 8013 1114
rect 8013 1062 8059 1114
rect 7763 1060 7819 1062
rect 7843 1060 7899 1062
rect 7923 1060 7979 1062
rect 8003 1060 8059 1062
rect 6826 584 6882 640
<< metal3 >>
rect 5574 9148 5580 9212
rect 5644 9210 5650 9212
rect 8200 9210 9000 9240
rect 5644 9150 9000 9210
rect 5644 9148 5650 9150
rect 8200 9120 9000 9150
rect 0 9074 800 9104
rect 3325 9074 3391 9077
rect 0 9072 3391 9074
rect 0 9016 3330 9072
rect 3386 9016 3391 9072
rect 0 9014 3391 9016
rect 0 8984 800 9014
rect 3325 9011 3391 9014
rect 7465 8938 7531 8941
rect 7465 8936 8218 8938
rect 7465 8880 7470 8936
rect 7526 8880 8218 8936
rect 7465 8878 8218 8880
rect 7465 8875 7531 8878
rect 8158 8832 8218 8878
rect 8158 8742 9000 8832
rect 2578 8736 2894 8737
rect 2578 8672 2584 8736
rect 2648 8672 2664 8736
rect 2728 8672 2744 8736
rect 2808 8672 2824 8736
rect 2888 8672 2894 8736
rect 2578 8671 2894 8672
rect 4303 8736 4619 8737
rect 4303 8672 4309 8736
rect 4373 8672 4389 8736
rect 4453 8672 4469 8736
rect 4533 8672 4549 8736
rect 4613 8672 4619 8736
rect 4303 8671 4619 8672
rect 6028 8736 6344 8737
rect 6028 8672 6034 8736
rect 6098 8672 6114 8736
rect 6178 8672 6194 8736
rect 6258 8672 6274 8736
rect 6338 8672 6344 8736
rect 6028 8671 6344 8672
rect 7753 8736 8069 8737
rect 7753 8672 7759 8736
rect 7823 8672 7839 8736
rect 7903 8672 7919 8736
rect 7983 8672 7999 8736
rect 8063 8672 8069 8736
rect 8200 8712 9000 8742
rect 7753 8671 8069 8672
rect 0 8394 800 8424
rect 2405 8394 2471 8397
rect 0 8392 2471 8394
rect 0 8336 2410 8392
rect 2466 8336 2471 8392
rect 0 8334 2471 8336
rect 0 8304 800 8334
rect 2405 8331 2471 8334
rect 6545 8394 6611 8397
rect 8200 8394 9000 8424
rect 6545 8392 9000 8394
rect 6545 8336 6550 8392
rect 6606 8336 9000 8392
rect 6545 8334 9000 8336
rect 6545 8331 6611 8334
rect 8200 8304 9000 8334
rect 1716 8192 2032 8193
rect 1716 8128 1722 8192
rect 1786 8128 1802 8192
rect 1866 8128 1882 8192
rect 1946 8128 1962 8192
rect 2026 8128 2032 8192
rect 1716 8127 2032 8128
rect 3441 8192 3757 8193
rect 3441 8128 3447 8192
rect 3511 8128 3527 8192
rect 3591 8128 3607 8192
rect 3671 8128 3687 8192
rect 3751 8128 3757 8192
rect 3441 8127 3757 8128
rect 5166 8192 5482 8193
rect 5166 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5482 8192
rect 5166 8127 5482 8128
rect 6891 8192 7207 8193
rect 6891 8128 6897 8192
rect 6961 8128 6977 8192
rect 7041 8128 7057 8192
rect 7121 8128 7137 8192
rect 7201 8128 7207 8192
rect 6891 8127 7207 8128
rect 5349 7986 5415 7989
rect 8200 7986 9000 8016
rect 5349 7984 9000 7986
rect 5349 7928 5354 7984
rect 5410 7928 9000 7984
rect 5349 7926 9000 7928
rect 5349 7923 5415 7926
rect 8200 7896 9000 7926
rect 4245 7850 4311 7853
rect 4245 7848 4906 7850
rect 4245 7792 4250 7848
rect 4306 7792 4906 7848
rect 4245 7790 4906 7792
rect 4245 7787 4311 7790
rect 0 7714 800 7744
rect 1209 7714 1275 7717
rect 0 7712 1275 7714
rect 0 7656 1214 7712
rect 1270 7656 1275 7712
rect 0 7654 1275 7656
rect 0 7624 800 7654
rect 1209 7651 1275 7654
rect 2578 7648 2894 7649
rect 2578 7584 2584 7648
rect 2648 7584 2664 7648
rect 2728 7584 2744 7648
rect 2808 7584 2824 7648
rect 2888 7584 2894 7648
rect 2578 7583 2894 7584
rect 4303 7648 4619 7649
rect 4303 7584 4309 7648
rect 4373 7584 4389 7648
rect 4453 7584 4469 7648
rect 4533 7584 4549 7648
rect 4613 7584 4619 7648
rect 4303 7583 4619 7584
rect 4846 7442 4906 7790
rect 6028 7648 6344 7649
rect 6028 7584 6034 7648
rect 6098 7584 6114 7648
rect 6178 7584 6194 7648
rect 6258 7584 6274 7648
rect 6338 7584 6344 7648
rect 6028 7583 6344 7584
rect 7753 7648 8069 7649
rect 7753 7584 7759 7648
rect 7823 7584 7839 7648
rect 7903 7584 7919 7648
rect 7983 7584 7999 7648
rect 8063 7584 8069 7648
rect 7753 7583 8069 7584
rect 8200 7578 9000 7608
rect 8158 7488 9000 7578
rect 8158 7442 8218 7488
rect 4846 7382 8218 7442
rect 4153 7306 4219 7309
rect 4153 7304 7482 7306
rect 4153 7248 4158 7304
rect 4214 7248 7482 7304
rect 4153 7246 7482 7248
rect 4153 7243 4219 7246
rect 7422 7170 7482 7246
rect 8200 7170 9000 7200
rect 7422 7110 9000 7170
rect 1716 7104 2032 7105
rect 0 7034 800 7064
rect 1716 7040 1722 7104
rect 1786 7040 1802 7104
rect 1866 7040 1882 7104
rect 1946 7040 1962 7104
rect 2026 7040 2032 7104
rect 1716 7039 2032 7040
rect 3441 7104 3757 7105
rect 3441 7040 3447 7104
rect 3511 7040 3527 7104
rect 3591 7040 3607 7104
rect 3671 7040 3687 7104
rect 3751 7040 3757 7104
rect 3441 7039 3757 7040
rect 5166 7104 5482 7105
rect 5166 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5482 7104
rect 5166 7039 5482 7040
rect 6891 7104 7207 7105
rect 6891 7040 6897 7104
rect 6961 7040 6977 7104
rect 7041 7040 7057 7104
rect 7121 7040 7137 7104
rect 7201 7040 7207 7104
rect 8200 7080 9000 7110
rect 6891 7039 7207 7040
rect 1577 7034 1643 7037
rect 0 7032 1643 7034
rect 0 6976 1582 7032
rect 1638 6976 1643 7032
rect 0 6974 1643 6976
rect 0 6944 800 6974
rect 1577 6971 1643 6974
rect 4797 6762 4863 6765
rect 8200 6762 9000 6792
rect 4797 6760 9000 6762
rect 4797 6704 4802 6760
rect 4858 6704 9000 6760
rect 4797 6702 9000 6704
rect 4797 6699 4863 6702
rect 8200 6672 9000 6702
rect 2578 6560 2894 6561
rect 2578 6496 2584 6560
rect 2648 6496 2664 6560
rect 2728 6496 2744 6560
rect 2808 6496 2824 6560
rect 2888 6496 2894 6560
rect 2578 6495 2894 6496
rect 4303 6560 4619 6561
rect 4303 6496 4309 6560
rect 4373 6496 4389 6560
rect 4453 6496 4469 6560
rect 4533 6496 4549 6560
rect 4613 6496 4619 6560
rect 4303 6495 4619 6496
rect 6028 6560 6344 6561
rect 6028 6496 6034 6560
rect 6098 6496 6114 6560
rect 6178 6496 6194 6560
rect 6258 6496 6274 6560
rect 6338 6496 6344 6560
rect 6028 6495 6344 6496
rect 7753 6560 8069 6561
rect 7753 6496 7759 6560
rect 7823 6496 7839 6560
rect 7903 6496 7919 6560
rect 7983 6496 7999 6560
rect 8063 6496 8069 6560
rect 7753 6495 8069 6496
rect 0 6354 800 6384
rect 4102 6354 4108 6356
rect 0 6294 4108 6354
rect 0 6264 800 6294
rect 4102 6292 4108 6294
rect 4172 6292 4178 6356
rect 5901 6354 5967 6357
rect 8200 6354 9000 6384
rect 5901 6352 9000 6354
rect 5901 6296 5906 6352
rect 5962 6296 9000 6352
rect 5901 6294 9000 6296
rect 5901 6291 5967 6294
rect 8200 6264 9000 6294
rect 6361 6218 6427 6221
rect 6361 6216 7482 6218
rect 6361 6160 6366 6216
rect 6422 6160 7482 6216
rect 6361 6158 7482 6160
rect 6361 6155 6427 6158
rect 1716 6016 2032 6017
rect 1716 5952 1722 6016
rect 1786 5952 1802 6016
rect 1866 5952 1882 6016
rect 1946 5952 1962 6016
rect 2026 5952 2032 6016
rect 1716 5951 2032 5952
rect 3441 6016 3757 6017
rect 3441 5952 3447 6016
rect 3511 5952 3527 6016
rect 3591 5952 3607 6016
rect 3671 5952 3687 6016
rect 3751 5952 3757 6016
rect 3441 5951 3757 5952
rect 5166 6016 5482 6017
rect 5166 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5482 6016
rect 5166 5951 5482 5952
rect 6891 6016 7207 6017
rect 6891 5952 6897 6016
rect 6961 5952 6977 6016
rect 7041 5952 7057 6016
rect 7121 5952 7137 6016
rect 7201 5952 7207 6016
rect 6891 5951 7207 5952
rect 7422 5946 7482 6158
rect 8200 5946 9000 5976
rect 7422 5886 9000 5946
rect 8200 5856 9000 5886
rect 5441 5810 5507 5813
rect 5574 5810 5580 5812
rect 5441 5808 5580 5810
rect 5441 5752 5446 5808
rect 5502 5752 5580 5808
rect 5441 5750 5580 5752
rect 5441 5747 5507 5750
rect 5574 5748 5580 5750
rect 5644 5748 5650 5812
rect 0 5674 800 5704
rect 3233 5674 3299 5677
rect 0 5672 3299 5674
rect 0 5616 3238 5672
rect 3294 5616 3299 5672
rect 0 5614 3299 5616
rect 0 5584 800 5614
rect 3233 5611 3299 5614
rect 8017 5674 8083 5677
rect 8017 5672 8218 5674
rect 8017 5616 8022 5672
rect 8078 5616 8218 5672
rect 8017 5614 8218 5616
rect 8017 5611 8083 5614
rect 8158 5568 8218 5614
rect 8158 5478 9000 5568
rect 2578 5472 2894 5473
rect 2578 5408 2584 5472
rect 2648 5408 2664 5472
rect 2728 5408 2744 5472
rect 2808 5408 2824 5472
rect 2888 5408 2894 5472
rect 2578 5407 2894 5408
rect 4303 5472 4619 5473
rect 4303 5408 4309 5472
rect 4373 5408 4389 5472
rect 4453 5408 4469 5472
rect 4533 5408 4549 5472
rect 4613 5408 4619 5472
rect 4303 5407 4619 5408
rect 6028 5472 6344 5473
rect 6028 5408 6034 5472
rect 6098 5408 6114 5472
rect 6178 5408 6194 5472
rect 6258 5408 6274 5472
rect 6338 5408 6344 5472
rect 6028 5407 6344 5408
rect 7753 5472 8069 5473
rect 7753 5408 7759 5472
rect 7823 5408 7839 5472
rect 7903 5408 7919 5472
rect 7983 5408 7999 5472
rect 8063 5408 8069 5472
rect 8200 5448 9000 5478
rect 7753 5407 8069 5408
rect 5533 5130 5599 5133
rect 8200 5130 9000 5160
rect 5533 5128 9000 5130
rect 5533 5072 5538 5128
rect 5594 5072 9000 5128
rect 5533 5070 9000 5072
rect 5533 5067 5599 5070
rect 8200 5040 9000 5070
rect 0 4994 800 5024
rect 0 4934 1640 4994
rect 0 4904 800 4934
rect 1580 4722 1640 4934
rect 1716 4928 2032 4929
rect 1716 4864 1722 4928
rect 1786 4864 1802 4928
rect 1866 4864 1882 4928
rect 1946 4864 1962 4928
rect 2026 4864 2032 4928
rect 1716 4863 2032 4864
rect 3441 4928 3757 4929
rect 3441 4864 3447 4928
rect 3511 4864 3527 4928
rect 3591 4864 3607 4928
rect 3671 4864 3687 4928
rect 3751 4864 3757 4928
rect 3441 4863 3757 4864
rect 5166 4928 5482 4929
rect 5166 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5482 4928
rect 5166 4863 5482 4864
rect 6891 4928 7207 4929
rect 6891 4864 6897 4928
rect 6961 4864 6977 4928
rect 7041 4864 7057 4928
rect 7121 4864 7137 4928
rect 7201 4864 7207 4928
rect 6891 4863 7207 4864
rect 3877 4722 3943 4725
rect 1580 4720 3943 4722
rect 1580 4664 3882 4720
rect 3938 4664 3943 4720
rect 1580 4662 3943 4664
rect 3877 4659 3943 4662
rect 7281 4722 7347 4725
rect 8200 4722 9000 4752
rect 7281 4720 9000 4722
rect 7281 4664 7286 4720
rect 7342 4664 9000 4720
rect 7281 4662 9000 4664
rect 7281 4659 7347 4662
rect 8200 4632 9000 4662
rect 2578 4384 2894 4385
rect 0 4314 800 4344
rect 2578 4320 2584 4384
rect 2648 4320 2664 4384
rect 2728 4320 2744 4384
rect 2808 4320 2824 4384
rect 2888 4320 2894 4384
rect 2578 4319 2894 4320
rect 4303 4384 4619 4385
rect 4303 4320 4309 4384
rect 4373 4320 4389 4384
rect 4453 4320 4469 4384
rect 4533 4320 4549 4384
rect 4613 4320 4619 4384
rect 4303 4319 4619 4320
rect 6028 4384 6344 4385
rect 6028 4320 6034 4384
rect 6098 4320 6114 4384
rect 6178 4320 6194 4384
rect 6258 4320 6274 4384
rect 6338 4320 6344 4384
rect 6028 4319 6344 4320
rect 7753 4384 8069 4385
rect 7753 4320 7759 4384
rect 7823 4320 7839 4384
rect 7903 4320 7919 4384
rect 7983 4320 7999 4384
rect 8063 4320 8069 4384
rect 7753 4319 8069 4320
rect 8200 4314 9000 4344
rect 0 4254 2514 4314
rect 0 4224 800 4254
rect 2454 4178 2514 4254
rect 8158 4224 9000 4314
rect 3601 4178 3667 4181
rect 2454 4176 3667 4178
rect 2454 4120 3606 4176
rect 3662 4120 3667 4176
rect 2454 4118 3667 4120
rect 3601 4115 3667 4118
rect 6545 4178 6611 4181
rect 8158 4178 8218 4224
rect 6545 4176 8218 4178
rect 6545 4120 6550 4176
rect 6606 4120 8218 4176
rect 6545 4118 8218 4120
rect 6545 4115 6611 4118
rect 6729 4042 6795 4045
rect 6729 4040 7482 4042
rect 6729 3984 6734 4040
rect 6790 3984 7482 4040
rect 6729 3982 7482 3984
rect 6729 3979 6795 3982
rect 7422 3906 7482 3982
rect 8200 3906 9000 3936
rect 7422 3846 9000 3906
rect 1716 3840 2032 3841
rect 1716 3776 1722 3840
rect 1786 3776 1802 3840
rect 1866 3776 1882 3840
rect 1946 3776 1962 3840
rect 2026 3776 2032 3840
rect 1716 3775 2032 3776
rect 3441 3840 3757 3841
rect 3441 3776 3447 3840
rect 3511 3776 3527 3840
rect 3591 3776 3607 3840
rect 3671 3776 3687 3840
rect 3751 3776 3757 3840
rect 3441 3775 3757 3776
rect 5166 3840 5482 3841
rect 5166 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5482 3840
rect 5166 3775 5482 3776
rect 6891 3840 7207 3841
rect 6891 3776 6897 3840
rect 6961 3776 6977 3840
rect 7041 3776 7057 3840
rect 7121 3776 7137 3840
rect 7201 3776 7207 3840
rect 8200 3816 9000 3846
rect 6891 3775 7207 3776
rect 0 3634 800 3664
rect 4061 3634 4127 3637
rect 0 3632 4127 3634
rect 0 3576 4066 3632
rect 4122 3576 4127 3632
rect 0 3574 4127 3576
rect 0 3544 800 3574
rect 4061 3571 4127 3574
rect 4705 3634 4771 3637
rect 4705 3632 4906 3634
rect 4705 3576 4710 3632
rect 4766 3576 4906 3632
rect 4705 3574 4906 3576
rect 4705 3571 4771 3574
rect 4846 3498 4906 3574
rect 8200 3498 9000 3528
rect 4846 3438 9000 3498
rect 8200 3408 9000 3438
rect 2578 3296 2894 3297
rect 2578 3232 2584 3296
rect 2648 3232 2664 3296
rect 2728 3232 2744 3296
rect 2808 3232 2824 3296
rect 2888 3232 2894 3296
rect 2578 3231 2894 3232
rect 4303 3296 4619 3297
rect 4303 3232 4309 3296
rect 4373 3232 4389 3296
rect 4453 3232 4469 3296
rect 4533 3232 4549 3296
rect 4613 3232 4619 3296
rect 4303 3231 4619 3232
rect 6028 3296 6344 3297
rect 6028 3232 6034 3296
rect 6098 3232 6114 3296
rect 6178 3232 6194 3296
rect 6258 3232 6274 3296
rect 6338 3232 6344 3296
rect 6028 3231 6344 3232
rect 7753 3296 8069 3297
rect 7753 3232 7759 3296
rect 7823 3232 7839 3296
rect 7903 3232 7919 3296
rect 7983 3232 7999 3296
rect 8063 3232 8069 3296
rect 7753 3231 8069 3232
rect 4102 3028 4108 3092
rect 4172 3090 4178 3092
rect 4705 3090 4771 3093
rect 4172 3088 4771 3090
rect 4172 3032 4710 3088
rect 4766 3032 4771 3088
rect 4172 3030 4771 3032
rect 4172 3028 4178 3030
rect 4705 3027 4771 3030
rect 6637 3090 6703 3093
rect 8200 3090 9000 3120
rect 6637 3088 9000 3090
rect 6637 3032 6642 3088
rect 6698 3032 9000 3088
rect 6637 3030 9000 3032
rect 6637 3027 6703 3030
rect 8200 3000 9000 3030
rect 0 2954 800 2984
rect 2957 2954 3023 2957
rect 0 2952 3023 2954
rect 0 2896 2962 2952
rect 3018 2896 3023 2952
rect 0 2894 3023 2896
rect 0 2864 800 2894
rect 2957 2891 3023 2894
rect 1716 2752 2032 2753
rect 1716 2688 1722 2752
rect 1786 2688 1802 2752
rect 1866 2688 1882 2752
rect 1946 2688 1962 2752
rect 2026 2688 2032 2752
rect 1716 2687 2032 2688
rect 3441 2752 3757 2753
rect 3441 2688 3447 2752
rect 3511 2688 3527 2752
rect 3591 2688 3607 2752
rect 3671 2688 3687 2752
rect 3751 2688 3757 2752
rect 3441 2687 3757 2688
rect 5166 2752 5482 2753
rect 5166 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5482 2752
rect 5166 2687 5482 2688
rect 6891 2752 7207 2753
rect 6891 2688 6897 2752
rect 6961 2688 6977 2752
rect 7041 2688 7057 2752
rect 7121 2688 7137 2752
rect 7201 2688 7207 2752
rect 6891 2687 7207 2688
rect 8200 2682 9000 2712
rect 7422 2622 9000 2682
rect 6361 2546 6427 2549
rect 7422 2546 7482 2622
rect 8200 2592 9000 2622
rect 6361 2544 7482 2546
rect 6361 2488 6366 2544
rect 6422 2488 7482 2544
rect 6361 2486 7482 2488
rect 6361 2483 6427 2486
rect 3325 2410 3391 2413
rect 2454 2408 3391 2410
rect 2454 2352 3330 2408
rect 3386 2352 3391 2408
rect 2454 2350 3391 2352
rect 0 2274 800 2304
rect 2454 2274 2514 2350
rect 3325 2347 3391 2350
rect 6453 2410 6519 2413
rect 6453 2408 8218 2410
rect 6453 2352 6458 2408
rect 6514 2352 8218 2408
rect 6453 2350 8218 2352
rect 6453 2347 6519 2350
rect 0 2214 2514 2274
rect 8158 2304 8218 2350
rect 8158 2214 9000 2304
rect 0 2184 800 2214
rect 2578 2208 2894 2209
rect 2578 2144 2584 2208
rect 2648 2144 2664 2208
rect 2728 2144 2744 2208
rect 2808 2144 2824 2208
rect 2888 2144 2894 2208
rect 2578 2143 2894 2144
rect 4303 2208 4619 2209
rect 4303 2144 4309 2208
rect 4373 2144 4389 2208
rect 4453 2144 4469 2208
rect 4533 2144 4549 2208
rect 4613 2144 4619 2208
rect 4303 2143 4619 2144
rect 6028 2208 6344 2209
rect 6028 2144 6034 2208
rect 6098 2144 6114 2208
rect 6178 2144 6194 2208
rect 6258 2144 6274 2208
rect 6338 2144 6344 2208
rect 6028 2143 6344 2144
rect 7753 2208 8069 2209
rect 7753 2144 7759 2208
rect 7823 2144 7839 2208
rect 7903 2144 7919 2208
rect 7983 2144 7999 2208
rect 8063 2144 8069 2208
rect 8200 2184 9000 2214
rect 7753 2143 8069 2144
rect 3233 1866 3299 1869
rect 1580 1864 3299 1866
rect 1580 1808 3238 1864
rect 3294 1808 3299 1864
rect 1580 1806 3299 1808
rect 0 1594 800 1624
rect 1580 1594 1640 1806
rect 3233 1803 3299 1806
rect 6545 1866 6611 1869
rect 8200 1866 9000 1896
rect 6545 1864 9000 1866
rect 6545 1808 6550 1864
rect 6606 1808 9000 1864
rect 6545 1806 9000 1808
rect 6545 1803 6611 1806
rect 8200 1776 9000 1806
rect 1716 1664 2032 1665
rect 1716 1600 1722 1664
rect 1786 1600 1802 1664
rect 1866 1600 1882 1664
rect 1946 1600 1962 1664
rect 2026 1600 2032 1664
rect 1716 1599 2032 1600
rect 3441 1664 3757 1665
rect 3441 1600 3447 1664
rect 3511 1600 3527 1664
rect 3591 1600 3607 1664
rect 3671 1600 3687 1664
rect 3751 1600 3757 1664
rect 3441 1599 3757 1600
rect 5166 1664 5482 1665
rect 5166 1600 5172 1664
rect 5236 1600 5252 1664
rect 5316 1600 5332 1664
rect 5396 1600 5412 1664
rect 5476 1600 5482 1664
rect 5166 1599 5482 1600
rect 6891 1664 7207 1665
rect 6891 1600 6897 1664
rect 6961 1600 6977 1664
rect 7041 1600 7057 1664
rect 7121 1600 7137 1664
rect 7201 1600 7207 1664
rect 6891 1599 7207 1600
rect 0 1534 1640 1594
rect 0 1504 800 1534
rect 5901 1458 5967 1461
rect 8200 1458 9000 1488
rect 5901 1456 9000 1458
rect 5901 1400 5906 1456
rect 5962 1400 9000 1456
rect 5901 1398 9000 1400
rect 5901 1395 5967 1398
rect 8200 1368 9000 1398
rect 2578 1120 2894 1121
rect 2578 1056 2584 1120
rect 2648 1056 2664 1120
rect 2728 1056 2744 1120
rect 2808 1056 2824 1120
rect 2888 1056 2894 1120
rect 2578 1055 2894 1056
rect 4303 1120 4619 1121
rect 4303 1056 4309 1120
rect 4373 1056 4389 1120
rect 4453 1056 4469 1120
rect 4533 1056 4549 1120
rect 4613 1056 4619 1120
rect 4303 1055 4619 1056
rect 6028 1120 6344 1121
rect 6028 1056 6034 1120
rect 6098 1056 6114 1120
rect 6178 1056 6194 1120
rect 6258 1056 6274 1120
rect 6338 1056 6344 1120
rect 6028 1055 6344 1056
rect 7753 1120 8069 1121
rect 7753 1056 7759 1120
rect 7823 1056 7839 1120
rect 7903 1056 7919 1120
rect 7983 1056 7999 1120
rect 8063 1056 8069 1120
rect 7753 1055 8069 1056
rect 8200 1050 9000 1080
rect 8158 960 9000 1050
rect 0 914 800 944
rect 2497 914 2563 917
rect 0 912 2563 914
rect 0 856 2502 912
rect 2558 856 2563 912
rect 0 854 2563 856
rect 0 824 800 854
rect 2497 851 2563 854
rect 7373 914 7439 917
rect 8158 914 8218 960
rect 7373 912 8218 914
rect 7373 856 7378 912
rect 7434 856 8218 912
rect 7373 854 8218 856
rect 7373 851 7439 854
rect 6821 642 6887 645
rect 8200 642 9000 672
rect 6821 640 9000 642
rect 6821 584 6826 640
rect 6882 584 9000 640
rect 6821 582 9000 584
rect 6821 579 6887 582
rect 8200 552 9000 582
<< via3 >>
rect 5580 9148 5644 9212
rect 2584 8732 2648 8736
rect 2584 8676 2588 8732
rect 2588 8676 2644 8732
rect 2644 8676 2648 8732
rect 2584 8672 2648 8676
rect 2664 8732 2728 8736
rect 2664 8676 2668 8732
rect 2668 8676 2724 8732
rect 2724 8676 2728 8732
rect 2664 8672 2728 8676
rect 2744 8732 2808 8736
rect 2744 8676 2748 8732
rect 2748 8676 2804 8732
rect 2804 8676 2808 8732
rect 2744 8672 2808 8676
rect 2824 8732 2888 8736
rect 2824 8676 2828 8732
rect 2828 8676 2884 8732
rect 2884 8676 2888 8732
rect 2824 8672 2888 8676
rect 4309 8732 4373 8736
rect 4309 8676 4313 8732
rect 4313 8676 4369 8732
rect 4369 8676 4373 8732
rect 4309 8672 4373 8676
rect 4389 8732 4453 8736
rect 4389 8676 4393 8732
rect 4393 8676 4449 8732
rect 4449 8676 4453 8732
rect 4389 8672 4453 8676
rect 4469 8732 4533 8736
rect 4469 8676 4473 8732
rect 4473 8676 4529 8732
rect 4529 8676 4533 8732
rect 4469 8672 4533 8676
rect 4549 8732 4613 8736
rect 4549 8676 4553 8732
rect 4553 8676 4609 8732
rect 4609 8676 4613 8732
rect 4549 8672 4613 8676
rect 6034 8732 6098 8736
rect 6034 8676 6038 8732
rect 6038 8676 6094 8732
rect 6094 8676 6098 8732
rect 6034 8672 6098 8676
rect 6114 8732 6178 8736
rect 6114 8676 6118 8732
rect 6118 8676 6174 8732
rect 6174 8676 6178 8732
rect 6114 8672 6178 8676
rect 6194 8732 6258 8736
rect 6194 8676 6198 8732
rect 6198 8676 6254 8732
rect 6254 8676 6258 8732
rect 6194 8672 6258 8676
rect 6274 8732 6338 8736
rect 6274 8676 6278 8732
rect 6278 8676 6334 8732
rect 6334 8676 6338 8732
rect 6274 8672 6338 8676
rect 7759 8732 7823 8736
rect 7759 8676 7763 8732
rect 7763 8676 7819 8732
rect 7819 8676 7823 8732
rect 7759 8672 7823 8676
rect 7839 8732 7903 8736
rect 7839 8676 7843 8732
rect 7843 8676 7899 8732
rect 7899 8676 7903 8732
rect 7839 8672 7903 8676
rect 7919 8732 7983 8736
rect 7919 8676 7923 8732
rect 7923 8676 7979 8732
rect 7979 8676 7983 8732
rect 7919 8672 7983 8676
rect 7999 8732 8063 8736
rect 7999 8676 8003 8732
rect 8003 8676 8059 8732
rect 8059 8676 8063 8732
rect 7999 8672 8063 8676
rect 1722 8188 1786 8192
rect 1722 8132 1726 8188
rect 1726 8132 1782 8188
rect 1782 8132 1786 8188
rect 1722 8128 1786 8132
rect 1802 8188 1866 8192
rect 1802 8132 1806 8188
rect 1806 8132 1862 8188
rect 1862 8132 1866 8188
rect 1802 8128 1866 8132
rect 1882 8188 1946 8192
rect 1882 8132 1886 8188
rect 1886 8132 1942 8188
rect 1942 8132 1946 8188
rect 1882 8128 1946 8132
rect 1962 8188 2026 8192
rect 1962 8132 1966 8188
rect 1966 8132 2022 8188
rect 2022 8132 2026 8188
rect 1962 8128 2026 8132
rect 3447 8188 3511 8192
rect 3447 8132 3451 8188
rect 3451 8132 3507 8188
rect 3507 8132 3511 8188
rect 3447 8128 3511 8132
rect 3527 8188 3591 8192
rect 3527 8132 3531 8188
rect 3531 8132 3587 8188
rect 3587 8132 3591 8188
rect 3527 8128 3591 8132
rect 3607 8188 3671 8192
rect 3607 8132 3611 8188
rect 3611 8132 3667 8188
rect 3667 8132 3671 8188
rect 3607 8128 3671 8132
rect 3687 8188 3751 8192
rect 3687 8132 3691 8188
rect 3691 8132 3747 8188
rect 3747 8132 3751 8188
rect 3687 8128 3751 8132
rect 5172 8188 5236 8192
rect 5172 8132 5176 8188
rect 5176 8132 5232 8188
rect 5232 8132 5236 8188
rect 5172 8128 5236 8132
rect 5252 8188 5316 8192
rect 5252 8132 5256 8188
rect 5256 8132 5312 8188
rect 5312 8132 5316 8188
rect 5252 8128 5316 8132
rect 5332 8188 5396 8192
rect 5332 8132 5336 8188
rect 5336 8132 5392 8188
rect 5392 8132 5396 8188
rect 5332 8128 5396 8132
rect 5412 8188 5476 8192
rect 5412 8132 5416 8188
rect 5416 8132 5472 8188
rect 5472 8132 5476 8188
rect 5412 8128 5476 8132
rect 6897 8188 6961 8192
rect 6897 8132 6901 8188
rect 6901 8132 6957 8188
rect 6957 8132 6961 8188
rect 6897 8128 6961 8132
rect 6977 8188 7041 8192
rect 6977 8132 6981 8188
rect 6981 8132 7037 8188
rect 7037 8132 7041 8188
rect 6977 8128 7041 8132
rect 7057 8188 7121 8192
rect 7057 8132 7061 8188
rect 7061 8132 7117 8188
rect 7117 8132 7121 8188
rect 7057 8128 7121 8132
rect 7137 8188 7201 8192
rect 7137 8132 7141 8188
rect 7141 8132 7197 8188
rect 7197 8132 7201 8188
rect 7137 8128 7201 8132
rect 2584 7644 2648 7648
rect 2584 7588 2588 7644
rect 2588 7588 2644 7644
rect 2644 7588 2648 7644
rect 2584 7584 2648 7588
rect 2664 7644 2728 7648
rect 2664 7588 2668 7644
rect 2668 7588 2724 7644
rect 2724 7588 2728 7644
rect 2664 7584 2728 7588
rect 2744 7644 2808 7648
rect 2744 7588 2748 7644
rect 2748 7588 2804 7644
rect 2804 7588 2808 7644
rect 2744 7584 2808 7588
rect 2824 7644 2888 7648
rect 2824 7588 2828 7644
rect 2828 7588 2884 7644
rect 2884 7588 2888 7644
rect 2824 7584 2888 7588
rect 4309 7644 4373 7648
rect 4309 7588 4313 7644
rect 4313 7588 4369 7644
rect 4369 7588 4373 7644
rect 4309 7584 4373 7588
rect 4389 7644 4453 7648
rect 4389 7588 4393 7644
rect 4393 7588 4449 7644
rect 4449 7588 4453 7644
rect 4389 7584 4453 7588
rect 4469 7644 4533 7648
rect 4469 7588 4473 7644
rect 4473 7588 4529 7644
rect 4529 7588 4533 7644
rect 4469 7584 4533 7588
rect 4549 7644 4613 7648
rect 4549 7588 4553 7644
rect 4553 7588 4609 7644
rect 4609 7588 4613 7644
rect 4549 7584 4613 7588
rect 6034 7644 6098 7648
rect 6034 7588 6038 7644
rect 6038 7588 6094 7644
rect 6094 7588 6098 7644
rect 6034 7584 6098 7588
rect 6114 7644 6178 7648
rect 6114 7588 6118 7644
rect 6118 7588 6174 7644
rect 6174 7588 6178 7644
rect 6114 7584 6178 7588
rect 6194 7644 6258 7648
rect 6194 7588 6198 7644
rect 6198 7588 6254 7644
rect 6254 7588 6258 7644
rect 6194 7584 6258 7588
rect 6274 7644 6338 7648
rect 6274 7588 6278 7644
rect 6278 7588 6334 7644
rect 6334 7588 6338 7644
rect 6274 7584 6338 7588
rect 7759 7644 7823 7648
rect 7759 7588 7763 7644
rect 7763 7588 7819 7644
rect 7819 7588 7823 7644
rect 7759 7584 7823 7588
rect 7839 7644 7903 7648
rect 7839 7588 7843 7644
rect 7843 7588 7899 7644
rect 7899 7588 7903 7644
rect 7839 7584 7903 7588
rect 7919 7644 7983 7648
rect 7919 7588 7923 7644
rect 7923 7588 7979 7644
rect 7979 7588 7983 7644
rect 7919 7584 7983 7588
rect 7999 7644 8063 7648
rect 7999 7588 8003 7644
rect 8003 7588 8059 7644
rect 8059 7588 8063 7644
rect 7999 7584 8063 7588
rect 1722 7100 1786 7104
rect 1722 7044 1726 7100
rect 1726 7044 1782 7100
rect 1782 7044 1786 7100
rect 1722 7040 1786 7044
rect 1802 7100 1866 7104
rect 1802 7044 1806 7100
rect 1806 7044 1862 7100
rect 1862 7044 1866 7100
rect 1802 7040 1866 7044
rect 1882 7100 1946 7104
rect 1882 7044 1886 7100
rect 1886 7044 1942 7100
rect 1942 7044 1946 7100
rect 1882 7040 1946 7044
rect 1962 7100 2026 7104
rect 1962 7044 1966 7100
rect 1966 7044 2022 7100
rect 2022 7044 2026 7100
rect 1962 7040 2026 7044
rect 3447 7100 3511 7104
rect 3447 7044 3451 7100
rect 3451 7044 3507 7100
rect 3507 7044 3511 7100
rect 3447 7040 3511 7044
rect 3527 7100 3591 7104
rect 3527 7044 3531 7100
rect 3531 7044 3587 7100
rect 3587 7044 3591 7100
rect 3527 7040 3591 7044
rect 3607 7100 3671 7104
rect 3607 7044 3611 7100
rect 3611 7044 3667 7100
rect 3667 7044 3671 7100
rect 3607 7040 3671 7044
rect 3687 7100 3751 7104
rect 3687 7044 3691 7100
rect 3691 7044 3747 7100
rect 3747 7044 3751 7100
rect 3687 7040 3751 7044
rect 5172 7100 5236 7104
rect 5172 7044 5176 7100
rect 5176 7044 5232 7100
rect 5232 7044 5236 7100
rect 5172 7040 5236 7044
rect 5252 7100 5316 7104
rect 5252 7044 5256 7100
rect 5256 7044 5312 7100
rect 5312 7044 5316 7100
rect 5252 7040 5316 7044
rect 5332 7100 5396 7104
rect 5332 7044 5336 7100
rect 5336 7044 5392 7100
rect 5392 7044 5396 7100
rect 5332 7040 5396 7044
rect 5412 7100 5476 7104
rect 5412 7044 5416 7100
rect 5416 7044 5472 7100
rect 5472 7044 5476 7100
rect 5412 7040 5476 7044
rect 6897 7100 6961 7104
rect 6897 7044 6901 7100
rect 6901 7044 6957 7100
rect 6957 7044 6961 7100
rect 6897 7040 6961 7044
rect 6977 7100 7041 7104
rect 6977 7044 6981 7100
rect 6981 7044 7037 7100
rect 7037 7044 7041 7100
rect 6977 7040 7041 7044
rect 7057 7100 7121 7104
rect 7057 7044 7061 7100
rect 7061 7044 7117 7100
rect 7117 7044 7121 7100
rect 7057 7040 7121 7044
rect 7137 7100 7201 7104
rect 7137 7044 7141 7100
rect 7141 7044 7197 7100
rect 7197 7044 7201 7100
rect 7137 7040 7201 7044
rect 2584 6556 2648 6560
rect 2584 6500 2588 6556
rect 2588 6500 2644 6556
rect 2644 6500 2648 6556
rect 2584 6496 2648 6500
rect 2664 6556 2728 6560
rect 2664 6500 2668 6556
rect 2668 6500 2724 6556
rect 2724 6500 2728 6556
rect 2664 6496 2728 6500
rect 2744 6556 2808 6560
rect 2744 6500 2748 6556
rect 2748 6500 2804 6556
rect 2804 6500 2808 6556
rect 2744 6496 2808 6500
rect 2824 6556 2888 6560
rect 2824 6500 2828 6556
rect 2828 6500 2884 6556
rect 2884 6500 2888 6556
rect 2824 6496 2888 6500
rect 4309 6556 4373 6560
rect 4309 6500 4313 6556
rect 4313 6500 4369 6556
rect 4369 6500 4373 6556
rect 4309 6496 4373 6500
rect 4389 6556 4453 6560
rect 4389 6500 4393 6556
rect 4393 6500 4449 6556
rect 4449 6500 4453 6556
rect 4389 6496 4453 6500
rect 4469 6556 4533 6560
rect 4469 6500 4473 6556
rect 4473 6500 4529 6556
rect 4529 6500 4533 6556
rect 4469 6496 4533 6500
rect 4549 6556 4613 6560
rect 4549 6500 4553 6556
rect 4553 6500 4609 6556
rect 4609 6500 4613 6556
rect 4549 6496 4613 6500
rect 6034 6556 6098 6560
rect 6034 6500 6038 6556
rect 6038 6500 6094 6556
rect 6094 6500 6098 6556
rect 6034 6496 6098 6500
rect 6114 6556 6178 6560
rect 6114 6500 6118 6556
rect 6118 6500 6174 6556
rect 6174 6500 6178 6556
rect 6114 6496 6178 6500
rect 6194 6556 6258 6560
rect 6194 6500 6198 6556
rect 6198 6500 6254 6556
rect 6254 6500 6258 6556
rect 6194 6496 6258 6500
rect 6274 6556 6338 6560
rect 6274 6500 6278 6556
rect 6278 6500 6334 6556
rect 6334 6500 6338 6556
rect 6274 6496 6338 6500
rect 7759 6556 7823 6560
rect 7759 6500 7763 6556
rect 7763 6500 7819 6556
rect 7819 6500 7823 6556
rect 7759 6496 7823 6500
rect 7839 6556 7903 6560
rect 7839 6500 7843 6556
rect 7843 6500 7899 6556
rect 7899 6500 7903 6556
rect 7839 6496 7903 6500
rect 7919 6556 7983 6560
rect 7919 6500 7923 6556
rect 7923 6500 7979 6556
rect 7979 6500 7983 6556
rect 7919 6496 7983 6500
rect 7999 6556 8063 6560
rect 7999 6500 8003 6556
rect 8003 6500 8059 6556
rect 8059 6500 8063 6556
rect 7999 6496 8063 6500
rect 4108 6292 4172 6356
rect 1722 6012 1786 6016
rect 1722 5956 1726 6012
rect 1726 5956 1782 6012
rect 1782 5956 1786 6012
rect 1722 5952 1786 5956
rect 1802 6012 1866 6016
rect 1802 5956 1806 6012
rect 1806 5956 1862 6012
rect 1862 5956 1866 6012
rect 1802 5952 1866 5956
rect 1882 6012 1946 6016
rect 1882 5956 1886 6012
rect 1886 5956 1942 6012
rect 1942 5956 1946 6012
rect 1882 5952 1946 5956
rect 1962 6012 2026 6016
rect 1962 5956 1966 6012
rect 1966 5956 2022 6012
rect 2022 5956 2026 6012
rect 1962 5952 2026 5956
rect 3447 6012 3511 6016
rect 3447 5956 3451 6012
rect 3451 5956 3507 6012
rect 3507 5956 3511 6012
rect 3447 5952 3511 5956
rect 3527 6012 3591 6016
rect 3527 5956 3531 6012
rect 3531 5956 3587 6012
rect 3587 5956 3591 6012
rect 3527 5952 3591 5956
rect 3607 6012 3671 6016
rect 3607 5956 3611 6012
rect 3611 5956 3667 6012
rect 3667 5956 3671 6012
rect 3607 5952 3671 5956
rect 3687 6012 3751 6016
rect 3687 5956 3691 6012
rect 3691 5956 3747 6012
rect 3747 5956 3751 6012
rect 3687 5952 3751 5956
rect 5172 6012 5236 6016
rect 5172 5956 5176 6012
rect 5176 5956 5232 6012
rect 5232 5956 5236 6012
rect 5172 5952 5236 5956
rect 5252 6012 5316 6016
rect 5252 5956 5256 6012
rect 5256 5956 5312 6012
rect 5312 5956 5316 6012
rect 5252 5952 5316 5956
rect 5332 6012 5396 6016
rect 5332 5956 5336 6012
rect 5336 5956 5392 6012
rect 5392 5956 5396 6012
rect 5332 5952 5396 5956
rect 5412 6012 5476 6016
rect 5412 5956 5416 6012
rect 5416 5956 5472 6012
rect 5472 5956 5476 6012
rect 5412 5952 5476 5956
rect 6897 6012 6961 6016
rect 6897 5956 6901 6012
rect 6901 5956 6957 6012
rect 6957 5956 6961 6012
rect 6897 5952 6961 5956
rect 6977 6012 7041 6016
rect 6977 5956 6981 6012
rect 6981 5956 7037 6012
rect 7037 5956 7041 6012
rect 6977 5952 7041 5956
rect 7057 6012 7121 6016
rect 7057 5956 7061 6012
rect 7061 5956 7117 6012
rect 7117 5956 7121 6012
rect 7057 5952 7121 5956
rect 7137 6012 7201 6016
rect 7137 5956 7141 6012
rect 7141 5956 7197 6012
rect 7197 5956 7201 6012
rect 7137 5952 7201 5956
rect 5580 5748 5644 5812
rect 2584 5468 2648 5472
rect 2584 5412 2588 5468
rect 2588 5412 2644 5468
rect 2644 5412 2648 5468
rect 2584 5408 2648 5412
rect 2664 5468 2728 5472
rect 2664 5412 2668 5468
rect 2668 5412 2724 5468
rect 2724 5412 2728 5468
rect 2664 5408 2728 5412
rect 2744 5468 2808 5472
rect 2744 5412 2748 5468
rect 2748 5412 2804 5468
rect 2804 5412 2808 5468
rect 2744 5408 2808 5412
rect 2824 5468 2888 5472
rect 2824 5412 2828 5468
rect 2828 5412 2884 5468
rect 2884 5412 2888 5468
rect 2824 5408 2888 5412
rect 4309 5468 4373 5472
rect 4309 5412 4313 5468
rect 4313 5412 4369 5468
rect 4369 5412 4373 5468
rect 4309 5408 4373 5412
rect 4389 5468 4453 5472
rect 4389 5412 4393 5468
rect 4393 5412 4449 5468
rect 4449 5412 4453 5468
rect 4389 5408 4453 5412
rect 4469 5468 4533 5472
rect 4469 5412 4473 5468
rect 4473 5412 4529 5468
rect 4529 5412 4533 5468
rect 4469 5408 4533 5412
rect 4549 5468 4613 5472
rect 4549 5412 4553 5468
rect 4553 5412 4609 5468
rect 4609 5412 4613 5468
rect 4549 5408 4613 5412
rect 6034 5468 6098 5472
rect 6034 5412 6038 5468
rect 6038 5412 6094 5468
rect 6094 5412 6098 5468
rect 6034 5408 6098 5412
rect 6114 5468 6178 5472
rect 6114 5412 6118 5468
rect 6118 5412 6174 5468
rect 6174 5412 6178 5468
rect 6114 5408 6178 5412
rect 6194 5468 6258 5472
rect 6194 5412 6198 5468
rect 6198 5412 6254 5468
rect 6254 5412 6258 5468
rect 6194 5408 6258 5412
rect 6274 5468 6338 5472
rect 6274 5412 6278 5468
rect 6278 5412 6334 5468
rect 6334 5412 6338 5468
rect 6274 5408 6338 5412
rect 7759 5468 7823 5472
rect 7759 5412 7763 5468
rect 7763 5412 7819 5468
rect 7819 5412 7823 5468
rect 7759 5408 7823 5412
rect 7839 5468 7903 5472
rect 7839 5412 7843 5468
rect 7843 5412 7899 5468
rect 7899 5412 7903 5468
rect 7839 5408 7903 5412
rect 7919 5468 7983 5472
rect 7919 5412 7923 5468
rect 7923 5412 7979 5468
rect 7979 5412 7983 5468
rect 7919 5408 7983 5412
rect 7999 5468 8063 5472
rect 7999 5412 8003 5468
rect 8003 5412 8059 5468
rect 8059 5412 8063 5468
rect 7999 5408 8063 5412
rect 1722 4924 1786 4928
rect 1722 4868 1726 4924
rect 1726 4868 1782 4924
rect 1782 4868 1786 4924
rect 1722 4864 1786 4868
rect 1802 4924 1866 4928
rect 1802 4868 1806 4924
rect 1806 4868 1862 4924
rect 1862 4868 1866 4924
rect 1802 4864 1866 4868
rect 1882 4924 1946 4928
rect 1882 4868 1886 4924
rect 1886 4868 1942 4924
rect 1942 4868 1946 4924
rect 1882 4864 1946 4868
rect 1962 4924 2026 4928
rect 1962 4868 1966 4924
rect 1966 4868 2022 4924
rect 2022 4868 2026 4924
rect 1962 4864 2026 4868
rect 3447 4924 3511 4928
rect 3447 4868 3451 4924
rect 3451 4868 3507 4924
rect 3507 4868 3511 4924
rect 3447 4864 3511 4868
rect 3527 4924 3591 4928
rect 3527 4868 3531 4924
rect 3531 4868 3587 4924
rect 3587 4868 3591 4924
rect 3527 4864 3591 4868
rect 3607 4924 3671 4928
rect 3607 4868 3611 4924
rect 3611 4868 3667 4924
rect 3667 4868 3671 4924
rect 3607 4864 3671 4868
rect 3687 4924 3751 4928
rect 3687 4868 3691 4924
rect 3691 4868 3747 4924
rect 3747 4868 3751 4924
rect 3687 4864 3751 4868
rect 5172 4924 5236 4928
rect 5172 4868 5176 4924
rect 5176 4868 5232 4924
rect 5232 4868 5236 4924
rect 5172 4864 5236 4868
rect 5252 4924 5316 4928
rect 5252 4868 5256 4924
rect 5256 4868 5312 4924
rect 5312 4868 5316 4924
rect 5252 4864 5316 4868
rect 5332 4924 5396 4928
rect 5332 4868 5336 4924
rect 5336 4868 5392 4924
rect 5392 4868 5396 4924
rect 5332 4864 5396 4868
rect 5412 4924 5476 4928
rect 5412 4868 5416 4924
rect 5416 4868 5472 4924
rect 5472 4868 5476 4924
rect 5412 4864 5476 4868
rect 6897 4924 6961 4928
rect 6897 4868 6901 4924
rect 6901 4868 6957 4924
rect 6957 4868 6961 4924
rect 6897 4864 6961 4868
rect 6977 4924 7041 4928
rect 6977 4868 6981 4924
rect 6981 4868 7037 4924
rect 7037 4868 7041 4924
rect 6977 4864 7041 4868
rect 7057 4924 7121 4928
rect 7057 4868 7061 4924
rect 7061 4868 7117 4924
rect 7117 4868 7121 4924
rect 7057 4864 7121 4868
rect 7137 4924 7201 4928
rect 7137 4868 7141 4924
rect 7141 4868 7197 4924
rect 7197 4868 7201 4924
rect 7137 4864 7201 4868
rect 2584 4380 2648 4384
rect 2584 4324 2588 4380
rect 2588 4324 2644 4380
rect 2644 4324 2648 4380
rect 2584 4320 2648 4324
rect 2664 4380 2728 4384
rect 2664 4324 2668 4380
rect 2668 4324 2724 4380
rect 2724 4324 2728 4380
rect 2664 4320 2728 4324
rect 2744 4380 2808 4384
rect 2744 4324 2748 4380
rect 2748 4324 2804 4380
rect 2804 4324 2808 4380
rect 2744 4320 2808 4324
rect 2824 4380 2888 4384
rect 2824 4324 2828 4380
rect 2828 4324 2884 4380
rect 2884 4324 2888 4380
rect 2824 4320 2888 4324
rect 4309 4380 4373 4384
rect 4309 4324 4313 4380
rect 4313 4324 4369 4380
rect 4369 4324 4373 4380
rect 4309 4320 4373 4324
rect 4389 4380 4453 4384
rect 4389 4324 4393 4380
rect 4393 4324 4449 4380
rect 4449 4324 4453 4380
rect 4389 4320 4453 4324
rect 4469 4380 4533 4384
rect 4469 4324 4473 4380
rect 4473 4324 4529 4380
rect 4529 4324 4533 4380
rect 4469 4320 4533 4324
rect 4549 4380 4613 4384
rect 4549 4324 4553 4380
rect 4553 4324 4609 4380
rect 4609 4324 4613 4380
rect 4549 4320 4613 4324
rect 6034 4380 6098 4384
rect 6034 4324 6038 4380
rect 6038 4324 6094 4380
rect 6094 4324 6098 4380
rect 6034 4320 6098 4324
rect 6114 4380 6178 4384
rect 6114 4324 6118 4380
rect 6118 4324 6174 4380
rect 6174 4324 6178 4380
rect 6114 4320 6178 4324
rect 6194 4380 6258 4384
rect 6194 4324 6198 4380
rect 6198 4324 6254 4380
rect 6254 4324 6258 4380
rect 6194 4320 6258 4324
rect 6274 4380 6338 4384
rect 6274 4324 6278 4380
rect 6278 4324 6334 4380
rect 6334 4324 6338 4380
rect 6274 4320 6338 4324
rect 7759 4380 7823 4384
rect 7759 4324 7763 4380
rect 7763 4324 7819 4380
rect 7819 4324 7823 4380
rect 7759 4320 7823 4324
rect 7839 4380 7903 4384
rect 7839 4324 7843 4380
rect 7843 4324 7899 4380
rect 7899 4324 7903 4380
rect 7839 4320 7903 4324
rect 7919 4380 7983 4384
rect 7919 4324 7923 4380
rect 7923 4324 7979 4380
rect 7979 4324 7983 4380
rect 7919 4320 7983 4324
rect 7999 4380 8063 4384
rect 7999 4324 8003 4380
rect 8003 4324 8059 4380
rect 8059 4324 8063 4380
rect 7999 4320 8063 4324
rect 1722 3836 1786 3840
rect 1722 3780 1726 3836
rect 1726 3780 1782 3836
rect 1782 3780 1786 3836
rect 1722 3776 1786 3780
rect 1802 3836 1866 3840
rect 1802 3780 1806 3836
rect 1806 3780 1862 3836
rect 1862 3780 1866 3836
rect 1802 3776 1866 3780
rect 1882 3836 1946 3840
rect 1882 3780 1886 3836
rect 1886 3780 1942 3836
rect 1942 3780 1946 3836
rect 1882 3776 1946 3780
rect 1962 3836 2026 3840
rect 1962 3780 1966 3836
rect 1966 3780 2022 3836
rect 2022 3780 2026 3836
rect 1962 3776 2026 3780
rect 3447 3836 3511 3840
rect 3447 3780 3451 3836
rect 3451 3780 3507 3836
rect 3507 3780 3511 3836
rect 3447 3776 3511 3780
rect 3527 3836 3591 3840
rect 3527 3780 3531 3836
rect 3531 3780 3587 3836
rect 3587 3780 3591 3836
rect 3527 3776 3591 3780
rect 3607 3836 3671 3840
rect 3607 3780 3611 3836
rect 3611 3780 3667 3836
rect 3667 3780 3671 3836
rect 3607 3776 3671 3780
rect 3687 3836 3751 3840
rect 3687 3780 3691 3836
rect 3691 3780 3747 3836
rect 3747 3780 3751 3836
rect 3687 3776 3751 3780
rect 5172 3836 5236 3840
rect 5172 3780 5176 3836
rect 5176 3780 5232 3836
rect 5232 3780 5236 3836
rect 5172 3776 5236 3780
rect 5252 3836 5316 3840
rect 5252 3780 5256 3836
rect 5256 3780 5312 3836
rect 5312 3780 5316 3836
rect 5252 3776 5316 3780
rect 5332 3836 5396 3840
rect 5332 3780 5336 3836
rect 5336 3780 5392 3836
rect 5392 3780 5396 3836
rect 5332 3776 5396 3780
rect 5412 3836 5476 3840
rect 5412 3780 5416 3836
rect 5416 3780 5472 3836
rect 5472 3780 5476 3836
rect 5412 3776 5476 3780
rect 6897 3836 6961 3840
rect 6897 3780 6901 3836
rect 6901 3780 6957 3836
rect 6957 3780 6961 3836
rect 6897 3776 6961 3780
rect 6977 3836 7041 3840
rect 6977 3780 6981 3836
rect 6981 3780 7037 3836
rect 7037 3780 7041 3836
rect 6977 3776 7041 3780
rect 7057 3836 7121 3840
rect 7057 3780 7061 3836
rect 7061 3780 7117 3836
rect 7117 3780 7121 3836
rect 7057 3776 7121 3780
rect 7137 3836 7201 3840
rect 7137 3780 7141 3836
rect 7141 3780 7197 3836
rect 7197 3780 7201 3836
rect 7137 3776 7201 3780
rect 2584 3292 2648 3296
rect 2584 3236 2588 3292
rect 2588 3236 2644 3292
rect 2644 3236 2648 3292
rect 2584 3232 2648 3236
rect 2664 3292 2728 3296
rect 2664 3236 2668 3292
rect 2668 3236 2724 3292
rect 2724 3236 2728 3292
rect 2664 3232 2728 3236
rect 2744 3292 2808 3296
rect 2744 3236 2748 3292
rect 2748 3236 2804 3292
rect 2804 3236 2808 3292
rect 2744 3232 2808 3236
rect 2824 3292 2888 3296
rect 2824 3236 2828 3292
rect 2828 3236 2884 3292
rect 2884 3236 2888 3292
rect 2824 3232 2888 3236
rect 4309 3292 4373 3296
rect 4309 3236 4313 3292
rect 4313 3236 4369 3292
rect 4369 3236 4373 3292
rect 4309 3232 4373 3236
rect 4389 3292 4453 3296
rect 4389 3236 4393 3292
rect 4393 3236 4449 3292
rect 4449 3236 4453 3292
rect 4389 3232 4453 3236
rect 4469 3292 4533 3296
rect 4469 3236 4473 3292
rect 4473 3236 4529 3292
rect 4529 3236 4533 3292
rect 4469 3232 4533 3236
rect 4549 3292 4613 3296
rect 4549 3236 4553 3292
rect 4553 3236 4609 3292
rect 4609 3236 4613 3292
rect 4549 3232 4613 3236
rect 6034 3292 6098 3296
rect 6034 3236 6038 3292
rect 6038 3236 6094 3292
rect 6094 3236 6098 3292
rect 6034 3232 6098 3236
rect 6114 3292 6178 3296
rect 6114 3236 6118 3292
rect 6118 3236 6174 3292
rect 6174 3236 6178 3292
rect 6114 3232 6178 3236
rect 6194 3292 6258 3296
rect 6194 3236 6198 3292
rect 6198 3236 6254 3292
rect 6254 3236 6258 3292
rect 6194 3232 6258 3236
rect 6274 3292 6338 3296
rect 6274 3236 6278 3292
rect 6278 3236 6334 3292
rect 6334 3236 6338 3292
rect 6274 3232 6338 3236
rect 7759 3292 7823 3296
rect 7759 3236 7763 3292
rect 7763 3236 7819 3292
rect 7819 3236 7823 3292
rect 7759 3232 7823 3236
rect 7839 3292 7903 3296
rect 7839 3236 7843 3292
rect 7843 3236 7899 3292
rect 7899 3236 7903 3292
rect 7839 3232 7903 3236
rect 7919 3292 7983 3296
rect 7919 3236 7923 3292
rect 7923 3236 7979 3292
rect 7979 3236 7983 3292
rect 7919 3232 7983 3236
rect 7999 3292 8063 3296
rect 7999 3236 8003 3292
rect 8003 3236 8059 3292
rect 8059 3236 8063 3292
rect 7999 3232 8063 3236
rect 4108 3028 4172 3092
rect 1722 2748 1786 2752
rect 1722 2692 1726 2748
rect 1726 2692 1782 2748
rect 1782 2692 1786 2748
rect 1722 2688 1786 2692
rect 1802 2748 1866 2752
rect 1802 2692 1806 2748
rect 1806 2692 1862 2748
rect 1862 2692 1866 2748
rect 1802 2688 1866 2692
rect 1882 2748 1946 2752
rect 1882 2692 1886 2748
rect 1886 2692 1942 2748
rect 1942 2692 1946 2748
rect 1882 2688 1946 2692
rect 1962 2748 2026 2752
rect 1962 2692 1966 2748
rect 1966 2692 2022 2748
rect 2022 2692 2026 2748
rect 1962 2688 2026 2692
rect 3447 2748 3511 2752
rect 3447 2692 3451 2748
rect 3451 2692 3507 2748
rect 3507 2692 3511 2748
rect 3447 2688 3511 2692
rect 3527 2748 3591 2752
rect 3527 2692 3531 2748
rect 3531 2692 3587 2748
rect 3587 2692 3591 2748
rect 3527 2688 3591 2692
rect 3607 2748 3671 2752
rect 3607 2692 3611 2748
rect 3611 2692 3667 2748
rect 3667 2692 3671 2748
rect 3607 2688 3671 2692
rect 3687 2748 3751 2752
rect 3687 2692 3691 2748
rect 3691 2692 3747 2748
rect 3747 2692 3751 2748
rect 3687 2688 3751 2692
rect 5172 2748 5236 2752
rect 5172 2692 5176 2748
rect 5176 2692 5232 2748
rect 5232 2692 5236 2748
rect 5172 2688 5236 2692
rect 5252 2748 5316 2752
rect 5252 2692 5256 2748
rect 5256 2692 5312 2748
rect 5312 2692 5316 2748
rect 5252 2688 5316 2692
rect 5332 2748 5396 2752
rect 5332 2692 5336 2748
rect 5336 2692 5392 2748
rect 5392 2692 5396 2748
rect 5332 2688 5396 2692
rect 5412 2748 5476 2752
rect 5412 2692 5416 2748
rect 5416 2692 5472 2748
rect 5472 2692 5476 2748
rect 5412 2688 5476 2692
rect 6897 2748 6961 2752
rect 6897 2692 6901 2748
rect 6901 2692 6957 2748
rect 6957 2692 6961 2748
rect 6897 2688 6961 2692
rect 6977 2748 7041 2752
rect 6977 2692 6981 2748
rect 6981 2692 7037 2748
rect 7037 2692 7041 2748
rect 6977 2688 7041 2692
rect 7057 2748 7121 2752
rect 7057 2692 7061 2748
rect 7061 2692 7117 2748
rect 7117 2692 7121 2748
rect 7057 2688 7121 2692
rect 7137 2748 7201 2752
rect 7137 2692 7141 2748
rect 7141 2692 7197 2748
rect 7197 2692 7201 2748
rect 7137 2688 7201 2692
rect 2584 2204 2648 2208
rect 2584 2148 2588 2204
rect 2588 2148 2644 2204
rect 2644 2148 2648 2204
rect 2584 2144 2648 2148
rect 2664 2204 2728 2208
rect 2664 2148 2668 2204
rect 2668 2148 2724 2204
rect 2724 2148 2728 2204
rect 2664 2144 2728 2148
rect 2744 2204 2808 2208
rect 2744 2148 2748 2204
rect 2748 2148 2804 2204
rect 2804 2148 2808 2204
rect 2744 2144 2808 2148
rect 2824 2204 2888 2208
rect 2824 2148 2828 2204
rect 2828 2148 2884 2204
rect 2884 2148 2888 2204
rect 2824 2144 2888 2148
rect 4309 2204 4373 2208
rect 4309 2148 4313 2204
rect 4313 2148 4369 2204
rect 4369 2148 4373 2204
rect 4309 2144 4373 2148
rect 4389 2204 4453 2208
rect 4389 2148 4393 2204
rect 4393 2148 4449 2204
rect 4449 2148 4453 2204
rect 4389 2144 4453 2148
rect 4469 2204 4533 2208
rect 4469 2148 4473 2204
rect 4473 2148 4529 2204
rect 4529 2148 4533 2204
rect 4469 2144 4533 2148
rect 4549 2204 4613 2208
rect 4549 2148 4553 2204
rect 4553 2148 4609 2204
rect 4609 2148 4613 2204
rect 4549 2144 4613 2148
rect 6034 2204 6098 2208
rect 6034 2148 6038 2204
rect 6038 2148 6094 2204
rect 6094 2148 6098 2204
rect 6034 2144 6098 2148
rect 6114 2204 6178 2208
rect 6114 2148 6118 2204
rect 6118 2148 6174 2204
rect 6174 2148 6178 2204
rect 6114 2144 6178 2148
rect 6194 2204 6258 2208
rect 6194 2148 6198 2204
rect 6198 2148 6254 2204
rect 6254 2148 6258 2204
rect 6194 2144 6258 2148
rect 6274 2204 6338 2208
rect 6274 2148 6278 2204
rect 6278 2148 6334 2204
rect 6334 2148 6338 2204
rect 6274 2144 6338 2148
rect 7759 2204 7823 2208
rect 7759 2148 7763 2204
rect 7763 2148 7819 2204
rect 7819 2148 7823 2204
rect 7759 2144 7823 2148
rect 7839 2204 7903 2208
rect 7839 2148 7843 2204
rect 7843 2148 7899 2204
rect 7899 2148 7903 2204
rect 7839 2144 7903 2148
rect 7919 2204 7983 2208
rect 7919 2148 7923 2204
rect 7923 2148 7979 2204
rect 7979 2148 7983 2204
rect 7919 2144 7983 2148
rect 7999 2204 8063 2208
rect 7999 2148 8003 2204
rect 8003 2148 8059 2204
rect 8059 2148 8063 2204
rect 7999 2144 8063 2148
rect 1722 1660 1786 1664
rect 1722 1604 1726 1660
rect 1726 1604 1782 1660
rect 1782 1604 1786 1660
rect 1722 1600 1786 1604
rect 1802 1660 1866 1664
rect 1802 1604 1806 1660
rect 1806 1604 1862 1660
rect 1862 1604 1866 1660
rect 1802 1600 1866 1604
rect 1882 1660 1946 1664
rect 1882 1604 1886 1660
rect 1886 1604 1942 1660
rect 1942 1604 1946 1660
rect 1882 1600 1946 1604
rect 1962 1660 2026 1664
rect 1962 1604 1966 1660
rect 1966 1604 2022 1660
rect 2022 1604 2026 1660
rect 1962 1600 2026 1604
rect 3447 1660 3511 1664
rect 3447 1604 3451 1660
rect 3451 1604 3507 1660
rect 3507 1604 3511 1660
rect 3447 1600 3511 1604
rect 3527 1660 3591 1664
rect 3527 1604 3531 1660
rect 3531 1604 3587 1660
rect 3587 1604 3591 1660
rect 3527 1600 3591 1604
rect 3607 1660 3671 1664
rect 3607 1604 3611 1660
rect 3611 1604 3667 1660
rect 3667 1604 3671 1660
rect 3607 1600 3671 1604
rect 3687 1660 3751 1664
rect 3687 1604 3691 1660
rect 3691 1604 3747 1660
rect 3747 1604 3751 1660
rect 3687 1600 3751 1604
rect 5172 1660 5236 1664
rect 5172 1604 5176 1660
rect 5176 1604 5232 1660
rect 5232 1604 5236 1660
rect 5172 1600 5236 1604
rect 5252 1660 5316 1664
rect 5252 1604 5256 1660
rect 5256 1604 5312 1660
rect 5312 1604 5316 1660
rect 5252 1600 5316 1604
rect 5332 1660 5396 1664
rect 5332 1604 5336 1660
rect 5336 1604 5392 1660
rect 5392 1604 5396 1660
rect 5332 1600 5396 1604
rect 5412 1660 5476 1664
rect 5412 1604 5416 1660
rect 5416 1604 5472 1660
rect 5472 1604 5476 1660
rect 5412 1600 5476 1604
rect 6897 1660 6961 1664
rect 6897 1604 6901 1660
rect 6901 1604 6957 1660
rect 6957 1604 6961 1660
rect 6897 1600 6961 1604
rect 6977 1660 7041 1664
rect 6977 1604 6981 1660
rect 6981 1604 7037 1660
rect 7037 1604 7041 1660
rect 6977 1600 7041 1604
rect 7057 1660 7121 1664
rect 7057 1604 7061 1660
rect 7061 1604 7117 1660
rect 7117 1604 7121 1660
rect 7057 1600 7121 1604
rect 7137 1660 7201 1664
rect 7137 1604 7141 1660
rect 7141 1604 7197 1660
rect 7197 1604 7201 1660
rect 7137 1600 7201 1604
rect 2584 1116 2648 1120
rect 2584 1060 2588 1116
rect 2588 1060 2644 1116
rect 2644 1060 2648 1116
rect 2584 1056 2648 1060
rect 2664 1116 2728 1120
rect 2664 1060 2668 1116
rect 2668 1060 2724 1116
rect 2724 1060 2728 1116
rect 2664 1056 2728 1060
rect 2744 1116 2808 1120
rect 2744 1060 2748 1116
rect 2748 1060 2804 1116
rect 2804 1060 2808 1116
rect 2744 1056 2808 1060
rect 2824 1116 2888 1120
rect 2824 1060 2828 1116
rect 2828 1060 2884 1116
rect 2884 1060 2888 1116
rect 2824 1056 2888 1060
rect 4309 1116 4373 1120
rect 4309 1060 4313 1116
rect 4313 1060 4369 1116
rect 4369 1060 4373 1116
rect 4309 1056 4373 1060
rect 4389 1116 4453 1120
rect 4389 1060 4393 1116
rect 4393 1060 4449 1116
rect 4449 1060 4453 1116
rect 4389 1056 4453 1060
rect 4469 1116 4533 1120
rect 4469 1060 4473 1116
rect 4473 1060 4529 1116
rect 4529 1060 4533 1116
rect 4469 1056 4533 1060
rect 4549 1116 4613 1120
rect 4549 1060 4553 1116
rect 4553 1060 4609 1116
rect 4609 1060 4613 1116
rect 4549 1056 4613 1060
rect 6034 1116 6098 1120
rect 6034 1060 6038 1116
rect 6038 1060 6094 1116
rect 6094 1060 6098 1116
rect 6034 1056 6098 1060
rect 6114 1116 6178 1120
rect 6114 1060 6118 1116
rect 6118 1060 6174 1116
rect 6174 1060 6178 1116
rect 6114 1056 6178 1060
rect 6194 1116 6258 1120
rect 6194 1060 6198 1116
rect 6198 1060 6254 1116
rect 6254 1060 6258 1116
rect 6194 1056 6258 1060
rect 6274 1116 6338 1120
rect 6274 1060 6278 1116
rect 6278 1060 6334 1116
rect 6334 1060 6338 1116
rect 6274 1056 6338 1060
rect 7759 1116 7823 1120
rect 7759 1060 7763 1116
rect 7763 1060 7819 1116
rect 7819 1060 7823 1116
rect 7759 1056 7823 1060
rect 7839 1116 7903 1120
rect 7839 1060 7843 1116
rect 7843 1060 7899 1116
rect 7899 1060 7903 1116
rect 7839 1056 7903 1060
rect 7919 1116 7983 1120
rect 7919 1060 7923 1116
rect 7923 1060 7979 1116
rect 7979 1060 7983 1116
rect 7919 1056 7983 1060
rect 7999 1116 8063 1120
rect 7999 1060 8003 1116
rect 8003 1060 8059 1116
rect 8059 1060 8063 1116
rect 7999 1056 8063 1060
<< metal4 >>
rect 5579 9212 5645 9213
rect 5579 9148 5580 9212
rect 5644 9148 5645 9212
rect 5579 9147 5645 9148
rect 1714 8192 2034 8752
rect 1714 8128 1722 8192
rect 1786 8128 1802 8192
rect 1866 8128 1882 8192
rect 1946 8128 1962 8192
rect 2026 8128 2034 8192
rect 1714 7104 2034 8128
rect 1714 7040 1722 7104
rect 1786 7040 1802 7104
rect 1866 7040 1882 7104
rect 1946 7040 1962 7104
rect 2026 7040 2034 7104
rect 1714 6016 2034 7040
rect 1714 5952 1722 6016
rect 1786 5952 1802 6016
rect 1866 5952 1882 6016
rect 1946 5952 1962 6016
rect 2026 5952 2034 6016
rect 1714 4928 2034 5952
rect 1714 4864 1722 4928
rect 1786 4864 1802 4928
rect 1866 4864 1882 4928
rect 1946 4864 1962 4928
rect 2026 4864 2034 4928
rect 1714 3840 2034 4864
rect 1714 3776 1722 3840
rect 1786 3776 1802 3840
rect 1866 3776 1882 3840
rect 1946 3776 1962 3840
rect 2026 3776 2034 3840
rect 1714 2752 2034 3776
rect 1714 2688 1722 2752
rect 1786 2688 1802 2752
rect 1866 2688 1882 2752
rect 1946 2688 1962 2752
rect 2026 2688 2034 2752
rect 1714 1664 2034 2688
rect 1714 1600 1722 1664
rect 1786 1600 1802 1664
rect 1866 1600 1882 1664
rect 1946 1600 1962 1664
rect 2026 1600 2034 1664
rect 1714 1040 2034 1600
rect 2576 8736 2896 8752
rect 2576 8672 2584 8736
rect 2648 8672 2664 8736
rect 2728 8672 2744 8736
rect 2808 8672 2824 8736
rect 2888 8672 2896 8736
rect 2576 7648 2896 8672
rect 2576 7584 2584 7648
rect 2648 7584 2664 7648
rect 2728 7584 2744 7648
rect 2808 7584 2824 7648
rect 2888 7584 2896 7648
rect 2576 6560 2896 7584
rect 2576 6496 2584 6560
rect 2648 6496 2664 6560
rect 2728 6496 2744 6560
rect 2808 6496 2824 6560
rect 2888 6496 2896 6560
rect 2576 5472 2896 6496
rect 2576 5408 2584 5472
rect 2648 5408 2664 5472
rect 2728 5408 2744 5472
rect 2808 5408 2824 5472
rect 2888 5408 2896 5472
rect 2576 4384 2896 5408
rect 2576 4320 2584 4384
rect 2648 4320 2664 4384
rect 2728 4320 2744 4384
rect 2808 4320 2824 4384
rect 2888 4320 2896 4384
rect 2576 3296 2896 4320
rect 2576 3232 2584 3296
rect 2648 3232 2664 3296
rect 2728 3232 2744 3296
rect 2808 3232 2824 3296
rect 2888 3232 2896 3296
rect 2576 2208 2896 3232
rect 2576 2144 2584 2208
rect 2648 2144 2664 2208
rect 2728 2144 2744 2208
rect 2808 2144 2824 2208
rect 2888 2144 2896 2208
rect 2576 1120 2896 2144
rect 2576 1056 2584 1120
rect 2648 1056 2664 1120
rect 2728 1056 2744 1120
rect 2808 1056 2824 1120
rect 2888 1056 2896 1120
rect 2576 1040 2896 1056
rect 3439 8192 3759 8752
rect 3439 8128 3447 8192
rect 3511 8128 3527 8192
rect 3591 8128 3607 8192
rect 3671 8128 3687 8192
rect 3751 8128 3759 8192
rect 3439 7104 3759 8128
rect 3439 7040 3447 7104
rect 3511 7040 3527 7104
rect 3591 7040 3607 7104
rect 3671 7040 3687 7104
rect 3751 7040 3759 7104
rect 3439 6016 3759 7040
rect 4301 8736 4621 8752
rect 4301 8672 4309 8736
rect 4373 8672 4389 8736
rect 4453 8672 4469 8736
rect 4533 8672 4549 8736
rect 4613 8672 4621 8736
rect 4301 7648 4621 8672
rect 4301 7584 4309 7648
rect 4373 7584 4389 7648
rect 4453 7584 4469 7648
rect 4533 7584 4549 7648
rect 4613 7584 4621 7648
rect 4301 6560 4621 7584
rect 4301 6496 4309 6560
rect 4373 6496 4389 6560
rect 4453 6496 4469 6560
rect 4533 6496 4549 6560
rect 4613 6496 4621 6560
rect 4107 6356 4173 6357
rect 4107 6292 4108 6356
rect 4172 6292 4173 6356
rect 4107 6291 4173 6292
rect 3439 5952 3447 6016
rect 3511 5952 3527 6016
rect 3591 5952 3607 6016
rect 3671 5952 3687 6016
rect 3751 5952 3759 6016
rect 3439 4928 3759 5952
rect 3439 4864 3447 4928
rect 3511 4864 3527 4928
rect 3591 4864 3607 4928
rect 3671 4864 3687 4928
rect 3751 4864 3759 4928
rect 3439 3840 3759 4864
rect 3439 3776 3447 3840
rect 3511 3776 3527 3840
rect 3591 3776 3607 3840
rect 3671 3776 3687 3840
rect 3751 3776 3759 3840
rect 3439 2752 3759 3776
rect 4110 3093 4170 6291
rect 4301 5472 4621 6496
rect 4301 5408 4309 5472
rect 4373 5408 4389 5472
rect 4453 5408 4469 5472
rect 4533 5408 4549 5472
rect 4613 5408 4621 5472
rect 4301 4384 4621 5408
rect 4301 4320 4309 4384
rect 4373 4320 4389 4384
rect 4453 4320 4469 4384
rect 4533 4320 4549 4384
rect 4613 4320 4621 4384
rect 4301 3296 4621 4320
rect 4301 3232 4309 3296
rect 4373 3232 4389 3296
rect 4453 3232 4469 3296
rect 4533 3232 4549 3296
rect 4613 3232 4621 3296
rect 4107 3092 4173 3093
rect 4107 3028 4108 3092
rect 4172 3028 4173 3092
rect 4107 3027 4173 3028
rect 3439 2688 3447 2752
rect 3511 2688 3527 2752
rect 3591 2688 3607 2752
rect 3671 2688 3687 2752
rect 3751 2688 3759 2752
rect 3439 1664 3759 2688
rect 3439 1600 3447 1664
rect 3511 1600 3527 1664
rect 3591 1600 3607 1664
rect 3671 1600 3687 1664
rect 3751 1600 3759 1664
rect 3439 1040 3759 1600
rect 4301 2208 4621 3232
rect 4301 2144 4309 2208
rect 4373 2144 4389 2208
rect 4453 2144 4469 2208
rect 4533 2144 4549 2208
rect 4613 2144 4621 2208
rect 4301 1120 4621 2144
rect 4301 1056 4309 1120
rect 4373 1056 4389 1120
rect 4453 1056 4469 1120
rect 4533 1056 4549 1120
rect 4613 1056 4621 1120
rect 4301 1040 4621 1056
rect 5164 8192 5484 8752
rect 5164 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5484 8192
rect 5164 7104 5484 8128
rect 5164 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5484 7104
rect 5164 6016 5484 7040
rect 5164 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5484 6016
rect 5164 4928 5484 5952
rect 5582 5813 5642 9147
rect 6026 8736 6346 8752
rect 6026 8672 6034 8736
rect 6098 8672 6114 8736
rect 6178 8672 6194 8736
rect 6258 8672 6274 8736
rect 6338 8672 6346 8736
rect 6026 7648 6346 8672
rect 6026 7584 6034 7648
rect 6098 7584 6114 7648
rect 6178 7584 6194 7648
rect 6258 7584 6274 7648
rect 6338 7584 6346 7648
rect 6026 6560 6346 7584
rect 6026 6496 6034 6560
rect 6098 6496 6114 6560
rect 6178 6496 6194 6560
rect 6258 6496 6274 6560
rect 6338 6496 6346 6560
rect 5579 5812 5645 5813
rect 5579 5748 5580 5812
rect 5644 5748 5645 5812
rect 5579 5747 5645 5748
rect 5164 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5484 4928
rect 5164 3840 5484 4864
rect 5164 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5484 3840
rect 5164 2752 5484 3776
rect 5164 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5484 2752
rect 5164 1664 5484 2688
rect 5164 1600 5172 1664
rect 5236 1600 5252 1664
rect 5316 1600 5332 1664
rect 5396 1600 5412 1664
rect 5476 1600 5484 1664
rect 5164 1040 5484 1600
rect 6026 5472 6346 6496
rect 6026 5408 6034 5472
rect 6098 5408 6114 5472
rect 6178 5408 6194 5472
rect 6258 5408 6274 5472
rect 6338 5408 6346 5472
rect 6026 4384 6346 5408
rect 6026 4320 6034 4384
rect 6098 4320 6114 4384
rect 6178 4320 6194 4384
rect 6258 4320 6274 4384
rect 6338 4320 6346 4384
rect 6026 3296 6346 4320
rect 6026 3232 6034 3296
rect 6098 3232 6114 3296
rect 6178 3232 6194 3296
rect 6258 3232 6274 3296
rect 6338 3232 6346 3296
rect 6026 2208 6346 3232
rect 6026 2144 6034 2208
rect 6098 2144 6114 2208
rect 6178 2144 6194 2208
rect 6258 2144 6274 2208
rect 6338 2144 6346 2208
rect 6026 1120 6346 2144
rect 6026 1056 6034 1120
rect 6098 1056 6114 1120
rect 6178 1056 6194 1120
rect 6258 1056 6274 1120
rect 6338 1056 6346 1120
rect 6026 1040 6346 1056
rect 6889 8192 7209 8752
rect 6889 8128 6897 8192
rect 6961 8128 6977 8192
rect 7041 8128 7057 8192
rect 7121 8128 7137 8192
rect 7201 8128 7209 8192
rect 6889 7104 7209 8128
rect 6889 7040 6897 7104
rect 6961 7040 6977 7104
rect 7041 7040 7057 7104
rect 7121 7040 7137 7104
rect 7201 7040 7209 7104
rect 6889 6016 7209 7040
rect 6889 5952 6897 6016
rect 6961 5952 6977 6016
rect 7041 5952 7057 6016
rect 7121 5952 7137 6016
rect 7201 5952 7209 6016
rect 6889 4928 7209 5952
rect 6889 4864 6897 4928
rect 6961 4864 6977 4928
rect 7041 4864 7057 4928
rect 7121 4864 7137 4928
rect 7201 4864 7209 4928
rect 6889 3840 7209 4864
rect 6889 3776 6897 3840
rect 6961 3776 6977 3840
rect 7041 3776 7057 3840
rect 7121 3776 7137 3840
rect 7201 3776 7209 3840
rect 6889 2752 7209 3776
rect 6889 2688 6897 2752
rect 6961 2688 6977 2752
rect 7041 2688 7057 2752
rect 7121 2688 7137 2752
rect 7201 2688 7209 2752
rect 6889 1664 7209 2688
rect 6889 1600 6897 1664
rect 6961 1600 6977 1664
rect 7041 1600 7057 1664
rect 7121 1600 7137 1664
rect 7201 1600 7209 1664
rect 6889 1040 7209 1600
rect 7751 8736 8071 8752
rect 7751 8672 7759 8736
rect 7823 8672 7839 8736
rect 7903 8672 7919 8736
rect 7983 8672 7999 8736
rect 8063 8672 8071 8736
rect 7751 7648 8071 8672
rect 7751 7584 7759 7648
rect 7823 7584 7839 7648
rect 7903 7584 7919 7648
rect 7983 7584 7999 7648
rect 8063 7584 8071 7648
rect 7751 6560 8071 7584
rect 7751 6496 7759 6560
rect 7823 6496 7839 6560
rect 7903 6496 7919 6560
rect 7983 6496 7999 6560
rect 8063 6496 8071 6560
rect 7751 5472 8071 6496
rect 7751 5408 7759 5472
rect 7823 5408 7839 5472
rect 7903 5408 7919 5472
rect 7983 5408 7999 5472
rect 8063 5408 8071 5472
rect 7751 4384 8071 5408
rect 7751 4320 7759 4384
rect 7823 4320 7839 4384
rect 7903 4320 7919 4384
rect 7983 4320 7999 4384
rect 8063 4320 8071 4384
rect 7751 3296 8071 4320
rect 7751 3232 7759 3296
rect 7823 3232 7839 3296
rect 7903 3232 7919 3296
rect 7983 3232 7999 3296
rect 8063 3232 8071 3296
rect 7751 2208 8071 3232
rect 7751 2144 7759 2208
rect 7823 2144 7839 2208
rect 7903 2144 7919 2208
rect 7983 2144 7999 2208
rect 8063 2144 8071 2208
rect 7751 1120 8071 2144
rect 7751 1056 7759 1120
rect 7823 1056 7839 1120
rect 7903 1056 7919 1120
rect 7983 1056 7999 1120
rect 8063 1056 8071 1120
rect 7751 1040 8071 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[0\]_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[1\]_A
timestamp 1673029049
transform 1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[2\]_A
timestamp 1673029049
transform -1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[3\]_A
timestamp 1673029049
transform 1 0 3864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[4\]_A
timestamp 1673029049
transform -1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[5\]_A
timestamp 1673029049
transform -1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[6\]_A
timestamp 1673029049
transform -1 0 7360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[7\]_A
timestamp 1673029049
transform -1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[8\]_A
timestamp 1673029049
transform -1 0 4140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[9\]_A
timestamp 1673029049
transform -1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[10\]_A
timestamp 1673029049
transform -1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[11\]_A
timestamp 1673029049
transform -1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[12\]_A
timestamp 1673029049
transform -1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[13\]_A
timestamp 1673029049
transform -1 0 2852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[14\]_A
timestamp 1673029049
transform -1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[15\]_A
timestamp 1673029049
transform -1 0 1656 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[16\]_A
timestamp 1673029049
transform -1 0 5428 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[17\]_A
timestamp 1673029049
transform 1 0 5336 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[18\]_A
timestamp 1673029049
transform -1 0 2024 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[19\]_A
timestamp 1673029049
transform -1 0 6808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[20\]_A
timestamp 1673029049
transform 1 0 7268 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[21\]_A
timestamp 1673029049
transform 1 0 5796 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[22\]_A
timestamp 1673029049
transform -1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[23\]_A
timestamp 1673029049
transform -1 0 6900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[24\]_A
timestamp 1673029049
transform -1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[25\]_A
timestamp 1673029049
transform -1 0 5980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[26\]_A
timestamp 1673029049
transform -1 0 5980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[27\]_A
timestamp 1673029049
transform -1 0 6900 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[28\]_A
timestamp 1673029049
transform -1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[29\]_A
timestamp 1673029049
transform -1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[30\]_A
timestamp 1673029049
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[31\]_A
timestamp 1673029049
transform -1 0 2024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[32\]_A
timestamp 1673029049
transform 1 0 3864 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[33\]_A
timestamp 1673029049
transform -1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[34\]_A
timestamp 1673029049
transform -1 0 1840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[35\]_A
timestamp 1673029049
transform -1 0 1656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[36\]_A
timestamp 1673029049
transform -1 0 2208 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[37\]_A
timestamp 1673029049
transform -1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[38\]_A
timestamp 1673029049
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[39\]_A
timestamp 1673029049
transform 1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_BUF\[40\]_A
timestamp 1673029049
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 4232 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[1\]
timestamp 1673029049
transform 1 0 3312 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[2\]
timestamp 1673029049
transform 1 0 4876 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[3\]
timestamp 1673029049
transform 1 0 4692 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[4\]
timestamp 1673029049
transform 1 0 4416 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[5\]
timestamp 1673029049
transform 1 0 4140 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[6\]
timestamp 1673029049
transform 1 0 3864 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[7\]
timestamp 1673029049
transform 1 0 2392 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[8\]
timestamp 1673029049
transform -1 0 4048 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[9\]
timestamp 1673029049
transform 1 0 1932 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[10\]
timestamp 1673029049
transform -1 0 3404 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[11\]
timestamp 1673029049
transform -1 0 3772 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[12\]
timestamp 1673029049
transform -1 0 3404 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[13\]
timestamp 1673029049
transform -1 0 2668 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[14\]
timestamp 1673029049
transform -1 0 3680 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[15\]
timestamp 1673029049
transform -1 0 3404 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[16\]
timestamp 1673029049
transform -1 0 4876 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[17\]
timestamp 1673029049
transform -1 0 4968 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[18\]
timestamp 1673029049
transform -1 0 3588 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[19\]
timestamp 1673029049
transform -1 0 6256 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[20\]
timestamp 1673029049
transform -1 0 7452 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[21\]
timestamp 1673029049
transform -1 0 3404 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[22\]
timestamp 1673029049
transform -1 0 7452 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[23\]
timestamp 1673029049
transform -1 0 7452 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[24\]
timestamp 1673029049
transform -1 0 7452 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[25\]
timestamp 1673029049
transform 1 0 6440 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[26\]
timestamp 1673029049
transform -1 0 5520 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[27\]
timestamp 1673029049
transform 1 0 6440 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[28\]
timestamp 1673029049
transform 1 0 5888 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[29\]
timestamp 1673029049
transform 1 0 6440 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[30\]
timestamp 1673029049
transform 1 0 4968 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[31\]
timestamp 1673029049
transform 1 0 6440 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[32\]
timestamp 1673029049
transform 1 0 5336 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[33\]
timestamp 1673029049
transform 1 0 4968 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[34\]
timestamp 1673029049
transform 1 0 3956 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[35\]
timestamp 1673029049
transform 1 0 2392 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[36\]
timestamp 1673029049
transform 1 0 2392 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[37\]
timestamp 1673029049
transform 1 0 2208 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[38\]
timestamp 1673029049
transform 1 0 3588 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[39\]
timestamp 1673029049
transform 1 0 4416 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[40\]
timestamp 1673029049
transform 1 0 4692 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 1288 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 2024 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3404 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1673029049
transform 1 0 3680 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42
timestamp 1673029049
transform 1 0 4876 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48
timestamp 1673029049
transform 1 0 5428 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1673029049
transform 1 0 5980 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6256 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6992 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1673029049
transform 1 0 7452 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1673029049
transform 1 0 1288 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1673029049
transform 1 0 1656 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1673029049
transform 1 0 2208 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1673029049
transform 1 0 3588 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1673029049
transform 1 0 4968 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1673029049
transform 1 0 5520 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 6072 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1673029049
transform 1 0 6256 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 1673029049
transform 1 0 7452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1673029049
transform 1 0 1288 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1673029049
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1673029049
transform 1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1673029049
transform 1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1673029049
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1673029049
transform 1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1673029049
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_69
timestamp 1673029049
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1673029049
transform 1 0 1288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1673029049
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1673029049
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1673029049
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_33
timestamp 1673029049
transform 1 0 4048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_45
timestamp 1673029049
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1673029049
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1673029049
transform 1 0 6072 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1673029049
transform 1 0 6256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_61
timestamp 1673029049
transform 1 0 6624 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1673029049
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1673029049
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1673029049
transform 1 0 1288 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1673029049
transform 1 0 2024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1673029049
transform 1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1673029049
transform 1 0 3680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_33
timestamp 1673029049
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_48
timestamp 1673029049
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_54
timestamp 1673029049
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_64
timestamp 1673029049
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1673029049
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1673029049
transform 1 0 1288 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1673029049
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1673029049
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1673029049
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_34
timestamp 1673029049
transform 1 0 4140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_46
timestamp 1673029049
transform 1 0 5244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1673029049
transform 1 0 5980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1673029049
transform 1 0 6256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_70
timestamp 1673029049
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1673029049
transform 1 0 1288 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1673029049
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1673029049
transform 1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1673029049
transform 1 0 3680 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1673029049
transform 1 0 4232 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_38
timestamp 1673029049
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_53
timestamp 1673029049
transform 1 0 5888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_70
timestamp 1673029049
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1673029049
transform 1 0 1288 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1673029049
transform 1 0 1840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_21
timestamp 1673029049
transform 1 0 2944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1673029049
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1673029049
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1673029049
transform 1 0 6072 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1673029049
transform 1 0 6256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_70
timestamp 1673029049
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1673029049
transform 1 0 1288 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_11
timestamp 1673029049
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1673029049
transform 1 0 3404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1673029049
transform 1 0 3680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_33
timestamp 1673029049
transform 1 0 4048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1673029049
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1673029049
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp 1673029049
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1673029049
transform 1 0 1288 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_18
timestamp 1673029049
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_33
timestamp 1673029049
transform 1 0 4048 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_48
timestamp 1673029049
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1673029049
transform 1 0 5980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1673029049
transform 1 0 6256 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1673029049
transform 1 0 7452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1673029049
transform 1 0 1288 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1673029049
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1673029049
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_17
timestamp 1673029049
transform 1 0 2576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_20
timestamp 1673029049
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1673029049
transform 1 0 3404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1673029049
transform 1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1673029049
transform 1 0 4140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_49
timestamp 1673029049
transform 1 0 5520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_64
timestamp 1673029049
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1673029049
transform 1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1673029049
transform 1 0 1288 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_9
timestamp 1673029049
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1673029049
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 1673029049
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1673029049
transform 1 0 5980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1673029049
transform 1 0 6256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1673029049
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1673029049
transform 1 0 1288 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1673029049
transform 1 0 2024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1673029049
transform 1 0 3404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1673029049
transform 1 0 3680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1673029049
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1673029049
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1673029049
transform 1 0 6900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_70
timestamp 1673029049
transform 1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1673029049
transform 1 0 1288 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1673029049
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1673029049
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1673029049
transform 1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp 1673029049
transform 1 0 4048 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_39
timestamp 1673029049
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1673029049
transform 1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1673029049
transform 1 0 6256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1673029049
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1673029049
transform 1 0 1012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1673029049
transform -1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1673029049
transform 1 0 1012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1673029049
transform -1 0 7912 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1673029049
transform 1 0 1012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1673029049
transform -1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1673029049
transform 1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1673029049
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1673029049
transform 1 0 1012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1673029049
transform -1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1673029049
transform 1 0 1012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1673029049
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1673029049
transform 1 0 1012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1673029049
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1673029049
transform 1 0 1012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1673029049
transform -1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1673029049
transform 1 0 1012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1673029049
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1673029049
transform 1 0 1012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1673029049
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1673029049
transform 1 0 1012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1673029049
transform -1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1673029049
transform 1 0 1012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1673029049
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1673029049
transform 1 0 1012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1673029049
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1673029049
transform 1 0 1012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1673029049
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1673029049
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1673029049
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1673029049
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1673029049
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1673029049
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1673029049
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1673029049
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1673029049
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1673029049
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1673029049
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1673029049
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1673029049
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1673029049
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1673029049
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1673029049
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1673029049
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 2576 1040 2896 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4301 1040 4621 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6026 1040 6346 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7751 1040 8071 8752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1714 1040 2034 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3439 1040 3759 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5164 1040 5484 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6889 1040 7209 8752 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 7930 9200 7986 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[0]
port 2 nsew signal input
flabel metal2 s 2410 9200 2466 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[10]
port 3 nsew signal input
flabel metal2 s 1858 9200 1914 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[11]
port 4 nsew signal input
flabel metal2 s 1306 9200 1362 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[12]
port 5 nsew signal input
flabel metal2 s 754 9200 810 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[13]
port 6 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 mgmt_gpio_in[14]
port 7 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 mgmt_gpio_in[15]
port 8 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 mgmt_gpio_in[16]
port 9 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 mgmt_gpio_in[17]
port 10 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 mgmt_gpio_in[18]
port 11 nsew signal input
flabel metal2 s 7378 9200 7434 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[1]
port 12 nsew signal input
flabel metal2 s 6826 9200 6882 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[2]
port 13 nsew signal input
flabel metal2 s 6274 9200 6330 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[3]
port 14 nsew signal input
flabel metal2 s 5722 9200 5778 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[4]
port 15 nsew signal input
flabel metal2 s 5170 9200 5226 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[5]
port 16 nsew signal input
flabel metal2 s 4618 9200 4674 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[6]
port 17 nsew signal input
flabel metal2 s 4066 9200 4122 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[7]
port 18 nsew signal input
flabel metal2 s 3514 9200 3570 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[8]
port 19 nsew signal input
flabel metal2 s 2962 9200 3018 10000 0 FreeSans 224 90 0 0 mgmt_gpio_in[9]
port 20 nsew signal input
flabel metal3 s 8200 1776 9000 1896 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[0]
port 21 nsew signal tristate
flabel metal3 s 8200 5856 9000 5976 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[10]
port 22 nsew signal tristate
flabel metal3 s 8200 6264 9000 6384 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[11]
port 23 nsew signal tristate
flabel metal3 s 8200 6672 9000 6792 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[12]
port 24 nsew signal tristate
flabel metal3 s 8200 7080 9000 7200 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[13]
port 25 nsew signal tristate
flabel metal3 s 8200 7488 9000 7608 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[14]
port 26 nsew signal tristate
flabel metal3 s 8200 7896 9000 8016 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[15]
port 27 nsew signal tristate
flabel metal3 s 8200 8304 9000 8424 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[16]
port 28 nsew signal tristate
flabel metal3 s 8200 8712 9000 8832 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[17]
port 29 nsew signal tristate
flabel metal3 s 8200 9120 9000 9240 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[18]
port 30 nsew signal tristate
flabel metal3 s 8200 2184 9000 2304 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[1]
port 31 nsew signal tristate
flabel metal3 s 8200 2592 9000 2712 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[2]
port 32 nsew signal tristate
flabel metal3 s 8200 3000 9000 3120 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[3]
port 33 nsew signal tristate
flabel metal3 s 8200 3408 9000 3528 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[4]
port 34 nsew signal tristate
flabel metal3 s 8200 3816 9000 3936 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[5]
port 35 nsew signal tristate
flabel metal3 s 8200 4224 9000 4344 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[6]
port 36 nsew signal tristate
flabel metal3 s 8200 4632 9000 4752 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[7]
port 37 nsew signal tristate
flabel metal3 s 8200 5040 9000 5160 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[8]
port 38 nsew signal tristate
flabel metal3 s 8200 5448 9000 5568 0 FreeSans 480 0 0 0 mgmt_gpio_in_buf[9]
port 39 nsew signal tristate
flabel metal3 s 8200 552 9000 672 0 FreeSans 480 0 0 0 mgmt_gpio_oeb[0]
port 40 nsew signal input
flabel metal3 s 8200 960 9000 1080 0 FreeSans 480 0 0 0 mgmt_gpio_oeb[1]
port 41 nsew signal input
flabel metal3 s 8200 1368 9000 1488 0 FreeSans 480 0 0 0 mgmt_gpio_oeb[2]
port 42 nsew signal input
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 mgmt_gpio_oeb_buf[0]
port 43 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 mgmt_gpio_oeb_buf[1]
port 44 nsew signal tristate
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 mgmt_gpio_oeb_buf[2]
port 45 nsew signal tristate
flabel metal2 s 294 0 350 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[0]
port 46 nsew signal input
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[10]
port 47 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[11]
port 48 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[12]
port 49 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[13]
port 50 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[14]
port 51 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[15]
port 52 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[16]
port 53 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[17]
port 54 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[18]
port 55 nsew signal input
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[1]
port 56 nsew signal input
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[2]
port 57 nsew signal input
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[3]
port 58 nsew signal input
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[4]
port 59 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[5]
port 60 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[6]
port 61 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[7]
port 62 nsew signal input
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[8]
port 63 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 mgmt_gpio_out[9]
port 64 nsew signal input
flabel metal2 s 8206 9200 8262 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[0]
port 65 nsew signal tristate
flabel metal2 s 2686 9200 2742 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[10]
port 66 nsew signal tristate
flabel metal2 s 2134 9200 2190 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[11]
port 67 nsew signal tristate
flabel metal2 s 1582 9200 1638 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[12]
port 68 nsew signal tristate
flabel metal2 s 1030 9200 1086 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[13]
port 69 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[14]
port 70 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[15]
port 71 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[16]
port 72 nsew signal tristate
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[17]
port 73 nsew signal tristate
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 mgmt_gpio_out_buf[18]
port 74 nsew signal tristate
flabel metal2 s 7654 9200 7710 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[1]
port 75 nsew signal tristate
flabel metal2 s 7102 9200 7158 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[2]
port 76 nsew signal tristate
flabel metal2 s 6550 9200 6606 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[3]
port 77 nsew signal tristate
flabel metal2 s 5998 9200 6054 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[4]
port 78 nsew signal tristate
flabel metal2 s 5446 9200 5502 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[5]
port 79 nsew signal tristate
flabel metal2 s 4894 9200 4950 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[6]
port 80 nsew signal tristate
flabel metal2 s 4342 9200 4398 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[7]
port 81 nsew signal tristate
flabel metal2 s 3790 9200 3846 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[8]
port 82 nsew signal tristate
flabel metal2 s 3238 9200 3294 10000 0 FreeSans 224 90 0 0 mgmt_gpio_out_buf[9]
port 83 nsew signal tristate
rlabel via1 4541 8704 4541 8704 0 VGND
rlabel metal1 4462 8160 4462 8160 0 VPWR
rlabel metal1 7544 4182 7544 4182 0 mgmt_gpio_in[0]
rlabel metal2 2346 8483 2346 8483 0 mgmt_gpio_in[10]
rlabel metal2 1886 8952 1886 8952 0 mgmt_gpio_in[11]
rlabel metal1 1518 7514 1518 7514 0 mgmt_gpio_in[12]
rlabel metal2 1518 7650 1518 7650 0 mgmt_gpio_in[13]
rlabel metal1 2254 2074 2254 2074 0 mgmt_gpio_in[14]
rlabel metal1 1840 6970 1840 6970 0 mgmt_gpio_in[15]
rlabel metal2 3266 6137 3266 6137 0 mgmt_gpio_in[16]
rlabel metal2 4186 5457 4186 5457 0 mgmt_gpio_in[17]
rlabel metal3 2438 1836 2438 1836 0 mgmt_gpio_in[18]
rlabel metal1 7452 4590 7452 4590 0 mgmt_gpio_in[1]
rlabel metal2 7406 5814 7406 5814 0 mgmt_gpio_in[2]
rlabel metal2 6486 7497 6486 7497 0 mgmt_gpio_in[3]
rlabel metal1 5612 6766 5612 6766 0 mgmt_gpio_in[4]
rlabel metal1 6716 8058 6716 8058 0 mgmt_gpio_in[5]
rlabel metal1 5474 6698 5474 6698 0 mgmt_gpio_in[6]
rlabel metal1 6026 7446 6026 7446 0 mgmt_gpio_in[7]
rlabel metal1 4094 8602 4094 8602 0 mgmt_gpio_in[8]
rlabel metal2 3910 8262 3910 8262 0 mgmt_gpio_in[9]
rlabel metal3 7460 1836 7460 1836 0 mgmt_gpio_in_buf[0]
rlabel metal1 6302 7786 6302 7786 0 mgmt_gpio_in_buf[10]
rlabel metal1 5888 8398 5888 8398 0 mgmt_gpio_in_buf[11]
rlabel metal2 4830 7259 4830 7259 0 mgmt_gpio_in_buf[12]
rlabel metal1 3726 7786 3726 7786 0 mgmt_gpio_in_buf[13]
rlabel metal1 3772 8398 3772 8398 0 mgmt_gpio_in_buf[14]
rlabel metal1 3082 7480 3082 7480 0 mgmt_gpio_in_buf[15]
rlabel metal1 5520 7378 5520 7378 0 mgmt_gpio_in_buf[16]
rlabel metal2 5290 6494 5290 6494 0 mgmt_gpio_in_buf[17]
rlabel via2 5474 5763 5474 5763 0 mgmt_gpio_in_buf[18]
rlabel metal3 8188 2312 8188 2312 0 mgmt_gpio_in_buf[1]
rlabel metal3 7452 2584 7452 2584 0 mgmt_gpio_in_buf[2]
rlabel metal1 6946 5610 6946 5610 0 mgmt_gpio_in_buf[3]
rlabel metal1 4738 6664 4738 6664 0 mgmt_gpio_in_buf[4]
rlabel metal1 6992 6222 6992 6222 0 mgmt_gpio_in_buf[5]
rlabel metal1 6624 6698 6624 6698 0 mgmt_gpio_in_buf[6]
rlabel metal2 7314 6001 7314 6001 0 mgmt_gpio_in_buf[7]
rlabel metal1 5658 7310 5658 7310 0 mgmt_gpio_in_buf[8]
rlabel metal1 7728 8398 7728 8398 0 mgmt_gpio_in_buf[9]
rlabel metal2 6762 1921 6762 1921 0 mgmt_gpio_oeb[0]
rlabel metal2 7406 1037 7406 1037 0 mgmt_gpio_oeb[1]
rlabel metal2 5934 1377 5934 1377 0 mgmt_gpio_oeb[2]
rlabel metal3 1579 4284 1579 4284 0 mgmt_gpio_oeb_buf[0]
rlabel metal3 1579 2244 1579 2244 0 mgmt_gpio_oeb_buf[1]
rlabel metal3 1602 884 1602 884 0 mgmt_gpio_oeb_buf[2]
rlabel metal1 1288 3978 1288 3978 0 mgmt_gpio_out[0]
rlabel metal2 4968 2380 4968 2380 0 mgmt_gpio_out[10]
rlabel metal2 5382 823 5382 823 0 mgmt_gpio_out[11]
rlabel metal2 1702 3298 1702 3298 0 mgmt_gpio_out[12]
rlabel metal2 6348 2380 6348 2380 0 mgmt_gpio_out[13]
rlabel metal2 6716 1428 6716 1428 0 mgmt_gpio_out[14]
rlabel metal1 3358 2380 3358 2380 0 mgmt_gpio_out[15]
rlabel metal1 5106 1258 5106 1258 0 mgmt_gpio_out[16]
rlabel metal1 5198 1938 5198 1938 0 mgmt_gpio_out[17]
rlabel metal1 3680 1938 3680 1938 0 mgmt_gpio_out[18]
rlabel via1 1334 4454 1334 4454 0 mgmt_gpio_out[1]
rlabel metal1 5842 3434 5842 3434 0 mgmt_gpio_out[2]
rlabel metal1 2990 3706 2990 3706 0 mgmt_gpio_out[3]
rlabel metal2 2162 2132 2162 2132 0 mgmt_gpio_out[4]
rlabel metal1 2346 2822 2346 2822 0 mgmt_gpio_out[5]
rlabel metal1 3910 2312 3910 2312 0 mgmt_gpio_out[6]
rlabel metal2 3772 748 3772 748 0 mgmt_gpio_out[7]
rlabel metal2 4002 6460 4002 6460 0 mgmt_gpio_out[8]
rlabel metal2 4278 748 4278 748 0 mgmt_gpio_out[9]
rlabel metal1 5290 4114 5290 4114 0 mgmt_gpio_out_buf[0]
rlabel metal2 2615 9316 2615 9316 0 mgmt_gpio_out_buf[10]
rlabel metal2 2162 7422 2162 7422 0 mgmt_gpio_out_buf[11]
rlabel metal2 1511 9316 1511 9316 0 mgmt_gpio_out_buf[12]
rlabel metal1 1426 6358 1426 6358 0 mgmt_gpio_out_buf[13]
rlabel metal2 3358 6035 3358 6035 0 mgmt_gpio_out_buf[14]
rlabel metal3 958 7684 958 7684 0 mgmt_gpio_out_buf[15]
rlabel metal1 4416 1394 4416 1394 0 mgmt_gpio_out_buf[16]
rlabel metal3 1142 4964 1142 4964 0 mgmt_gpio_out_buf[17]
rlabel metal1 2898 2006 2898 2006 0 mgmt_gpio_out_buf[18]
rlabel metal1 4094 5304 4094 5304 0 mgmt_gpio_out_buf[1]
rlabel metal1 6670 4658 6670 4658 0 mgmt_gpio_out_buf[2]
rlabel metal1 5566 5270 5566 5270 0 mgmt_gpio_out_buf[3]
rlabel metal1 5566 3570 5566 3570 0 mgmt_gpio_out_buf[4]
rlabel metal1 5060 3094 5060 3094 0 mgmt_gpio_out_buf[5]
rlabel metal1 4830 2482 4830 2482 0 mgmt_gpio_out_buf[6]
rlabel metal1 3680 5746 3680 5746 0 mgmt_gpio_out_buf[7]
rlabel metal1 3542 6358 3542 6358 0 mgmt_gpio_out_buf[8]
rlabel metal2 3174 7293 3174 7293 0 mgmt_gpio_out_buf[9]
<< properties >>
string FIXED_BBOX 0 0 9000 10000
<< end >>
