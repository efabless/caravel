magic
tech sky130A
magscale 1 2
timestamp 1663176679
<< viali >>
rect 3801 11305 3835 11339
rect 8033 11305 8067 11339
rect 9229 11305 9263 11339
rect 6193 11237 6227 11271
rect 6653 11237 6687 11271
rect 8309 11169 8343 11203
rect 8493 11169 8527 11203
rect 9413 11169 9447 11203
rect 3065 11101 3099 11135
rect 4077 11101 4111 11135
rect 4353 11101 4387 11135
rect 5181 11101 5215 11135
rect 6009 11101 6043 11135
rect 7941 11101 7975 11135
rect 8861 11101 8895 11135
rect 3433 11033 3467 11067
rect 3709 11033 3743 11067
rect 4261 11033 4295 11067
rect 4905 11033 4939 11067
rect 2973 10965 3007 10999
rect 4629 10965 4663 10999
rect 5917 10965 5951 10999
rect 6469 10965 6503 10999
rect 6929 10965 6963 10999
rect 7297 10965 7331 10999
rect 7573 10965 7607 10999
rect 7849 10965 7883 10999
rect 9045 10965 9079 10999
rect 7941 10693 7975 10727
rect 2789 10625 2823 10659
rect 4629 10625 4663 10659
rect 5365 10625 5399 10659
rect 5549 10625 5583 10659
rect 5825 10625 5859 10659
rect 6285 10625 6319 10659
rect 6561 10625 6595 10659
rect 6837 10625 6871 10659
rect 7021 10625 7055 10659
rect 7481 10625 7515 10659
rect 7665 10625 7699 10659
rect 2053 10557 2087 10591
rect 3157 10557 3191 10591
rect 2697 10421 2731 10455
rect 5189 10421 5223 10455
rect 5641 10421 5675 10455
rect 5917 10421 5951 10455
rect 6377 10421 6411 10455
rect 7113 10421 7147 10455
rect 7389 10421 7423 10455
rect 9413 10421 9447 10455
rect 4721 10217 4755 10251
rect 5365 10217 5399 10251
rect 1869 10081 1903 10115
rect 3341 10081 3375 10115
rect 4169 10081 4203 10115
rect 4813 10081 4847 10115
rect 5457 10081 5491 10115
rect 1593 10013 1627 10047
rect 4537 10013 4571 10047
rect 5089 10013 5123 10047
rect 5825 10013 5859 10047
rect 7297 10013 7331 10047
rect 8125 10013 8159 10047
rect 8493 10013 8527 10047
rect 9137 10013 9171 10047
rect 8309 9945 8343 9979
rect 8769 9945 8803 9979
rect 8953 9945 8987 9979
rect 3617 9877 3651 9911
rect 4445 9877 4479 9911
rect 7861 9877 7895 9911
rect 9321 9877 9355 9911
rect 9413 9877 9447 9911
rect 6193 9673 6227 9707
rect 6009 9605 6043 9639
rect 3249 9537 3283 9571
rect 3341 9537 3375 9571
rect 5181 9537 5215 9571
rect 7021 9537 7055 9571
rect 8861 9537 8895 9571
rect 1501 9469 1535 9503
rect 2973 9469 3007 9503
rect 3709 9469 3743 9503
rect 6745 9469 6779 9503
rect 7389 9469 7423 9503
rect 5745 9401 5779 9435
rect 9421 9333 9455 9367
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 4077 9129 4111 9163
rect 4629 9129 4663 9163
rect 8217 9129 8251 9163
rect 9505 9129 9539 9163
rect 3433 9061 3467 9095
rect 8493 9061 8527 9095
rect 6377 8993 6411 9027
rect 6469 8993 6503 9027
rect 2605 8925 2639 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 3801 8925 3835 8959
rect 3985 8925 4019 8959
rect 8861 8925 8895 8959
rect 3065 8857 3099 8891
rect 3709 8857 3743 8891
rect 6101 8857 6135 8891
rect 6745 8857 6779 8891
rect 4353 8789 4387 8823
rect 9045 8789 9079 8823
rect 9321 8789 9355 8823
rect 4721 8585 4755 8619
rect 7481 8585 7515 8619
rect 8033 8585 8067 8619
rect 1777 8517 1811 8551
rect 6193 8517 6227 8551
rect 9137 8517 9171 8551
rect 1501 8449 1535 8483
rect 6009 8449 6043 8483
rect 8585 8449 8619 8483
rect 8953 8449 8987 8483
rect 9229 8449 9263 8483
rect 3249 8381 3283 8415
rect 3985 8381 4019 8415
rect 8769 8313 8803 8347
rect 9413 8313 9447 8347
rect 3433 8245 3467 8279
rect 2789 8041 2823 8075
rect 3433 8041 3467 8075
rect 9413 8041 9447 8075
rect 4721 7973 4755 8007
rect 9045 7973 9079 8007
rect 6101 7905 6135 7939
rect 9321 7905 9355 7939
rect 3065 7837 3099 7871
rect 3617 7837 3651 7871
rect 4077 7837 4111 7871
rect 6469 7837 6503 7871
rect 7941 7837 7975 7871
rect 3249 7769 3283 7803
rect 3893 7769 3927 7803
rect 6009 7769 6043 7803
rect 8505 7769 8539 7803
rect 2973 7701 3007 7735
rect 8861 7701 8895 7735
rect 2513 7497 2547 7531
rect 9413 7497 9447 7531
rect 7941 7429 7975 7463
rect 9045 7429 9079 7463
rect 2789 7361 2823 7395
rect 3157 7361 3191 7395
rect 4629 7361 4663 7395
rect 5549 7361 5583 7395
rect 6009 7361 6043 7395
rect 9229 7361 9263 7395
rect 6193 7293 6227 7327
rect 8585 7293 8619 7327
rect 8953 7293 8987 7327
rect 5193 7225 5227 7259
rect 2697 7157 2731 7191
rect 5917 7157 5951 7191
rect 8033 7157 8067 7191
rect 1764 6953 1798 6987
rect 1501 6817 1535 6851
rect 3249 6817 3283 6851
rect 4169 6817 4203 6851
rect 8401 6817 8435 6851
rect 8953 6817 8987 6851
rect 4353 6749 4387 6783
rect 4813 6749 4847 6783
rect 5089 6749 5123 6783
rect 5457 6749 5491 6783
rect 6929 6749 6963 6783
rect 7849 6749 7883 6783
rect 8125 6749 8159 6783
rect 4629 6681 4663 6715
rect 7757 6681 7791 6715
rect 8309 6681 8343 6715
rect 9137 6681 9171 6715
rect 3617 6613 3651 6647
rect 7493 6613 7527 6647
rect 9045 6613 9079 6647
rect 9505 6613 9539 6647
rect 2237 6409 2271 6443
rect 8125 6409 8159 6443
rect 8953 6409 8987 6443
rect 9045 6409 9079 6443
rect 9505 6409 9539 6443
rect 2053 6341 2087 6375
rect 2421 6341 2455 6375
rect 8309 6341 8343 6375
rect 8769 6341 8803 6375
rect 9137 6341 9171 6375
rect 2697 6273 2731 6307
rect 3157 6273 3191 6307
rect 4629 6273 4663 6307
rect 5365 6273 5399 6307
rect 6193 6273 6227 6307
rect 8493 6273 8527 6307
rect 8677 6273 8711 6307
rect 2605 6205 2639 6239
rect 2789 6205 2823 6239
rect 5917 6205 5951 6239
rect 6469 6205 6503 6239
rect 7941 6205 7975 6239
rect 9321 6137 9355 6171
rect 5193 6069 5227 6103
rect 1501 5865 1535 5899
rect 1856 5865 1890 5899
rect 3985 5865 4019 5899
rect 5917 5865 5951 5899
rect 8217 5865 8251 5899
rect 8585 5865 8619 5899
rect 8401 5797 8435 5831
rect 1593 5729 1627 5763
rect 4445 5729 4479 5763
rect 6193 5729 6227 5763
rect 6469 5729 6503 5763
rect 7941 5729 7975 5763
rect 4169 5661 4203 5695
rect 3709 5593 3743 5627
rect 3893 5593 3927 5627
rect 8861 5593 8895 5627
rect 8953 5593 8987 5627
rect 9505 5593 9539 5627
rect 3341 5525 3375 5559
rect 5273 5321 5307 5355
rect 8309 5321 8343 5355
rect 3617 5253 3651 5287
rect 8125 5253 8159 5287
rect 9045 5253 9079 5287
rect 3341 5185 3375 5219
rect 6009 5185 6043 5219
rect 9229 5185 9263 5219
rect 5825 5117 5859 5151
rect 6285 5117 6319 5151
rect 7757 5117 7791 5151
rect 8861 5117 8895 5151
rect 5089 4981 5123 5015
rect 9321 4981 9355 5015
rect 5733 4777 5767 4811
rect 9413 4777 9447 4811
rect 3341 4641 3375 4675
rect 5365 4641 5399 4675
rect 6285 4641 6319 4675
rect 5457 4573 5491 4607
rect 6561 4573 6595 4607
rect 6929 4573 6963 4607
rect 8401 4573 8435 4607
rect 9321 4573 9355 4607
rect 3617 4505 3651 4539
rect 5089 4437 5123 4471
rect 8961 4437 8995 4471
rect 9229 4437 9263 4471
rect 6377 4233 6411 4267
rect 9045 4233 9079 4267
rect 9229 4233 9263 4267
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 5365 4097 5399 4131
rect 6285 4097 6319 4131
rect 8125 4097 8159 4131
rect 9505 4097 9539 4131
rect 3893 4029 3927 4063
rect 6561 4029 6595 4063
rect 8309 4029 8343 4063
rect 8861 4029 8895 4063
rect 8033 3961 8067 3995
rect 5925 3893 5959 3927
rect 6193 3893 6227 3927
rect 5457 3689 5491 3723
rect 5825 3689 5859 3723
rect 9413 3689 9447 3723
rect 3433 3553 3467 3587
rect 7205 3553 7239 3587
rect 5089 3485 5123 3519
rect 5733 3485 5767 3519
rect 6193 3485 6227 3519
rect 6745 3485 6779 3519
rect 6837 3485 6871 3519
rect 8677 3485 8711 3519
rect 5181 3417 5215 3451
rect 5365 3417 5399 3451
rect 6377 3417 6411 3451
rect 6561 3417 6595 3451
rect 9241 3417 9275 3451
rect 8861 3349 8895 3383
rect 4169 3145 4203 3179
rect 7941 3145 7975 3179
rect 8493 3145 8527 3179
rect 8953 3145 8987 3179
rect 9413 3145 9447 3179
rect 3433 3077 3467 3111
rect 7481 3077 7515 3111
rect 8125 3077 8159 3111
rect 8309 3077 8343 3111
rect 4445 3009 4479 3043
rect 6469 3009 6503 3043
rect 7267 3009 7301 3043
rect 7757 3009 7791 3043
rect 9045 3009 9079 3043
rect 3617 2941 3651 2975
rect 4629 2941 4663 2975
rect 4997 2941 5031 2975
rect 8861 2941 8895 2975
rect 7033 2873 7067 2907
rect 4353 2805 4387 2839
rect 4813 2601 4847 2635
rect 6101 2601 6135 2635
rect 6653 2601 6687 2635
rect 7021 2601 7055 2635
rect 7297 2601 7331 2635
rect 7941 2601 7975 2635
rect 9045 2601 9079 2635
rect 9229 2601 9263 2635
rect 5089 2533 5123 2567
rect 6469 2533 6503 2567
rect 6837 2533 6871 2567
rect 8493 2533 8527 2567
rect 9413 2533 9447 2567
rect 3433 2465 3467 2499
rect 5365 2465 5399 2499
rect 5549 2465 5583 2499
rect 3617 2397 3651 2431
rect 3985 2397 4019 2431
rect 4169 2397 4203 2431
rect 4353 2397 4387 2431
rect 4905 2397 4939 2431
rect 5917 2397 5951 2431
rect 6193 2397 6227 2431
rect 6929 2397 6963 2431
rect 7573 2397 7607 2431
rect 7849 2397 7883 2431
rect 8125 2397 8159 2431
rect 8677 2397 8711 2431
rect 3801 2329 3835 2363
rect 4537 2329 4571 2363
rect 8309 2329 8343 2363
rect 9091 2329 9125 2363
rect 5745 2057 5779 2091
rect 8309 2057 8343 2091
rect 8585 2057 8619 2091
rect 8769 2057 8803 2091
rect 9321 2057 9355 2091
rect 6009 1989 6043 2023
rect 7297 1989 7331 2023
rect 7941 1989 7975 2023
rect 9413 1989 9447 2023
rect 3341 1921 3375 1955
rect 5181 1921 5215 1955
rect 3709 1853 3743 1887
rect 9137 1853 9171 1887
rect 8953 1717 8987 1751
rect 5365 1513 5399 1547
rect 9505 1513 9539 1547
rect 5273 1445 5307 1479
rect 5089 1309 5123 1343
rect 3801 1173 3835 1207
<< obsli1 >>
rect 0 12986 853 13014
rect 0 12969 9963 12986
rect 0 11481 33962 12969
rect 0 6005 853 11481
rect 0 5899 3359 6005
rect 0 5865 1501 5899
rect 1535 5865 1856 5899
rect 1890 5865 3359 5899
rect 0 5763 3359 5865
rect 0 5729 1593 5763
rect 1627 5729 3359 5763
rect 0 5559 3359 5729
rect 0 5525 3341 5559
rect 0 5219 3359 5525
rect 0 5185 3341 5219
rect 0 4675 3359 5185
rect 0 4641 3341 4675
rect 0 4131 3359 4641
rect 0 4097 3341 4131
rect 0 1955 3359 4097
rect 0 1921 3341 1955
rect 0 0 3359 1921
rect 9800 1048 33962 11481
rect 3366 0 33962 1048
<< metal1 >>
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 1820 11308 3801 11336
rect 1820 11296 1826 11308
rect 3789 11305 3801 11308
rect 3835 11336 3847 11339
rect 4338 11336 4344 11348
rect 3835 11308 4344 11336
rect 3835 11305 3847 11308
rect 3789 11299 3847 11305
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 6512 11308 8033 11336
rect 6512 11296 6518 11308
rect 8021 11305 8033 11308
rect 8067 11336 8079 11339
rect 8110 11336 8116 11348
rect 8067 11308 8116 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8110 11296 8116 11308
rect 8168 11336 8174 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 8168 11308 9229 11336
rect 8168 11296 8174 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 1210 11228 1216 11280
rect 1268 11268 1274 11280
rect 6181 11271 6239 11277
rect 6181 11268 6193 11271
rect 1268 11240 6193 11268
rect 1268 11228 1274 11240
rect 6181 11237 6193 11240
rect 6227 11268 6239 11271
rect 6546 11268 6552 11280
rect 6227 11240 6552 11268
rect 6227 11237 6239 11240
rect 6181 11231 6239 11237
rect 6546 11228 6552 11240
rect 6604 11268 6610 11280
rect 6641 11271 6699 11277
rect 6641 11268 6653 11271
rect 6604 11240 6653 11268
rect 6604 11228 6610 11240
rect 6641 11237 6653 11240
rect 6687 11237 6699 11271
rect 6641 11231 6699 11237
rect 4706 11200 4712 11212
rect 3068 11172 4712 11200
rect 3068 11141 3096 11172
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 6270 11200 6276 11212
rect 5592 11172 6276 11200
rect 5592 11160 5598 11172
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 7340 11172 8309 11200
rect 7340 11160 7346 11172
rect 8297 11169 8309 11172
rect 8343 11200 8355 11203
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 8343 11172 8493 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 8481 11169 8493 11172
rect 8527 11200 8539 11203
rect 9401 11203 9459 11209
rect 9401 11200 9413 11203
rect 8527 11172 9413 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 9401 11169 9413 11172
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4338 11132 4344 11144
rect 4299 11104 4344 11132
rect 4065 11095 4123 11101
rect 3421 11067 3479 11073
rect 3421 11033 3433 11067
rect 3467 11064 3479 11067
rect 3697 11067 3755 11073
rect 3697 11064 3709 11067
rect 3467 11036 3709 11064
rect 3467 11033 3479 11036
rect 3421 11027 3479 11033
rect 3697 11033 3709 11036
rect 3743 11033 3755 11067
rect 3697 11027 3755 11033
rect 2958 10996 2964 11008
rect 2919 10968 2964 10996
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 3712 10996 3740 11027
rect 4080 10996 4108 11095
rect 4338 11092 4344 11104
rect 4396 11132 4402 11144
rect 4982 11132 4988 11144
rect 4396 11104 4988 11132
rect 4396 11092 4402 11104
rect 4982 11092 4988 11104
rect 5040 11132 5046 11144
rect 5169 11135 5227 11141
rect 5169 11132 5181 11135
rect 5040 11104 5181 11132
rect 5040 11092 5046 11104
rect 5169 11101 5181 11104
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 4246 11064 4252 11076
rect 4207 11036 4252 11064
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 4893 11067 4951 11073
rect 4893 11064 4905 11067
rect 4448 11036 4905 11064
rect 4448 10996 4476 11036
rect 4893 11033 4905 11036
rect 4939 11064 4951 11067
rect 5626 11064 5632 11076
rect 4939 11036 5632 11064
rect 4939 11033 4951 11036
rect 4893 11027 4951 11033
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 6012 11064 6040 11095
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 6880 11104 7941 11132
rect 6880 11092 6886 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11101 8907 11135
rect 8849 11095 8907 11101
rect 7466 11064 7472 11076
rect 6012 11036 7472 11064
rect 7466 11024 7472 11036
rect 7524 11064 7530 11076
rect 8864 11064 8892 11095
rect 16574 11064 16580 11076
rect 7524 11036 8892 11064
rect 9048 11036 16580 11064
rect 7524 11024 7530 11036
rect 4614 10996 4620 11008
rect 3712 10968 4476 10996
rect 4575 10968 4620 10996
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 5905 10999 5963 11005
rect 5905 10996 5917 10999
rect 5592 10968 5917 10996
rect 5592 10956 5598 10968
rect 5905 10965 5917 10968
rect 5951 10965 5963 10999
rect 5905 10959 5963 10965
rect 6457 10999 6515 11005
rect 6457 10965 6469 10999
rect 6503 10996 6515 10999
rect 6917 10999 6975 11005
rect 6917 10996 6929 10999
rect 6503 10968 6929 10996
rect 6503 10965 6515 10968
rect 6457 10959 6515 10965
rect 6917 10965 6929 10968
rect 6963 10996 6975 10999
rect 7282 10996 7288 11008
rect 6963 10968 7288 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 7282 10956 7288 10968
rect 7340 10996 7346 11008
rect 7561 10999 7619 11005
rect 7561 10996 7573 10999
rect 7340 10968 7573 10996
rect 7340 10956 7346 10968
rect 7561 10965 7573 10968
rect 7607 10965 7619 10999
rect 7561 10959 7619 10965
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 9048 11005 9076 11036
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 7708 10968 7849 10996
rect 7708 10956 7714 10968
rect 7837 10965 7849 10968
rect 7883 10965 7895 10999
rect 7837 10959 7895 10965
rect 9033 10999 9091 11005
rect 9033 10965 9045 10999
rect 9079 10965 9091 10999
rect 9033 10959 9091 10965
rect 920 10906 9844 10928
rect 920 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 5194 10906
rect 5246 10854 5258 10906
rect 5310 10854 5322 10906
rect 5374 10854 9844 10906
rect 920 10832 9844 10854
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6454 10792 6460 10804
rect 6052 10764 6460 10792
rect 6052 10752 6058 10764
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 4522 10724 4528 10736
rect 4278 10696 4528 10724
rect 4522 10684 4528 10696
rect 4580 10684 4586 10736
rect 4706 10684 4712 10736
rect 4764 10724 4770 10736
rect 7929 10727 7987 10733
rect 4764 10696 7512 10724
rect 4764 10684 4770 10696
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 2958 10656 2964 10668
rect 2823 10628 2964 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4617 10659 4675 10665
rect 4617 10656 4629 10659
rect 4396 10628 4629 10656
rect 4396 10616 4402 10628
rect 4617 10625 4629 10628
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5828 10665 5856 10696
rect 7484 10668 7512 10696
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 8202 10724 8208 10736
rect 7975 10696 8208 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5040 10628 5365 10656
rect 5040 10616 5046 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 6273 10659 6331 10665
rect 6273 10625 6285 10659
rect 6319 10625 6331 10659
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 6273 10619 6331 10625
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 2041 10591 2099 10597
rect 2041 10588 2053 10591
rect 1636 10560 2053 10588
rect 1636 10548 1642 10560
rect 2041 10557 2053 10560
rect 2087 10557 2099 10591
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 2041 10551 2099 10557
rect 2700 10560 3157 10588
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 2700 10461 2728 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 5552 10588 5580 10619
rect 5626 10588 5632 10600
rect 5539 10560 5632 10588
rect 3145 10551 3203 10557
rect 5626 10548 5632 10560
rect 5684 10588 5690 10600
rect 6288 10588 6316 10619
rect 6546 10616 6552 10628
rect 6604 10656 6610 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6604 10628 6837 10656
rect 6604 10616 6610 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 7009 10619 7067 10625
rect 7024 10588 7052 10619
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7650 10656 7656 10668
rect 7611 10628 7656 10656
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 9398 10656 9404 10668
rect 9062 10642 9404 10656
rect 9048 10628 9404 10642
rect 7282 10588 7288 10600
rect 5684 10560 7288 10588
rect 5684 10548 5690 10560
rect 6288 10520 6316 10560
rect 7282 10548 7288 10560
rect 7340 10588 7346 10600
rect 9048 10588 9076 10628
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 7340 10560 9076 10588
rect 7340 10548 7346 10560
rect 6104 10492 6316 10520
rect 2685 10455 2743 10461
rect 2685 10452 2697 10455
rect 1820 10424 2697 10452
rect 1820 10412 1826 10424
rect 2685 10421 2697 10424
rect 2731 10421 2743 10455
rect 2685 10415 2743 10421
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 5177 10455 5235 10461
rect 5177 10452 5189 10455
rect 4948 10424 5189 10452
rect 4948 10412 4954 10424
rect 5177 10421 5189 10424
rect 5223 10421 5235 10455
rect 5626 10452 5632 10464
rect 5587 10424 5632 10452
rect 5177 10415 5235 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5902 10452 5908 10464
rect 5863 10424 5908 10452
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6104 10452 6132 10492
rect 6362 10452 6368 10464
rect 6052 10424 6132 10452
rect 6323 10424 6368 10452
rect 6052 10412 6058 10424
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 7098 10452 7104 10464
rect 7059 10424 7104 10452
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 7377 10455 7435 10461
rect 7377 10452 7389 10455
rect 7248 10424 7389 10452
rect 7248 10412 7254 10424
rect 7377 10421 7389 10424
rect 7423 10421 7435 10455
rect 7377 10415 7435 10421
rect 9401 10455 9459 10461
rect 9401 10421 9413 10455
rect 9447 10452 9459 10455
rect 16574 10452 16580 10464
rect 9447 10424 16580 10452
rect 9447 10421 9459 10424
rect 9401 10415 9459 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 4522 10208 4528 10260
rect 4580 10248 4586 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 4580 10220 4721 10248
rect 4580 10208 4586 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 5353 10251 5411 10257
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 5994 10248 6000 10260
rect 5399 10220 6000 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 3329 10115 3387 10121
rect 1903 10084 3280 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 1486 10004 1492 10056
rect 1544 10044 1550 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 1544 10016 1593 10044
rect 1544 10004 1550 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 2314 9936 2320 9988
rect 2372 9936 2378 9988
rect 3252 9976 3280 10084
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 4157 10115 4215 10121
rect 4157 10112 4169 10115
rect 3375 10084 4169 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 4157 10081 4169 10084
rect 4203 10081 4215 10115
rect 4157 10075 4215 10081
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 4672 10084 4813 10112
rect 4672 10072 4678 10084
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 5368 10112 5396 10211
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 4801 10075 4859 10081
rect 5092 10084 5396 10112
rect 5445 10115 5503 10121
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 4706 10044 4712 10056
rect 4571 10016 4712 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 5092 10053 5120 10084
rect 5445 10081 5457 10115
rect 5491 10112 5503 10115
rect 5534 10112 5540 10124
rect 5491 10084 5540 10112
rect 5491 10081 5503 10084
rect 5445 10075 5503 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 8128 10084 9168 10112
rect 8128 10056 8156 10084
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5810 10044 5816 10056
rect 5077 10007 5135 10013
rect 5184 10016 5816 10044
rect 5184 9976 5212 10016
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 7285 10047 7343 10053
rect 7285 10044 7297 10047
rect 7156 10016 7297 10044
rect 7156 10004 7162 10016
rect 7285 10013 7297 10016
rect 7331 10013 7343 10047
rect 8110 10044 8116 10056
rect 8071 10016 8116 10044
rect 7285 10007 7343 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 9140 10053 9168 10084
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10044 8539 10047
rect 9125 10047 9183 10053
rect 8527 10016 8984 10044
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 3252 9948 5212 9976
rect 6362 9936 6368 9988
rect 6420 9936 6426 9988
rect 8294 9976 8300 9988
rect 8255 9948 8300 9976
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 8757 9979 8815 9985
rect 8757 9945 8769 9979
rect 8803 9976 8815 9979
rect 8846 9976 8852 9988
rect 8803 9948 8852 9976
rect 8803 9945 8815 9948
rect 8757 9939 8815 9945
rect 8846 9936 8852 9948
rect 8904 9936 8910 9988
rect 8956 9985 8984 10016
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 8941 9979 8999 9985
rect 8941 9945 8953 9979
rect 8987 9976 8999 9979
rect 8987 9948 9352 9976
rect 8987 9945 8999 9948
rect 8941 9939 8999 9945
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9908 3663 9911
rect 3694 9908 3700 9920
rect 3651 9880 3700 9908
rect 3651 9877 3663 9880
rect 3605 9871 3663 9877
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4433 9911 4491 9917
rect 4433 9908 4445 9911
rect 4212 9880 4445 9908
rect 4212 9868 4218 9880
rect 4433 9877 4445 9880
rect 4479 9877 4491 9911
rect 4433 9871 4491 9877
rect 7849 9911 7907 9917
rect 7849 9877 7861 9911
rect 7895 9908 7907 9911
rect 9122 9908 9128 9920
rect 7895 9880 9128 9908
rect 7895 9877 7907 9880
rect 7849 9871 7907 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9324 9917 9352 9948
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9398 9908 9404 9920
rect 9355 9880 9404 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 920 9818 9844 9840
rect 920 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 5194 9818
rect 5246 9766 5258 9818
rect 5310 9766 5322 9818
rect 5374 9766 9844 9818
rect 920 9744 9844 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 1544 9676 2728 9704
rect 1544 9664 1550 9676
rect 2314 9596 2320 9648
rect 2372 9596 2378 9648
rect 2700 9636 2728 9676
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4890 9704 4896 9716
rect 4580 9676 4896 9704
rect 4580 9664 4586 9676
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 6181 9707 6239 9713
rect 6181 9704 6193 9707
rect 5868 9676 6193 9704
rect 5868 9664 5874 9676
rect 6181 9673 6193 9676
rect 6227 9673 6239 9707
rect 6181 9667 6239 9673
rect 2700 9608 3280 9636
rect 3252 9577 3280 9608
rect 4246 9596 4252 9648
rect 4304 9596 4310 9648
rect 5994 9636 6000 9648
rect 5955 9608 6000 9636
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 8294 9596 8300 9648
rect 8352 9596 8358 9648
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9568 3387 9571
rect 5169 9571 5227 9577
rect 3375 9540 3832 9568
rect 3375 9537 3387 9540
rect 3329 9531 3387 9537
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9500 1547 9503
rect 1578 9500 1584 9512
rect 1535 9472 1584 9500
rect 1535 9469 1547 9472
rect 1489 9463 1547 9469
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9500 3019 9503
rect 3694 9500 3700 9512
rect 3007 9472 3700 9500
rect 3007 9469 3019 9472
rect 2961 9463 3019 9469
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 3804 9500 3832 9540
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5626 9568 5632 9580
rect 5215 9540 5632 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9568 7067 9571
rect 7190 9568 7196 9580
rect 7055 9540 7196 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 8846 9568 8852 9580
rect 8807 9540 8852 9568
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 4154 9500 4160 9512
rect 3804 9472 4160 9500
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 6730 9500 6736 9512
rect 6691 9472 6736 9500
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 8018 9500 8024 9512
rect 7423 9472 8024 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 5733 9435 5791 9441
rect 5733 9401 5745 9435
rect 5779 9432 5791 9435
rect 5779 9404 7144 9432
rect 5779 9401 5791 9404
rect 5733 9395 5791 9401
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 6638 9364 6644 9376
rect 4488 9336 6644 9364
rect 4488 9324 4494 9336
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7116 9364 7144 9404
rect 8386 9364 8392 9376
rect 7116 9336 8392 9364
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 9409 9367 9467 9373
rect 9409 9364 9421 9367
rect 8720 9336 9421 9364
rect 8720 9324 8726 9336
rect 9409 9333 9421 9336
rect 9455 9333 9467 9367
rect 9409 9327 9467 9333
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2004 9132 2329 9160
rect 2004 9120 2010 9132
rect 2317 9129 2329 9132
rect 2363 9129 2375 9163
rect 2317 9123 2375 9129
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2464 9132 2789 9160
rect 2464 9120 2470 9132
rect 2777 9129 2789 9132
rect 2823 9160 2835 9163
rect 2958 9160 2964 9172
rect 2823 9132 2964 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 2958 9120 2964 9132
rect 3016 9160 3022 9172
rect 3602 9160 3608 9172
rect 3016 9132 3608 9160
rect 3016 9120 3022 9132
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 4065 9163 4123 9169
rect 4065 9129 4077 9163
rect 4111 9160 4123 9163
rect 4154 9160 4160 9172
rect 4111 9132 4160 9160
rect 4111 9129 4123 9132
rect 4065 9123 4123 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4617 9163 4675 9169
rect 4617 9129 4629 9163
rect 4663 9160 4675 9163
rect 6730 9160 6736 9172
rect 4663 9132 6736 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 8202 9160 8208 9172
rect 8163 9132 8208 9160
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 9490 9160 9496 9172
rect 9451 9132 9496 9160
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 3421 9095 3479 9101
rect 3421 9061 3433 9095
rect 3467 9092 3479 9095
rect 4338 9092 4344 9104
rect 3467 9064 4344 9092
rect 3467 9061 3479 9064
rect 3421 9055 3479 9061
rect 4338 9052 4344 9064
rect 4396 9052 4402 9104
rect 8481 9095 8539 9101
rect 8481 9061 8493 9095
rect 8527 9092 8539 9095
rect 8527 9064 16574 9092
rect 8527 9061 8539 9064
rect 8481 9055 8539 9061
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 9024 6423 9027
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 6411 8996 6469 9024
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 6457 8993 6469 8996
rect 6503 9024 6515 9027
rect 6822 9024 6828 9036
rect 6503 8996 6828 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 6822 8984 6828 8996
rect 6880 9024 6886 9036
rect 6880 8996 8892 9024
rect 6880 8984 6886 8996
rect 2314 8916 2320 8968
rect 2372 8956 2378 8968
rect 2593 8959 2651 8965
rect 2593 8956 2605 8959
rect 2372 8928 2605 8956
rect 2372 8916 2378 8928
rect 2593 8925 2605 8928
rect 2639 8956 2651 8959
rect 2866 8956 2872 8968
rect 2639 8928 2872 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2866 8916 2872 8928
rect 2924 8956 2930 8968
rect 2961 8959 3019 8965
rect 2961 8956 2973 8959
rect 2924 8928 2973 8956
rect 2924 8916 2930 8928
rect 2961 8925 2973 8928
rect 3007 8956 3019 8959
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3007 8928 3249 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3053 8891 3111 8897
rect 3053 8857 3065 8891
rect 3099 8888 3111 8891
rect 3142 8888 3148 8900
rect 3099 8860 3148 8888
rect 3099 8857 3111 8860
rect 3053 8851 3111 8857
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 3252 8888 3280 8919
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 8864 8965 8892 8996
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3660 8928 3801 8956
rect 3660 8916 3666 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8956 4031 8959
rect 8849 8959 8907 8965
rect 4019 8928 4384 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 3697 8891 3755 8897
rect 3697 8888 3709 8891
rect 3252 8860 3709 8888
rect 3697 8857 3709 8860
rect 3743 8888 3755 8891
rect 3988 8888 4016 8919
rect 3743 8860 4016 8888
rect 3743 8857 3755 8860
rect 3697 8851 3755 8857
rect 4356 8829 4384 8928
rect 8849 8925 8861 8959
rect 8895 8925 8907 8959
rect 8849 8919 8907 8925
rect 5626 8848 5632 8900
rect 5684 8888 5690 8900
rect 5994 8888 6000 8900
rect 5684 8860 6000 8888
rect 5684 8848 5690 8860
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8820 4399 8823
rect 5736 8820 5764 8860
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 6089 8891 6147 8897
rect 6089 8857 6101 8891
rect 6135 8857 6147 8891
rect 6089 8851 6147 8857
rect 6733 8891 6791 8897
rect 6733 8857 6745 8891
rect 6779 8888 6791 8891
rect 7006 8888 7012 8900
rect 6779 8860 7012 8888
rect 6779 8857 6791 8860
rect 6733 8851 6791 8857
rect 4387 8792 5764 8820
rect 6104 8820 6132 8851
rect 7006 8848 7012 8860
rect 7064 8848 7070 8900
rect 8754 8888 8760 8900
rect 7958 8860 8760 8888
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 8956 8820 8984 9064
rect 16546 9024 16574 9064
rect 16758 9024 16764 9036
rect 16546 8996 16764 9024
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 9048 8860 16574 8888
rect 9048 8829 9076 8860
rect 16546 8832 16574 8860
rect 6104 8792 8984 8820
rect 9033 8823 9091 8829
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 9033 8789 9045 8823
rect 9079 8789 9091 8823
rect 9306 8820 9312 8832
rect 9267 8792 9312 8820
rect 9033 8783 9091 8789
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 16546 8792 16580 8832
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 920 8730 9844 8752
rect 920 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 5194 8730
rect 5246 8678 5258 8730
rect 5310 8678 5322 8730
rect 5374 8678 9844 8730
rect 920 8656 9844 8678
rect 4706 8616 4712 8628
rect 4667 8588 4712 8616
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 5442 8576 5448 8628
rect 5500 8616 5506 8628
rect 5500 8588 6776 8616
rect 5500 8576 5506 8588
rect 1762 8548 1768 8560
rect 1723 8520 1768 8548
rect 1762 8508 1768 8520
rect 1820 8508 1826 8560
rect 4798 8508 4804 8560
rect 4856 8548 4862 8560
rect 6181 8551 6239 8557
rect 6181 8548 6193 8551
rect 4856 8520 6193 8548
rect 4856 8508 4862 8520
rect 6181 8517 6193 8520
rect 6227 8517 6239 8551
rect 6748 8548 6776 8588
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 6880 8588 7481 8616
rect 6880 8576 6886 8588
rect 7469 8585 7481 8588
rect 7515 8585 7527 8619
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 7469 8579 7527 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 9125 8551 9183 8557
rect 9125 8548 9137 8551
rect 6748 8520 9137 8548
rect 6181 8511 6239 8517
rect 9125 8517 9137 8520
rect 9171 8548 9183 8551
rect 9306 8548 9312 8560
rect 9171 8520 9312 8548
rect 9171 8517 9183 8520
rect 9125 8511 9183 8517
rect 9306 8508 9312 8520
rect 9364 8508 9370 8560
rect 1486 8480 1492 8492
rect 1447 8452 1492 8480
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 2866 8440 2872 8492
rect 2924 8440 2930 8492
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8480 6055 8483
rect 6086 8480 6092 8492
rect 6043 8452 6092 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8573 8483 8631 8489
rect 8573 8480 8585 8483
rect 8260 8452 8585 8480
rect 8260 8440 8266 8452
rect 8573 8449 8585 8452
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 8941 8483 8999 8489
rect 8941 8480 8953 8483
rect 8812 8452 8953 8480
rect 8812 8440 8818 8452
rect 8941 8449 8953 8452
rect 8987 8480 8999 8483
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 8987 8452 9229 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 9217 8449 9229 8452
rect 9263 8480 9275 8483
rect 9398 8480 9404 8492
rect 9263 8452 9404 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3283 8384 3985 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 4430 8344 4436 8356
rect 3844 8316 4436 8344
rect 3844 8304 3850 8316
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 8478 8344 8484 8356
rect 6512 8316 8484 8344
rect 6512 8304 6518 8316
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8754 8344 8760 8356
rect 8715 8316 8760 8344
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8344 9459 8347
rect 16574 8344 16580 8356
rect 9447 8316 16580 8344
rect 9447 8313 9459 8316
rect 9401 8307 9459 8313
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 3421 8279 3479 8285
rect 3421 8276 3433 8279
rect 3200 8248 3433 8276
rect 3200 8236 3206 8248
rect 3421 8245 3433 8248
rect 3467 8245 3479 8279
rect 3421 8239 3479 8245
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 2958 8072 2964 8084
rect 2823 8044 2964 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3467 8044 8892 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 4709 8007 4767 8013
rect 4709 7973 4721 8007
rect 4755 8004 4767 8007
rect 4798 8004 4804 8016
rect 4755 7976 4804 8004
rect 4755 7973 4767 7976
rect 4709 7967 4767 7973
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 4614 7936 4620 7948
rect 3068 7908 4620 7936
rect 3068 7877 3096 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 5902 7896 5908 7948
rect 5960 7936 5966 7948
rect 6089 7939 6147 7945
rect 6089 7936 6101 7939
rect 5960 7908 6101 7936
rect 5960 7896 5966 7908
rect 6089 7905 6101 7908
rect 6135 7905 6147 7939
rect 6089 7899 6147 7905
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3602 7868 3608 7880
rect 3563 7840 3608 7868
rect 3053 7831 3111 7837
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3712 7840 4077 7868
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 3326 7800 3332 7812
rect 3283 7772 3332 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 3326 7760 3332 7772
rect 3384 7800 3390 7812
rect 3712 7800 3740 7840
rect 4065 7837 4077 7840
rect 4111 7868 4123 7871
rect 4890 7868 4896 7880
rect 4111 7840 4896 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 6196 7868 6224 8044
rect 8754 7936 8760 7948
rect 7944 7908 8760 7936
rect 6454 7868 6460 7880
rect 6012 7840 6224 7868
rect 6415 7840 6460 7868
rect 3878 7800 3884 7812
rect 3384 7772 3740 7800
rect 3839 7772 3884 7800
rect 3384 7760 3390 7772
rect 3878 7760 3884 7772
rect 3936 7760 3942 7812
rect 6012 7809 6040 7840
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 7944 7877 7972 7908
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 8864 7868 8892 8044
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 9364 8044 9413 8072
rect 9364 8032 9370 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 9033 8007 9091 8013
rect 9033 7973 9045 8007
rect 9079 8004 9091 8007
rect 9490 8004 9496 8016
rect 9079 7976 9496 8004
rect 9079 7973 9091 7976
rect 9033 7967 9091 7973
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 9180 7908 9321 7936
rect 9180 7896 9186 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 8864 7840 16574 7868
rect 7929 7831 7987 7837
rect 5997 7803 6055 7809
rect 5997 7769 6009 7803
rect 6043 7769 6055 7803
rect 8018 7800 8024 7812
rect 7590 7772 8024 7800
rect 5997 7763 6055 7769
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 8493 7803 8551 7809
rect 8493 7769 8505 7803
rect 8539 7800 8551 7803
rect 16546 7800 16574 7840
rect 16666 7800 16672 7812
rect 8539 7772 12572 7800
rect 16546 7772 16672 7800
rect 8539 7769 8551 7772
rect 8493 7763 8551 7769
rect 2958 7732 2964 7744
rect 2919 7704 2964 7732
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 8846 7732 8852 7744
rect 8807 7704 8852 7732
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 12544 7732 12572 7772
rect 16666 7760 16672 7772
rect 16724 7760 16730 7812
rect 16574 7732 16580 7744
rect 12544 7704 16580 7732
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 920 7642 9844 7664
rect 920 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 5194 7642
rect 5246 7590 5258 7642
rect 5310 7590 5322 7642
rect 5374 7590 9844 7642
rect 920 7568 9844 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 3050 7528 3056 7540
rect 2547 7500 3056 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 9398 7528 9404 7540
rect 9359 7500 9404 7528
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 3878 7420 3884 7472
rect 3936 7420 3942 7472
rect 7926 7460 7932 7472
rect 7887 7432 7932 7460
rect 7926 7420 7932 7432
rect 7984 7420 7990 7472
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 9033 7463 9091 7469
rect 9033 7460 9045 7463
rect 8076 7432 9045 7460
rect 8076 7420 8082 7432
rect 9033 7429 9045 7432
rect 9079 7429 9091 7463
rect 9033 7423 9091 7429
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 2958 7392 2964 7404
rect 2823 7364 2964 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4212 7364 4629 7392
rect 4212 7352 4218 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5626 7392 5632 7404
rect 5583 7364 5632 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 8294 7392 8300 7404
rect 6043 7364 8300 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 4982 7284 4988 7336
rect 5040 7324 5046 7336
rect 6012 7324 6040 7355
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9416 7392 9444 7488
rect 9263 7364 9444 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 6178 7324 6184 7336
rect 5040 7296 6040 7324
rect 6139 7296 6184 7324
rect 5040 7284 5046 7296
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 5092 7188 5120 7296
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 8570 7324 8576 7336
rect 8531 7296 8576 7324
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7324 8999 7327
rect 9306 7324 9312 7336
rect 8987 7296 9312 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 5181 7259 5239 7265
rect 5181 7225 5193 7259
rect 5227 7256 5239 7259
rect 6362 7256 6368 7268
rect 5227 7228 6368 7256
rect 5227 7225 5239 7228
rect 5181 7219 5239 7225
rect 6362 7216 6368 7228
rect 6420 7216 6426 7268
rect 5902 7188 5908 7200
rect 2731 7160 5120 7188
rect 5863 7160 5908 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 6512 7160 8033 7188
rect 6512 7148 6518 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 1752 6987 1810 6993
rect 1752 6953 1764 6987
rect 1798 6984 1810 6987
rect 3142 6984 3148 6996
rect 1798 6956 3148 6984
rect 1798 6953 1810 6956
rect 1752 6947 1810 6953
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 6362 6876 6368 6928
rect 6420 6916 6426 6928
rect 6420 6888 6960 6916
rect 6420 6876 6426 6888
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 3283 6820 4169 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 4157 6817 4169 6820
rect 4203 6817 4215 6851
rect 5626 6848 5632 6860
rect 4157 6811 4215 6817
rect 4816 6820 5632 6848
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3786 6780 3792 6792
rect 3108 6752 3792 6780
rect 3108 6740 3114 6752
rect 3786 6740 3792 6752
rect 3844 6780 3850 6792
rect 4816 6789 4844 6820
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 6932 6848 6960 6888
rect 8386 6848 8392 6860
rect 6932 6820 8156 6848
rect 8347 6820 8392 6848
rect 8128 6792 8156 6820
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 9122 6848 9128 6860
rect 8987 6820 9128 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 3844 6752 4353 6780
rect 3844 6740 3850 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6749 5135 6783
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5077 6743 5135 6749
rect 3326 6712 3332 6724
rect 2990 6684 3332 6712
rect 2406 6604 2412 6656
rect 2464 6644 2470 6656
rect 3068 6644 3096 6684
rect 3326 6672 3332 6684
rect 3384 6672 3390 6724
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4617 6715 4675 6721
rect 4617 6712 4629 6715
rect 4304 6684 4629 6712
rect 4304 6672 4310 6684
rect 4617 6681 4629 6684
rect 4663 6681 4675 6715
rect 4617 6675 4675 6681
rect 2464 6616 3096 6644
rect 2464 6604 2470 6616
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3200 6616 3617 6644
rect 3200 6604 3206 6616
rect 3605 6613 3617 6616
rect 3651 6613 3663 6647
rect 5092 6644 5120 6743
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 7374 6780 7380 6792
rect 6963 6752 7380 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7524 6752 7849 6780
rect 7524 6740 7530 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 8110 6780 8116 6792
rect 8071 6752 8116 6780
rect 7837 6743 7895 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 8570 6780 8576 6792
rect 8220 6752 8576 6780
rect 5902 6672 5908 6724
rect 5960 6672 5966 6724
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 6656 6684 7757 6712
rect 6656 6644 6684 6684
rect 7745 6681 7757 6684
rect 7791 6681 7803 6715
rect 7745 6675 7803 6681
rect 8018 6672 8024 6724
rect 8076 6712 8082 6724
rect 8220 6712 8248 6752
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 8076 6684 8248 6712
rect 8297 6715 8355 6721
rect 8076 6672 8082 6684
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 8938 6712 8944 6724
rect 8343 6684 8944 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 9125 6715 9183 6721
rect 9125 6681 9137 6715
rect 9171 6712 9183 6715
rect 9214 6712 9220 6724
rect 9171 6684 9220 6712
rect 9171 6681 9183 6684
rect 9125 6675 9183 6681
rect 9214 6672 9220 6684
rect 9272 6712 9278 6724
rect 9582 6712 9588 6724
rect 9272 6684 9588 6712
rect 9272 6672 9278 6684
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 5092 6616 6684 6644
rect 7481 6647 7539 6653
rect 3605 6607 3663 6613
rect 7481 6613 7493 6647
rect 7527 6644 7539 6647
rect 8202 6644 8208 6656
rect 7527 6616 8208 6644
rect 7527 6613 7539 6616
rect 7481 6607 7539 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 9030 6644 9036 6656
rect 8991 6616 9036 6644
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 9493 6647 9551 6653
rect 9493 6613 9505 6647
rect 9539 6644 9551 6647
rect 9539 6616 16574 6644
rect 9539 6613 9551 6616
rect 9493 6607 9551 6613
rect 920 6554 9844 6576
rect 920 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 5194 6554
rect 5246 6502 5258 6554
rect 5310 6502 5322 6554
rect 5374 6502 9844 6554
rect 920 6480 9844 6502
rect 16546 6452 16574 6616
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 3050 6440 3056 6452
rect 2271 6412 3056 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 7374 6400 7380 6452
rect 7432 6440 7438 6452
rect 7432 6412 7788 6440
rect 7432 6400 7438 6412
rect 4252 6384 4304 6390
rect 1578 6332 1584 6384
rect 1636 6372 1642 6384
rect 2041 6375 2099 6381
rect 2041 6372 2053 6375
rect 1636 6344 2053 6372
rect 1636 6332 1642 6344
rect 2041 6341 2053 6344
rect 2087 6372 2099 6375
rect 2406 6372 2412 6384
rect 2087 6344 2412 6372
rect 2087 6341 2099 6344
rect 2041 6335 2099 6341
rect 2406 6332 2412 6344
rect 2464 6332 2470 6384
rect 6730 6372 6736 6384
rect 4252 6326 4304 6332
rect 6196 6344 6736 6372
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 3142 6304 3148 6316
rect 2731 6276 2912 6304
rect 3103 6276 3148 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 2593 6239 2651 6245
rect 2593 6205 2605 6239
rect 2639 6236 2651 6239
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 2639 6208 2789 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 2777 6205 2789 6208
rect 2823 6205 2835 6239
rect 2777 6199 2835 6205
rect 2884 6100 2912 6276
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 4614 6304 4620 6316
rect 4575 6276 4620 6304
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6304 5411 6307
rect 5442 6304 5448 6316
rect 5399 6276 5448 6304
rect 5399 6273 5411 6276
rect 5353 6267 5411 6273
rect 5442 6264 5448 6276
rect 5500 6304 5506 6316
rect 5500 6276 6040 6304
rect 5500 6264 5506 6276
rect 5902 6236 5908 6248
rect 5863 6208 5908 6236
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 6012 6236 6040 6276
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 6196 6313 6224 6344
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 7760 6372 7788 6412
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 7984 6412 8125 6440
rect 7984 6400 7990 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 8113 6403 8171 6409
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8444 6412 8953 6440
rect 8444 6400 8450 6412
rect 8941 6409 8953 6412
rect 8987 6409 8999 6443
rect 8941 6403 8999 6409
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9398 6440 9404 6452
rect 9079 6412 9404 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 9490 6400 9496 6452
rect 9548 6440 9554 6452
rect 9548 6412 9593 6440
rect 16546 6412 16580 6452
rect 9548 6400 9554 6412
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 8297 6375 8355 6381
rect 8297 6372 8309 6375
rect 7760 6344 8309 6372
rect 8297 6341 8309 6344
rect 8343 6341 8355 6375
rect 8297 6335 8355 6341
rect 8757 6375 8815 6381
rect 8757 6341 8769 6375
rect 8803 6372 8815 6375
rect 8846 6372 8852 6384
rect 8803 6344 8852 6372
rect 8803 6341 8815 6344
rect 8757 6335 8815 6341
rect 8846 6332 8852 6344
rect 8904 6332 8910 6384
rect 9122 6372 9128 6384
rect 9083 6344 9128 6372
rect 9122 6332 9128 6344
rect 9180 6332 9186 6384
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 6144 6276 6193 6304
rect 6144 6264 6150 6276
rect 6181 6273 6193 6276
rect 6227 6273 6239 6307
rect 8202 6304 8208 6316
rect 7590 6276 8208 6304
rect 6181 6267 6239 6273
rect 8202 6264 8208 6276
rect 8260 6304 8266 6316
rect 8386 6304 8392 6316
rect 8260 6276 8392 6304
rect 8260 6264 8266 6276
rect 8386 6264 8392 6276
rect 8444 6304 8450 6316
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8444 6276 8493 6304
rect 8444 6264 8450 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8628 6276 8677 6304
rect 8628 6264 8634 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6012 6208 6469 6236
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8018 6236 8024 6248
rect 7975 6208 8024 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8294 6196 8300 6248
rect 8352 6236 8358 6248
rect 8680 6236 8708 6267
rect 8352 6208 8708 6236
rect 8352 6196 8358 6208
rect 9309 6171 9367 6177
rect 9309 6137 9321 6171
rect 9355 6168 9367 6171
rect 19426 6168 19432 6180
rect 9355 6140 19432 6168
rect 9355 6137 9367 6140
rect 9309 6131 9367 6137
rect 19426 6128 19432 6140
rect 19484 6128 19490 6180
rect 4982 6100 4988 6112
rect 2884 6072 4988 6100
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5181 6103 5239 6109
rect 5181 6069 5193 6103
rect 5227 6100 5239 6103
rect 5442 6100 5448 6112
rect 5227 6072 5448 6100
rect 5227 6069 5239 6072
rect 5181 6063 5239 6069
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 1489 5899 1547 5905
rect 1489 5865 1501 5899
rect 1535 5896 1547 5899
rect 1578 5896 1584 5908
rect 1535 5868 1584 5896
rect 1535 5865 1547 5868
rect 1489 5859 1547 5865
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 1844 5899 1902 5905
rect 1844 5865 1856 5899
rect 1890 5896 1902 5899
rect 3142 5896 3148 5908
rect 1890 5868 3148 5896
rect 1890 5865 1902 5868
rect 1844 5859 1902 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4614 5896 4620 5908
rect 4019 5868 4620 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5902 5896 5908 5908
rect 5863 5868 5908 5896
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 8202 5896 8208 5908
rect 8163 5868 8208 5896
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8389 5831 8447 5837
rect 8389 5828 8401 5831
rect 8168 5800 8401 5828
rect 8168 5788 8174 5800
rect 8389 5797 8401 5800
rect 8435 5828 8447 5831
rect 8435 5800 12434 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 1581 5763 1639 5769
rect 1581 5760 1593 5763
rect 1544 5732 1593 5760
rect 1544 5720 1550 5732
rect 1581 5729 1593 5732
rect 1627 5729 1639 5763
rect 1581 5723 1639 5729
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 5718 5760 5724 5772
rect 4479 5732 5724 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 6086 5720 6092 5772
rect 6144 5760 6150 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 6144 5732 6193 5760
rect 6144 5720 6150 5732
rect 6181 5729 6193 5732
rect 6227 5729 6239 5763
rect 6454 5760 6460 5772
rect 6415 5732 6460 5760
rect 6181 5723 6239 5729
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5760 7987 5763
rect 8846 5760 8852 5772
rect 7975 5732 8852 5760
rect 7975 5729 7987 5732
rect 7929 5723 7987 5729
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 3384 5664 4169 5692
rect 3384 5652 3390 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 3697 5627 3755 5633
rect 3082 5596 3648 5624
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 3418 5556 3424 5568
rect 3375 5528 3424 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 3620 5556 3648 5596
rect 3697 5593 3709 5627
rect 3743 5624 3755 5627
rect 3786 5624 3792 5636
rect 3743 5596 3792 5624
rect 3743 5593 3755 5596
rect 3697 5587 3755 5593
rect 3786 5584 3792 5596
rect 3844 5584 3850 5636
rect 3881 5627 3939 5633
rect 3881 5593 3893 5627
rect 3927 5624 3939 5627
rect 4890 5624 4896 5636
rect 3927 5596 4896 5624
rect 3927 5593 3939 5596
rect 3881 5587 3939 5593
rect 3896 5556 3924 5587
rect 4890 5584 4896 5596
rect 4948 5584 4954 5636
rect 8202 5624 8208 5636
rect 5658 5596 6500 5624
rect 7682 5596 8208 5624
rect 3620 5528 3924 5556
rect 6472 5556 6500 5596
rect 7760 5556 7788 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 8849 5627 8907 5633
rect 8849 5593 8861 5627
rect 8895 5593 8907 5627
rect 8849 5587 8907 5593
rect 6472 5528 7788 5556
rect 8864 5556 8892 5587
rect 8938 5584 8944 5636
rect 8996 5624 9002 5636
rect 9490 5624 9496 5636
rect 8996 5596 9041 5624
rect 9451 5596 9496 5624
rect 8996 5584 9002 5596
rect 9490 5584 9496 5596
rect 9548 5584 9554 5636
rect 9122 5556 9128 5568
rect 8864 5528 9128 5556
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 12406 5556 12434 5800
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 16666 5624 16672 5636
rect 13872 5596 16672 5624
rect 13872 5584 13878 5596
rect 16666 5584 16672 5596
rect 16724 5584 16730 5636
rect 16574 5556 16580 5568
rect 12406 5528 16580 5556
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 920 5466 9844 5488
rect 920 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 5194 5466
rect 5246 5414 5258 5466
rect 5310 5414 5322 5466
rect 5374 5414 9844 5466
rect 920 5392 9844 5414
rect 3878 5352 3884 5364
rect 3620 5324 3884 5352
rect 3620 5293 3648 5324
rect 3878 5312 3884 5324
rect 3936 5352 3942 5364
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 3936 5324 5273 5352
rect 3936 5312 3942 5324
rect 5261 5321 5273 5324
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 7064 5324 8309 5352
rect 7064 5312 7070 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 8297 5315 8355 5321
rect 3605 5287 3663 5293
rect 3605 5253 3617 5287
rect 3651 5253 3663 5287
rect 4890 5284 4896 5296
rect 4830 5256 4896 5284
rect 3605 5247 3663 5253
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 8113 5287 8171 5293
rect 8113 5284 8125 5287
rect 7498 5256 8125 5284
rect 8113 5253 8125 5256
rect 8159 5284 8171 5287
rect 8202 5284 8208 5296
rect 8159 5256 8208 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 8478 5244 8484 5296
rect 8536 5284 8542 5296
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 8536 5256 9045 5284
rect 8536 5244 8542 5256
rect 9033 5253 9045 5256
rect 9079 5253 9091 5287
rect 9033 5247 9091 5253
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 3326 5216 3332 5228
rect 1544 5188 3332 5216
rect 1544 5176 1550 5188
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 5994 5216 6000 5228
rect 5955 5188 6000 5216
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 8220 5216 8248 5244
rect 8754 5216 8760 5228
rect 8220 5188 8760 5216
rect 8754 5176 8760 5188
rect 8812 5216 8818 5228
rect 9214 5216 9220 5228
rect 8812 5188 9220 5216
rect 8812 5176 8818 5188
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 5166 5108 5172 5160
rect 5224 5148 5230 5160
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5224 5120 5825 5148
rect 5224 5108 5230 5120
rect 5813 5117 5825 5120
rect 5859 5117 5871 5151
rect 5813 5111 5871 5117
rect 6273 5151 6331 5157
rect 6273 5117 6285 5151
rect 6319 5148 6331 5151
rect 6914 5148 6920 5160
rect 6319 5120 6920 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5148 7803 5151
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 7791 5120 8861 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 5074 5012 5080 5024
rect 5035 4984 5080 5012
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 9309 5015 9367 5021
rect 9309 5012 9321 5015
rect 8444 4984 9321 5012
rect 8444 4972 8450 4984
rect 9309 4981 9321 4984
rect 9355 4981 9367 5015
rect 9309 4975 9367 4981
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 5718 4808 5724 4820
rect 5679 4780 5724 4808
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9272 4780 9413 4808
rect 9272 4768 9278 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 5074 4700 5080 4752
rect 5132 4740 5138 4752
rect 5132 4712 6316 4740
rect 5132 4700 5138 4712
rect 3326 4672 3332 4684
rect 3287 4644 3332 4672
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 6288 4681 6316 4712
rect 5353 4675 5411 4681
rect 5353 4672 5365 4675
rect 4212 4644 5365 4672
rect 4212 4632 4218 4644
rect 5353 4641 5365 4644
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 4982 4564 4988 4616
rect 5040 4604 5046 4616
rect 5442 4604 5448 4616
rect 5040 4576 5448 4604
rect 5040 4564 5046 4576
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7006 4604 7012 4616
rect 6963 4576 7012 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 8386 4604 8392 4616
rect 8347 4576 8392 4604
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9306 4604 9312 4616
rect 9180 4576 9312 4604
rect 9180 4564 9186 4576
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 3605 4539 3663 4545
rect 3605 4505 3617 4539
rect 3651 4505 3663 4539
rect 4890 4536 4896 4548
rect 4803 4508 4896 4536
rect 3605 4499 3663 4505
rect 3620 4468 3648 4499
rect 4890 4496 4896 4508
rect 4948 4536 4954 4548
rect 5534 4536 5540 4548
rect 4948 4508 5540 4536
rect 4948 4496 4954 4508
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 7466 4496 7472 4548
rect 7524 4496 7530 4548
rect 4338 4468 4344 4480
rect 3620 4440 4344 4468
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 5077 4471 5135 4477
rect 5077 4437 5089 4471
rect 5123 4468 5135 4471
rect 5166 4468 5172 4480
rect 5123 4440 5172 4468
rect 5123 4437 5135 4440
rect 5077 4431 5135 4437
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 8938 4428 8944 4480
rect 8996 4477 9002 4480
rect 8996 4468 9007 4477
rect 9214 4468 9220 4480
rect 8996 4440 9041 4468
rect 9175 4440 9220 4468
rect 8996 4431 9007 4440
rect 8996 4428 9002 4431
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 3036 4378 9844 4400
rect 3036 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 5194 4378
rect 5246 4326 5258 4378
rect 5310 4326 5322 4378
rect 5374 4326 9844 4378
rect 3036 4304 9844 4326
rect 6365 4267 6423 4273
rect 6365 4233 6377 4267
rect 6411 4264 6423 4267
rect 6546 4264 6552 4276
rect 6411 4236 6552 4264
rect 6411 4233 6423 4236
rect 6365 4227 6423 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 8754 4224 8760 4276
rect 8812 4264 8818 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 8812 4236 9045 4264
rect 8812 4224 8818 4236
rect 9033 4233 9045 4236
rect 9079 4264 9091 4267
rect 9217 4267 9275 4273
rect 9217 4264 9229 4267
rect 9079 4236 9229 4264
rect 9079 4233 9091 4236
rect 9033 4227 9091 4233
rect 9217 4233 9229 4236
rect 9263 4233 9275 4267
rect 9217 4227 9275 4233
rect 5810 4196 5816 4208
rect 5014 4168 5816 4196
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3292 4100 3341 4128
rect 3292 4088 3298 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 5350 4128 5356 4140
rect 3559 4100 4016 4128
rect 5311 4100 5356 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3878 4060 3884 4072
rect 3839 4032 3884 4060
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 3988 4060 4016 4100
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 6273 4131 6331 4137
rect 6273 4128 6285 4131
rect 5500 4100 6285 4128
rect 5500 4088 5506 4100
rect 6273 4097 6285 4100
rect 6319 4097 6331 4131
rect 6273 4091 6331 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 9214 4128 9220 4140
rect 8159 4100 9220 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4128 9551 4131
rect 9582 4128 9588 4140
rect 9539 4100 9588 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 4154 4060 4160 4072
rect 3988 4032 4160 4060
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 6549 4063 6607 4069
rect 6549 4029 6561 4063
rect 6595 4029 6607 4063
rect 6549 4023 6607 4029
rect 2682 3952 2688 4004
rect 2740 3992 2746 4004
rect 6564 3992 6592 4023
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 6972 4032 8309 4060
rect 6972 4020 6978 4032
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 8846 4060 8852 4072
rect 8807 4032 8852 4060
rect 8297 4023 8355 4029
rect 8846 4020 8852 4032
rect 8904 4020 8910 4072
rect 2740 3964 3648 3992
rect 2740 3952 2746 3964
rect 3620 3924 3648 3964
rect 4816 3964 6592 3992
rect 8021 3995 8079 4001
rect 4816 3924 4844 3964
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 13814 3992 13820 4004
rect 8067 3964 13820 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 5902 3924 5908 3936
rect 5960 3933 5966 3936
rect 3620 3896 4844 3924
rect 5871 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3887 5971 3933
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6546 3924 6552 3936
rect 6227 3896 6552 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 5960 3884 5966 3887
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 5445 3723 5503 3729
rect 5445 3720 5457 3723
rect 5408 3692 5457 3720
rect 5408 3680 5414 3692
rect 5445 3689 5457 3692
rect 5491 3689 5503 3723
rect 5810 3720 5816 3732
rect 5771 3692 5816 3720
rect 5445 3683 5503 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 9398 3720 9404 3732
rect 9359 3692 9404 3720
rect 9398 3680 9404 3692
rect 9456 3720 9462 3732
rect 9582 3720 9588 3732
rect 9456 3692 9588 3720
rect 9456 3680 9462 3692
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 3384 3556 3433 3584
rect 3384 3544 3390 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 6972 3556 7205 3584
rect 6972 3544 6978 3556
rect 7193 3553 7205 3556
rect 7239 3553 7251 3587
rect 7193 3547 7251 3553
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 4856 3488 5089 3516
rect 4856 3476 4862 3488
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5077 3479 5135 3485
rect 5184 3488 5733 3516
rect 4430 3408 4436 3460
rect 4488 3448 4494 3460
rect 5184 3457 5212 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3516 6239 3519
rect 6227 3488 6592 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 5169 3451 5227 3457
rect 5169 3448 5181 3451
rect 4488 3420 5181 3448
rect 4488 3408 4494 3420
rect 5169 3417 5181 3420
rect 5215 3417 5227 3451
rect 5169 3411 5227 3417
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 5534 3448 5540 3460
rect 5399 3420 5540 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 5534 3408 5540 3420
rect 5592 3448 5598 3460
rect 6196 3448 6224 3479
rect 6564 3460 6592 3488
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6696 3488 6745 3516
rect 6696 3476 6702 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7006 3516 7012 3528
rect 6871 3488 7012 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 8536 3488 8677 3516
rect 8536 3476 8542 3488
rect 8665 3485 8677 3488
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 5592 3420 6224 3448
rect 6365 3451 6423 3457
rect 5592 3408 5598 3420
rect 6365 3417 6377 3451
rect 6411 3448 6423 3451
rect 6454 3448 6460 3460
rect 6411 3420 6460 3448
rect 6411 3417 6423 3420
rect 6365 3411 6423 3417
rect 6454 3408 6460 3420
rect 6512 3408 6518 3460
rect 6546 3408 6552 3460
rect 6604 3448 6610 3460
rect 6604 3420 6649 3448
rect 6604 3408 6610 3420
rect 7926 3408 7932 3460
rect 7984 3408 7990 3460
rect 9229 3451 9287 3457
rect 9229 3417 9241 3451
rect 9275 3448 9287 3451
rect 9275 3420 16574 3448
rect 9275 3417 9287 3420
rect 9229 3411 9287 3417
rect 16546 3392 16574 3420
rect 8849 3383 8907 3389
rect 8849 3349 8861 3383
rect 8895 3380 8907 3383
rect 8938 3380 8944 3392
rect 8895 3352 8944 3380
rect 8895 3349 8907 3352
rect 8849 3343 8907 3349
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 16546 3352 16580 3392
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 3036 3290 9844 3312
rect 3036 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 5194 3290
rect 5246 3238 5258 3290
rect 5310 3238 5322 3290
rect 5374 3238 9844 3290
rect 3036 3216 9844 3238
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4338 3176 4344 3188
rect 4203 3148 4344 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 4430 3136 4436 3188
rect 4488 3136 4494 3188
rect 7929 3179 7987 3185
rect 7929 3176 7941 3179
rect 7760 3148 7941 3176
rect 3421 3111 3479 3117
rect 3421 3077 3433 3111
rect 3467 3108 3479 3111
rect 4448 3108 4476 3136
rect 3467 3080 4476 3108
rect 6092 3120 6144 3126
rect 3467 3077 3479 3080
rect 3421 3071 3479 3077
rect 7466 3108 7472 3120
rect 7427 3080 7472 3108
rect 7466 3068 7472 3080
rect 7524 3068 7530 3120
rect 6092 3062 6144 3068
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4890 3040 4896 3052
rect 4479 3012 4896 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 6454 3040 6460 3052
rect 6415 3012 6460 3040
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6546 3000 6552 3052
rect 6604 3040 6610 3052
rect 7760 3049 7788 3148
rect 7929 3145 7941 3148
rect 7975 3176 7987 3179
rect 8386 3176 8392 3188
rect 7975 3148 8392 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8386 3136 8392 3148
rect 8444 3176 8450 3188
rect 8481 3179 8539 3185
rect 8481 3176 8493 3179
rect 8444 3148 8493 3176
rect 8444 3136 8450 3148
rect 8481 3145 8493 3148
rect 8527 3145 8539 3179
rect 8938 3176 8944 3188
rect 8899 3148 8944 3176
rect 8481 3139 8539 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9088 3148 9413 3176
rect 9088 3136 9094 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 8110 3108 8116 3120
rect 8023 3080 8116 3108
rect 8110 3068 8116 3080
rect 8168 3108 8174 3120
rect 8297 3111 8355 3117
rect 8297 3108 8309 3111
rect 8168 3080 8309 3108
rect 8168 3068 8174 3080
rect 8297 3077 8309 3080
rect 8343 3108 8355 3111
rect 8754 3108 8760 3120
rect 8343 3080 8760 3108
rect 8343 3077 8355 3080
rect 8297 3071 8355 3077
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 7255 3043 7313 3049
rect 7255 3040 7267 3043
rect 6604 3012 7267 3040
rect 6604 3000 6610 3012
rect 7255 3009 7267 3012
rect 7301 3009 7313 3043
rect 7255 3003 7313 3009
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9306 3040 9312 3052
rect 9079 3012 9312 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 3476 2944 3617 2972
rect 3476 2932 3482 2944
rect 3605 2941 3617 2944
rect 3651 2941 3663 2975
rect 4614 2972 4620 2984
rect 4575 2944 4620 2972
rect 3605 2935 3663 2941
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 5626 2972 5632 2984
rect 5031 2944 5632 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2972 8907 2975
rect 9214 2972 9220 2984
rect 8895 2944 9220 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 7021 2907 7079 2913
rect 7021 2873 7033 2907
rect 7067 2904 7079 2907
rect 8202 2904 8208 2916
rect 7067 2876 8208 2904
rect 7067 2873 7079 2876
rect 7021 2867 7079 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 4338 2836 4344 2848
rect 4299 2808 4344 2836
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 3036 2672 9844 2694
rect 4614 2592 4620 2644
rect 4672 2632 4678 2644
rect 4801 2635 4859 2641
rect 4801 2632 4813 2635
rect 4672 2604 4813 2632
rect 4672 2592 4678 2604
rect 4801 2601 4813 2604
rect 4847 2601 4859 2635
rect 6086 2632 6092 2644
rect 6047 2604 6092 2632
rect 4801 2595 4859 2601
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 6641 2635 6699 2641
rect 6641 2601 6653 2635
rect 6687 2632 6699 2635
rect 6730 2632 6736 2644
rect 6687 2604 6736 2632
rect 6687 2601 6699 2604
rect 6641 2595 6699 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 7006 2632 7012 2644
rect 6967 2604 7012 2632
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2601 7343 2635
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7285 2595 7343 2601
rect 4430 2524 4436 2576
rect 4488 2564 4494 2576
rect 5077 2567 5135 2573
rect 5077 2564 5089 2567
rect 4488 2536 5089 2564
rect 4488 2524 4494 2536
rect 5077 2533 5089 2536
rect 5123 2533 5135 2567
rect 5077 2527 5135 2533
rect 6457 2567 6515 2573
rect 6457 2533 6469 2567
rect 6503 2564 6515 2567
rect 6546 2564 6552 2576
rect 6503 2536 6552 2564
rect 6503 2533 6515 2536
rect 6457 2527 6515 2533
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 3467 2468 5365 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3620 2437 3648 2468
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3605 2391 3663 2397
rect 3712 2400 3985 2428
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 3712 2360 3740 2400
rect 3973 2397 3985 2400
rect 4019 2428 4031 2431
rect 4154 2428 4160 2440
rect 4019 2400 4160 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 4356 2437 4384 2468
rect 5353 2465 5365 2468
rect 5399 2496 5411 2499
rect 5442 2496 5448 2508
rect 5399 2468 5448 2496
rect 5399 2465 5411 2468
rect 5353 2459 5411 2465
rect 5442 2456 5448 2468
rect 5500 2496 5506 2508
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 5500 2468 5549 2496
rect 5500 2456 5506 2468
rect 5537 2465 5549 2468
rect 5583 2496 5595 2499
rect 5583 2468 6224 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2397 4399 2431
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 4341 2391 4399 2397
rect 4890 2388 4896 2400
rect 4948 2428 4954 2440
rect 6196 2437 6224 2468
rect 5905 2431 5963 2437
rect 4948 2400 5304 2428
rect 4948 2388 4954 2400
rect 3292 2332 3740 2360
rect 3789 2363 3847 2369
rect 3292 2320 3298 2332
rect 3789 2329 3801 2363
rect 3835 2360 3847 2363
rect 4062 2360 4068 2372
rect 3835 2332 4068 2360
rect 3835 2329 3847 2332
rect 3789 2323 3847 2329
rect 4062 2320 4068 2332
rect 4120 2320 4126 2372
rect 4525 2363 4583 2369
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 4982 2360 4988 2372
rect 4571 2332 4988 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 5276 2292 5304 2400
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6472 2428 6500 2527
rect 6546 2524 6552 2536
rect 6604 2564 6610 2576
rect 6825 2567 6883 2573
rect 6825 2564 6837 2567
rect 6604 2536 6837 2564
rect 6604 2524 6610 2536
rect 6825 2533 6837 2536
rect 6871 2564 6883 2567
rect 7300 2564 7328 2595
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 9030 2632 9036 2644
rect 8991 2604 9036 2632
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9214 2632 9220 2644
rect 9175 2604 9220 2632
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 8110 2564 8116 2576
rect 6871 2536 8116 2564
rect 6871 2533 6883 2536
rect 6825 2527 6883 2533
rect 7576 2437 7604 2536
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 8478 2564 8484 2576
rect 8439 2536 8484 2564
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 9122 2524 9128 2576
rect 9180 2564 9186 2576
rect 9401 2567 9459 2573
rect 9401 2564 9413 2567
rect 9180 2536 9413 2564
rect 9180 2524 9186 2536
rect 9401 2533 9413 2536
rect 9447 2533 9459 2567
rect 9401 2527 9459 2533
rect 8128 2496 8156 2524
rect 8128 2468 8340 2496
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6227 2400 6500 2428
rect 6840 2400 6929 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 5920 2360 5948 2391
rect 5994 2360 6000 2372
rect 5907 2332 6000 2360
rect 5994 2320 6000 2332
rect 6052 2360 6058 2372
rect 6730 2360 6736 2372
rect 6052 2332 6736 2360
rect 6052 2320 6058 2332
rect 6730 2320 6736 2332
rect 6788 2320 6794 2372
rect 6840 2292 6868 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 7834 2428 7840 2440
rect 7795 2400 7840 2428
rect 7561 2391 7619 2397
rect 7834 2388 7840 2400
rect 7892 2428 7898 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7892 2400 8125 2428
rect 7892 2388 7898 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8312 2372 8340 2468
rect 8662 2428 8668 2440
rect 8623 2400 8668 2428
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 8294 2360 8300 2372
rect 8207 2332 8300 2360
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 9079 2363 9137 2369
rect 9079 2329 9091 2363
rect 9125 2360 9137 2363
rect 9582 2360 9588 2372
rect 9125 2332 9588 2360
rect 9125 2329 9137 2332
rect 9079 2323 9137 2329
rect 9582 2320 9588 2332
rect 9640 2320 9646 2372
rect 5276 2264 6868 2292
rect 3036 2202 9844 2224
rect 3036 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 5194 2202
rect 5246 2150 5258 2202
rect 5310 2150 5322 2202
rect 5374 2150 9844 2202
rect 3036 2128 9844 2150
rect 4338 2088 4344 2100
rect 3344 2060 4344 2088
rect 3344 1961 3372 2060
rect 4338 2048 4344 2060
rect 4396 2048 4402 2100
rect 5733 2091 5791 2097
rect 5733 2057 5745 2091
rect 5779 2088 5791 2091
rect 6822 2088 6828 2100
rect 5779 2060 6828 2088
rect 5779 2057 5791 2060
rect 5733 2051 5791 2057
rect 6822 2048 6828 2060
rect 6880 2048 6886 2100
rect 8294 2088 8300 2100
rect 8255 2060 8300 2088
rect 8294 2048 8300 2060
rect 8352 2088 8358 2100
rect 8573 2091 8631 2097
rect 8573 2088 8585 2091
rect 8352 2060 8585 2088
rect 8352 2048 8358 2060
rect 8573 2057 8585 2060
rect 8619 2057 8631 2091
rect 8573 2051 8631 2057
rect 8662 2048 8668 2100
rect 8720 2088 8726 2100
rect 8757 2091 8815 2097
rect 8757 2088 8769 2091
rect 8720 2060 8769 2088
rect 8720 2048 8726 2060
rect 8757 2057 8769 2060
rect 8803 2057 8815 2091
rect 9306 2088 9312 2100
rect 9267 2060 9312 2088
rect 8757 2051 8815 2057
rect 9306 2048 9312 2060
rect 9364 2048 9370 2100
rect 4062 1980 4068 2032
rect 4120 1980 4126 2032
rect 5994 2020 6000 2032
rect 5955 1992 6000 2020
rect 5994 1980 6000 1992
rect 6052 1980 6058 2032
rect 6270 1980 6276 2032
rect 6328 2020 6334 2032
rect 7285 2023 7343 2029
rect 7285 2020 7297 2023
rect 6328 1992 7297 2020
rect 6328 1980 6334 1992
rect 7285 1989 7297 1992
rect 7331 2020 7343 2023
rect 7834 2020 7840 2032
rect 7331 1992 7840 2020
rect 7331 1989 7343 1992
rect 7285 1983 7343 1989
rect 7834 1980 7840 1992
rect 7892 2020 7898 2032
rect 7929 2023 7987 2029
rect 7929 2020 7941 2023
rect 7892 1992 7941 2020
rect 7892 1980 7898 1992
rect 7929 1989 7941 1992
rect 7975 1989 7987 2023
rect 7929 1983 7987 1989
rect 9122 1980 9128 2032
rect 9180 2020 9186 2032
rect 9401 2023 9459 2029
rect 9401 2020 9413 2023
rect 9180 1992 9413 2020
rect 9180 1980 9186 1992
rect 9401 1989 9413 1992
rect 9447 1989 9459 2023
rect 9401 1983 9459 1989
rect 3329 1955 3387 1961
rect 3329 1921 3341 1955
rect 3375 1921 3387 1955
rect 3329 1915 3387 1921
rect 4982 1912 4988 1964
rect 5040 1952 5046 1964
rect 5169 1955 5227 1961
rect 5169 1952 5181 1955
rect 5040 1924 5181 1952
rect 5040 1912 5046 1924
rect 5169 1921 5181 1924
rect 5215 1921 5227 1955
rect 5169 1915 5227 1921
rect 3697 1887 3755 1893
rect 3697 1853 3709 1887
rect 3743 1884 3755 1887
rect 4246 1884 4252 1896
rect 3743 1856 4252 1884
rect 3743 1853 3755 1856
rect 3697 1847 3755 1853
rect 4246 1844 4252 1856
rect 4304 1844 4310 1896
rect 9122 1884 9128 1896
rect 9083 1856 9128 1884
rect 9122 1844 9128 1856
rect 9180 1844 9186 1896
rect 8938 1748 8944 1760
rect 8899 1720 8944 1748
rect 8938 1708 8944 1720
rect 8996 1708 9002 1760
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 4154 1504 4160 1556
rect 4212 1544 4218 1556
rect 5353 1547 5411 1553
rect 5353 1544 5365 1547
rect 4212 1516 5365 1544
rect 4212 1504 4218 1516
rect 5353 1513 5365 1516
rect 5399 1513 5411 1547
rect 5353 1507 5411 1513
rect 9493 1547 9551 1553
rect 9493 1513 9505 1547
rect 9539 1544 9551 1547
rect 9582 1544 9588 1556
rect 9539 1516 9588 1544
rect 9539 1513 9551 1516
rect 9493 1507 9551 1513
rect 9582 1504 9588 1516
rect 9640 1504 9646 1556
rect 5261 1479 5319 1485
rect 5261 1445 5273 1479
rect 5307 1476 5319 1479
rect 5442 1476 5448 1488
rect 5307 1448 5448 1476
rect 5307 1445 5319 1448
rect 5261 1439 5319 1445
rect 5442 1436 5448 1448
rect 5500 1436 5506 1488
rect 5077 1343 5135 1349
rect 5077 1309 5089 1343
rect 5123 1340 5135 1343
rect 6178 1340 6184 1352
rect 5123 1312 6184 1340
rect 5123 1309 5135 1312
rect 5077 1303 5135 1309
rect 6178 1300 6184 1312
rect 6236 1300 6242 1352
rect 3789 1207 3847 1213
rect 3789 1173 3801 1207
rect 3835 1204 3847 1207
rect 4890 1204 4896 1216
rect 3835 1176 4896 1204
rect 3835 1173 3847 1176
rect 3789 1167 3847 1173
rect 4890 1164 4896 1176
rect 4948 1164 4954 1216
rect 3036 1114 9844 1136
rect 3036 1062 5066 1114
rect 5118 1062 5130 1114
rect 5182 1062 5194 1114
rect 5246 1062 5258 1114
rect 5310 1062 5322 1114
rect 5374 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 1768 11296 1820 11348
rect 4344 11296 4396 11348
rect 6460 11296 6512 11348
rect 8116 11296 8168 11348
rect 1216 11228 1268 11280
rect 6552 11228 6604 11280
rect 4712 11160 4764 11212
rect 5540 11160 5592 11212
rect 6276 11160 6328 11212
rect 7288 11160 7340 11212
rect 4344 11135 4396 11144
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 4988 11092 5040 11144
rect 4252 11067 4304 11076
rect 4252 11033 4261 11067
rect 4261 11033 4295 11067
rect 4295 11033 4304 11067
rect 4252 11024 4304 11033
rect 5632 11024 5684 11076
rect 6828 11092 6880 11144
rect 7472 11024 7524 11076
rect 4620 10999 4672 11008
rect 4620 10965 4629 10999
rect 4629 10965 4663 10999
rect 4663 10965 4672 10999
rect 4620 10956 4672 10965
rect 5540 10956 5592 11008
rect 7288 10999 7340 11008
rect 7288 10965 7297 10999
rect 7297 10965 7331 10999
rect 7331 10965 7340 10999
rect 7288 10956 7340 10965
rect 7656 10956 7708 11008
rect 16580 11024 16632 11076
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5194 10854 5246 10906
rect 5258 10854 5310 10906
rect 5322 10854 5374 10906
rect 6000 10752 6052 10804
rect 6460 10752 6512 10804
rect 4528 10684 4580 10736
rect 4712 10684 4764 10736
rect 2964 10616 3016 10668
rect 4344 10616 4396 10668
rect 4988 10616 5040 10668
rect 8208 10684 8260 10736
rect 6552 10659 6604 10668
rect 1584 10548 1636 10600
rect 1768 10412 1820 10464
rect 5632 10548 5684 10600
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 7288 10548 7340 10600
rect 9404 10616 9456 10668
rect 4896 10412 4948 10464
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 6000 10412 6052 10464
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 7104 10455 7156 10464
rect 7104 10421 7113 10455
rect 7113 10421 7147 10455
rect 7147 10421 7156 10455
rect 7104 10412 7156 10421
rect 7196 10412 7248 10464
rect 16580 10412 16632 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 4528 10208 4580 10260
rect 1492 10004 1544 10056
rect 2320 9936 2372 9988
rect 4620 10072 4672 10124
rect 6000 10208 6052 10260
rect 4712 10004 4764 10056
rect 5540 10072 5592 10124
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 7104 10004 7156 10056
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 6368 9936 6420 9988
rect 8300 9979 8352 9988
rect 8300 9945 8309 9979
rect 8309 9945 8343 9979
rect 8343 9945 8352 9979
rect 8300 9936 8352 9945
rect 8852 9936 8904 9988
rect 3700 9868 3752 9920
rect 4160 9868 4212 9920
rect 9128 9868 9180 9920
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5194 9766 5246 9818
rect 5258 9766 5310 9818
rect 5322 9766 5374 9818
rect 1492 9664 1544 9716
rect 2320 9596 2372 9648
rect 4528 9664 4580 9716
rect 4896 9664 4948 9716
rect 5816 9664 5868 9716
rect 4252 9596 4304 9648
rect 6000 9639 6052 9648
rect 6000 9605 6009 9639
rect 6009 9605 6043 9639
rect 6043 9605 6052 9639
rect 6000 9596 6052 9605
rect 8300 9596 8352 9648
rect 1584 9460 1636 9512
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 5632 9528 5684 9580
rect 7196 9528 7248 9580
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 4160 9460 4212 9512
rect 6736 9503 6788 9512
rect 6736 9469 6745 9503
rect 6745 9469 6779 9503
rect 6779 9469 6788 9503
rect 6736 9460 6788 9469
rect 8024 9460 8076 9512
rect 4436 9324 4488 9376
rect 6644 9324 6696 9376
rect 8392 9324 8444 9376
rect 8668 9324 8720 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 1952 9120 2004 9172
rect 2412 9120 2464 9172
rect 2964 9120 3016 9172
rect 3608 9120 3660 9172
rect 4160 9120 4212 9172
rect 6736 9120 6788 9172
rect 8208 9163 8260 9172
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 4344 9052 4396 9104
rect 6828 8984 6880 9036
rect 2320 8916 2372 8968
rect 2872 8916 2924 8968
rect 3148 8848 3200 8900
rect 3608 8916 3660 8968
rect 5632 8848 5684 8900
rect 6000 8848 6052 8900
rect 7012 8848 7064 8900
rect 8760 8848 8812 8900
rect 16764 8984 16816 9036
rect 9312 8823 9364 8832
rect 9312 8789 9321 8823
rect 9321 8789 9355 8823
rect 9355 8789 9364 8823
rect 9312 8780 9364 8789
rect 16580 8780 16632 8832
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5194 8678 5246 8730
rect 5258 8678 5310 8730
rect 5322 8678 5374 8730
rect 4712 8619 4764 8628
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 5448 8576 5500 8628
rect 1768 8551 1820 8560
rect 1768 8517 1777 8551
rect 1777 8517 1811 8551
rect 1811 8517 1820 8551
rect 1768 8508 1820 8517
rect 4804 8508 4856 8560
rect 6828 8576 6880 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 9312 8508 9364 8560
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 2872 8440 2924 8492
rect 6092 8440 6144 8492
rect 8208 8440 8260 8492
rect 8760 8440 8812 8492
rect 9404 8440 9456 8492
rect 3792 8304 3844 8356
rect 4436 8304 4488 8356
rect 6460 8304 6512 8356
rect 8484 8304 8536 8356
rect 8760 8347 8812 8356
rect 8760 8313 8769 8347
rect 8769 8313 8803 8347
rect 8803 8313 8812 8347
rect 8760 8304 8812 8313
rect 16580 8304 16632 8356
rect 3148 8236 3200 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 2964 8032 3016 8084
rect 4804 7964 4856 8016
rect 4620 7896 4672 7948
rect 5908 7896 5960 7948
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 3332 7760 3384 7812
rect 4896 7828 4948 7880
rect 6460 7871 6512 7880
rect 3884 7803 3936 7812
rect 3884 7769 3893 7803
rect 3893 7769 3927 7803
rect 3927 7769 3936 7803
rect 3884 7760 3936 7769
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 8760 7896 8812 7948
rect 9312 8032 9364 8084
rect 9496 7964 9548 8016
rect 9128 7896 9180 7948
rect 8024 7760 8076 7812
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 8852 7735 8904 7744
rect 8852 7701 8861 7735
rect 8861 7701 8895 7735
rect 8895 7701 8904 7735
rect 8852 7692 8904 7701
rect 16672 7760 16724 7812
rect 16580 7692 16632 7744
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 5194 7590 5246 7642
rect 5258 7590 5310 7642
rect 5322 7590 5374 7642
rect 3056 7488 3108 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 3884 7420 3936 7472
rect 7932 7463 7984 7472
rect 7932 7429 7941 7463
rect 7941 7429 7975 7463
rect 7975 7429 7984 7463
rect 7932 7420 7984 7429
rect 8024 7420 8076 7472
rect 2964 7352 3016 7404
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 4160 7352 4212 7404
rect 5632 7352 5684 7404
rect 4988 7284 5040 7336
rect 8300 7352 8352 7404
rect 6184 7327 6236 7336
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 9312 7284 9364 7336
rect 6368 7216 6420 7268
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 6460 7148 6512 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 3148 6944 3200 6996
rect 6368 6876 6420 6928
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 3056 6740 3108 6792
rect 3792 6740 3844 6792
rect 5632 6808 5684 6860
rect 8392 6851 8444 6860
rect 8392 6817 8401 6851
rect 8401 6817 8435 6851
rect 8435 6817 8444 6851
rect 8392 6808 8444 6817
rect 9128 6808 9180 6860
rect 5448 6783 5500 6792
rect 2412 6604 2464 6656
rect 3332 6672 3384 6724
rect 4252 6672 4304 6724
rect 3148 6604 3200 6656
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 7380 6740 7432 6792
rect 7472 6740 7524 6792
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 5908 6672 5960 6724
rect 8024 6672 8076 6724
rect 8576 6740 8628 6792
rect 8944 6672 8996 6724
rect 9220 6672 9272 6724
rect 9588 6672 9640 6724
rect 8208 6604 8260 6656
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5194 6502 5246 6554
rect 5258 6502 5310 6554
rect 5322 6502 5374 6554
rect 3056 6400 3108 6452
rect 7380 6400 7432 6452
rect 1584 6332 1636 6384
rect 2412 6375 2464 6384
rect 2412 6341 2421 6375
rect 2421 6341 2455 6375
rect 2455 6341 2464 6375
rect 2412 6332 2464 6341
rect 4252 6332 4304 6384
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5448 6264 5500 6316
rect 5908 6239 5960 6248
rect 5908 6205 5917 6239
rect 5917 6205 5951 6239
rect 5951 6205 5960 6239
rect 5908 6196 5960 6205
rect 6092 6264 6144 6316
rect 6736 6332 6788 6384
rect 7932 6400 7984 6452
rect 8392 6400 8444 6452
rect 9404 6400 9456 6452
rect 9496 6443 9548 6452
rect 9496 6409 9505 6443
rect 9505 6409 9539 6443
rect 9539 6409 9548 6443
rect 9496 6400 9548 6409
rect 16580 6400 16632 6452
rect 8852 6332 8904 6384
rect 9128 6375 9180 6384
rect 9128 6341 9137 6375
rect 9137 6341 9171 6375
rect 9171 6341 9180 6375
rect 9128 6332 9180 6341
rect 8208 6264 8260 6316
rect 8392 6264 8444 6316
rect 8576 6264 8628 6316
rect 8024 6196 8076 6248
rect 8300 6196 8352 6248
rect 19432 6128 19484 6180
rect 4988 6060 5040 6112
rect 5448 6060 5500 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 1584 5856 1636 5908
rect 3148 5856 3200 5908
rect 4620 5856 4672 5908
rect 5908 5899 5960 5908
rect 5908 5865 5917 5899
rect 5917 5865 5951 5899
rect 5951 5865 5960 5899
rect 5908 5856 5960 5865
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 8116 5788 8168 5840
rect 1492 5720 1544 5772
rect 5724 5720 5776 5772
rect 6092 5720 6144 5772
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 8852 5720 8904 5772
rect 3332 5652 3384 5704
rect 3424 5516 3476 5568
rect 3792 5584 3844 5636
rect 4896 5584 4948 5636
rect 8208 5584 8260 5636
rect 8944 5627 8996 5636
rect 8944 5593 8953 5627
rect 8953 5593 8987 5627
rect 8987 5593 8996 5627
rect 9496 5627 9548 5636
rect 8944 5584 8996 5593
rect 9496 5593 9505 5627
rect 9505 5593 9539 5627
rect 9539 5593 9548 5627
rect 9496 5584 9548 5593
rect 9128 5516 9180 5568
rect 13820 5584 13872 5636
rect 16672 5584 16724 5636
rect 16580 5516 16632 5568
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5194 5414 5246 5466
rect 5258 5414 5310 5466
rect 5322 5414 5374 5466
rect 3884 5312 3936 5364
rect 7012 5312 7064 5364
rect 4896 5244 4948 5296
rect 8208 5244 8260 5296
rect 8484 5244 8536 5296
rect 1492 5176 1544 5228
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 8760 5176 8812 5228
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 5172 5108 5224 5160
rect 6920 5108 6972 5160
rect 5080 5015 5132 5024
rect 5080 4981 5089 5015
rect 5089 4981 5123 5015
rect 5123 4981 5132 5015
rect 5080 4972 5132 4981
rect 8392 4972 8444 5024
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 5724 4811 5776 4820
rect 5724 4777 5733 4811
rect 5733 4777 5767 4811
rect 5767 4777 5776 4811
rect 5724 4768 5776 4777
rect 9220 4768 9272 4820
rect 5080 4700 5132 4752
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 4160 4632 4212 4684
rect 4988 4564 5040 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7012 4564 7064 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 9128 4564 9180 4616
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 4896 4496 4948 4548
rect 5540 4496 5592 4548
rect 7472 4496 7524 4548
rect 4344 4428 4396 4480
rect 5172 4428 5224 4480
rect 8944 4471 8996 4480
rect 8944 4437 8961 4471
rect 8961 4437 8995 4471
rect 8995 4437 8996 4471
rect 9220 4471 9272 4480
rect 8944 4428 8996 4437
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 5194 4326 5246 4378
rect 5258 4326 5310 4378
rect 5322 4326 5374 4378
rect 6552 4224 6604 4276
rect 8760 4224 8812 4276
rect 5816 4156 5868 4208
rect 3240 4088 3292 4140
rect 5356 4131 5408 4140
rect 3884 4063 3936 4072
rect 3884 4029 3893 4063
rect 3893 4029 3927 4063
rect 3927 4029 3936 4063
rect 3884 4020 3936 4029
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5448 4088 5500 4140
rect 9220 4088 9272 4140
rect 9588 4088 9640 4140
rect 4160 4020 4212 4072
rect 2688 3952 2740 4004
rect 6920 4020 6972 4072
rect 8852 4063 8904 4072
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 13820 3952 13872 4004
rect 5908 3927 5960 3936
rect 5908 3893 5925 3927
rect 5925 3893 5959 3927
rect 5959 3893 5960 3927
rect 5908 3884 5960 3893
rect 6552 3884 6604 3936
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 5356 3680 5408 3732
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 9588 3680 9640 3732
rect 3332 3544 3384 3596
rect 6920 3544 6972 3596
rect 4804 3476 4856 3528
rect 4436 3408 4488 3460
rect 5540 3408 5592 3460
rect 6644 3476 6696 3528
rect 7012 3476 7064 3528
rect 8484 3476 8536 3528
rect 6460 3408 6512 3460
rect 6552 3451 6604 3460
rect 6552 3417 6561 3451
rect 6561 3417 6595 3451
rect 6595 3417 6604 3451
rect 6552 3408 6604 3417
rect 7932 3408 7984 3460
rect 8944 3340 8996 3392
rect 16580 3340 16632 3392
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5194 3238 5246 3290
rect 5258 3238 5310 3290
rect 5322 3238 5374 3290
rect 4344 3136 4396 3188
rect 4436 3136 4488 3188
rect 6092 3068 6144 3120
rect 7472 3111 7524 3120
rect 7472 3077 7481 3111
rect 7481 3077 7515 3111
rect 7515 3077 7524 3111
rect 7472 3068 7524 3077
rect 4896 3000 4948 3052
rect 6460 3043 6512 3052
rect 6460 3009 6469 3043
rect 6469 3009 6503 3043
rect 6503 3009 6512 3043
rect 6460 3000 6512 3009
rect 6552 3000 6604 3052
rect 8392 3136 8444 3188
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 9036 3136 9088 3188
rect 8116 3111 8168 3120
rect 8116 3077 8125 3111
rect 8125 3077 8159 3111
rect 8159 3077 8168 3111
rect 8116 3068 8168 3077
rect 8760 3068 8812 3120
rect 9312 3000 9364 3052
rect 3424 2932 3476 2984
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 5632 2932 5684 2984
rect 9220 2932 9272 2984
rect 8208 2864 8260 2916
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 4620 2592 4672 2644
rect 6092 2635 6144 2644
rect 6092 2601 6101 2635
rect 6101 2601 6135 2635
rect 6135 2601 6144 2635
rect 6092 2592 6144 2601
rect 6736 2592 6788 2644
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 7932 2635 7984 2644
rect 4436 2524 4488 2576
rect 3240 2320 3292 2372
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 5448 2456 5500 2508
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 4068 2320 4120 2372
rect 4988 2320 5040 2372
rect 6552 2524 6604 2576
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 9220 2635 9272 2644
rect 9220 2601 9229 2635
rect 9229 2601 9263 2635
rect 9263 2601 9272 2635
rect 9220 2592 9272 2601
rect 8116 2524 8168 2576
rect 8484 2567 8536 2576
rect 8484 2533 8493 2567
rect 8493 2533 8527 2567
rect 8527 2533 8536 2567
rect 8484 2524 8536 2533
rect 9128 2524 9180 2576
rect 6000 2320 6052 2372
rect 6736 2320 6788 2372
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 8300 2363 8352 2372
rect 8300 2329 8309 2363
rect 8309 2329 8343 2363
rect 8343 2329 8352 2363
rect 8300 2320 8352 2329
rect 9588 2320 9640 2372
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 5194 2150 5246 2202
rect 5258 2150 5310 2202
rect 5322 2150 5374 2202
rect 4344 2048 4396 2100
rect 6828 2048 6880 2100
rect 8300 2091 8352 2100
rect 8300 2057 8309 2091
rect 8309 2057 8343 2091
rect 8343 2057 8352 2091
rect 8300 2048 8352 2057
rect 8668 2048 8720 2100
rect 9312 2091 9364 2100
rect 9312 2057 9321 2091
rect 9321 2057 9355 2091
rect 9355 2057 9364 2091
rect 9312 2048 9364 2057
rect 4068 1980 4120 2032
rect 6000 2023 6052 2032
rect 6000 1989 6009 2023
rect 6009 1989 6043 2023
rect 6043 1989 6052 2023
rect 6000 1980 6052 1989
rect 6276 1980 6328 2032
rect 7840 1980 7892 2032
rect 9128 1980 9180 2032
rect 4988 1912 5040 1964
rect 4252 1844 4304 1896
rect 9128 1887 9180 1896
rect 9128 1853 9137 1887
rect 9137 1853 9171 1887
rect 9171 1853 9180 1887
rect 9128 1844 9180 1853
rect 8944 1751 8996 1760
rect 8944 1717 8953 1751
rect 8953 1717 8987 1751
rect 8987 1717 8996 1751
rect 8944 1708 8996 1717
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 4160 1504 4212 1556
rect 9588 1504 9640 1556
rect 5448 1436 5500 1488
rect 6184 1300 6236 1352
rect 4896 1164 4948 1216
rect 5066 1062 5118 1114
rect 5130 1062 5182 1114
rect 5194 1062 5246 1114
rect 5258 1062 5310 1114
rect 5322 1062 5374 1114
<< obsm1 >>
rect 24000 0 34000 13000
<< metal2 >>
rect 938 12322 994 13000
rect 1398 12322 1454 13000
rect 938 12294 1256 12322
rect 938 12200 994 12294
rect 1228 11286 1256 12294
rect 1398 12294 1808 12322
rect 1398 12200 1454 12294
rect 1780 11354 1808 12294
rect 1858 12200 1914 13000
rect 2318 12322 2374 13000
rect 2318 12294 2452 12322
rect 2318 12200 2374 12294
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1216 11280 1268 11286
rect 1216 11222 1268 11228
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 9722 1532 9998
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 1504 8498 1532 9658
rect 1596 9518 1624 10542
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1780 8566 1808 10406
rect 1872 9738 1900 12200
rect 2320 9988 2372 9994
rect 2320 9930 2372 9936
rect 1872 9710 1992 9738
rect 1964 9625 1992 9710
rect 2332 9654 2360 9930
rect 2320 9648 2372 9654
rect 1950 9616 2006 9625
rect 2320 9590 2372 9596
rect 1950 9551 2006 9560
rect 1964 9178 1992 9551
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2332 8974 2360 9590
rect 2424 9178 2452 12294
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12322 4214 13000
rect 4158 12294 4476 12322
rect 4158 12200 4214 12294
rect 2792 11642 2820 12200
rect 2792 11614 3096 11642
rect 2566 11452 2874 11461
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11387 2874 11396
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2976 10674 3004 10950
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2566 10364 2874 10373
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10299 2874 10308
rect 2566 9276 2874 9285
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9211 2874 9220
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 2884 8498 2912 8910
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 1504 6866 1532 8434
rect 2566 8188 2874 8197
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8123 2874 8132
rect 2976 8090 3004 9114
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 7410 3004 7686
rect 3068 7546 3096 11614
rect 3146 9616 3202 9625
rect 3146 9551 3202 9560
rect 3160 8906 3188 9551
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2566 7100 2874 7109
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7035 2874 7044
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 5778 1532 6802
rect 3068 6798 3096 7482
rect 3160 7410 3188 8230
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 7002 3188 7346
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 6390 2452 6598
rect 3068 6458 3096 6734
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 1584 6384 1636 6390
rect 1584 6326 1636 6332
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 1596 5914 1624 6326
rect 3160 6322 3188 6598
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2566 6012 2874 6021
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5947 2874 5956
rect 3160 5914 3188 6258
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1504 5234 1532 5714
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 3252 4146 3280 12200
rect 3712 10010 3740 12200
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4356 11150 4384 11290
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 3712 9982 3832 10010
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3712 9518 3740 9862
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3620 8974 3648 9114
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 7886 3648 8910
rect 3804 8362 3832 9982
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9518 4200 9862
rect 4264 9654 4292 11018
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3344 6730 3372 7754
rect 3896 7478 3924 7754
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 4172 7410 4200 9114
rect 4356 9110 4384 10610
rect 4448 9382 4476 12294
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 9218 12336 9274 12345
rect 9218 12271 9274 12280
rect 4632 11370 4660 12200
rect 4632 11342 4844 11370
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4540 10266 4568 10678
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4632 10130 4660 10950
rect 4724 10742 4752 11154
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5234 3372 5646
rect 3804 5642 3832 6734
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4264 6390 4292 6666
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3344 4690 3372 5170
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2700 3437 2728 3946
rect 2686 3428 2742 3437
rect 2686 3363 2742 3372
rect 3252 2378 3280 4082
rect 3344 3602 3372 4626
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3436 2990 3464 5510
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3896 4078 3924 5306
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4172 4078 4200 4626
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4356 3194 4384 4422
rect 4448 3466 4476 8298
rect 4540 5137 4568 9658
rect 4632 9625 4660 10066
rect 4724 10062 4752 10678
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4618 9616 4674 9625
rect 4618 9551 4674 9560
rect 4724 8634 4752 9998
rect 4816 8650 4844 11342
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5000 10674 5028 11086
rect 5092 10996 5120 12200
rect 5552 11218 5580 12200
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5540 11008 5592 11014
rect 5092 10968 5488 10996
rect 5066 10908 5374 10917
rect 5066 10906 5072 10908
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5368 10906 5374 10908
rect 5128 10854 5130 10906
rect 5310 10854 5312 10906
rect 5066 10852 5072 10854
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5368 10852 5374 10854
rect 5066 10843 5374 10852
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 9722 4936 10406
rect 5066 9820 5374 9829
rect 5066 9818 5072 9820
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5368 9818 5374 9820
rect 5128 9766 5130 9818
rect 5310 9766 5312 9818
rect 5066 9764 5072 9766
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5368 9764 5374 9766
rect 5066 9755 5374 9764
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5066 8732 5374 8741
rect 5066 8730 5072 8732
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5368 8730 5374 8732
rect 5128 8678 5130 8730
rect 5310 8678 5312 8730
rect 5066 8676 5072 8678
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5368 8676 5374 8678
rect 5066 8667 5374 8676
rect 4712 8628 4764 8634
rect 4816 8622 5028 8650
rect 5460 8634 5488 10968
rect 5540 10950 5592 10956
rect 5552 10130 5580 10950
rect 5644 10606 5672 11018
rect 6012 10810 6040 12200
rect 6472 11354 6500 12200
rect 7566 11452 7874 11461
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11387 7874 11396
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5644 9586 5672 10406
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5828 9722 5856 9998
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 4712 8570 4764 8576
rect 4724 7970 4752 8570
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4816 8022 4844 8502
rect 4632 7954 4752 7970
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4620 7948 4752 7954
rect 4672 7942 4752 7948
rect 4620 7890 4672 7896
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4632 5914 4660 6258
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4526 5128 4582 5137
rect 4526 5063 4582 5072
rect 4816 3534 4844 7958
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4908 5642 4936 7822
rect 5000 7342 5028 8622
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5066 7644 5374 7653
rect 5066 7642 5072 7644
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5368 7642 5374 7644
rect 5128 7590 5130 7642
rect 5310 7590 5312 7642
rect 5066 7588 5072 7590
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5368 7588 5374 7590
rect 5066 7579 5374 7588
rect 5644 7410 5672 8842
rect 5920 7954 5948 10406
rect 6012 10266 6040 10406
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6012 9654 6040 10202
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 6012 8906 6040 9590
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6104 8378 6132 8434
rect 6104 8350 6224 8378
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5644 6866 5672 7346
rect 6196 7342 6224 8350
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5066 6556 5374 6565
rect 5066 6554 5072 6556
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5368 6554 5374 6556
rect 5128 6502 5130 6554
rect 5310 6502 5312 6554
rect 5066 6500 5072 6502
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5368 6500 5374 6502
rect 5066 6491 5374 6500
rect 5460 6322 5488 6734
rect 5920 6730 5948 7142
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 4896 5636 4948 5642
rect 4896 5578 4948 5584
rect 4908 5302 4936 5578
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4908 4554 4936 5238
rect 5000 4622 5028 6054
rect 5066 5468 5374 5477
rect 5066 5466 5072 5468
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5368 5466 5374 5468
rect 5128 5414 5130 5466
rect 5310 5414 5312 5466
rect 5066 5412 5072 5414
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5368 5412 5374 5414
rect 5066 5403 5374 5412
rect 5460 5409 5488 6054
rect 5920 5914 5948 6190
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6104 5778 6132 6258
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 5446 5400 5502 5409
rect 5446 5335 5502 5344
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5092 4758 5120 4966
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4448 3194 4476 3402
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4356 3074 4384 3130
rect 4264 3046 4384 3074
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4080 2038 4108 2314
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 4172 1562 4200 2382
rect 4264 1902 4292 3046
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2106 4384 2790
rect 4448 2582 4476 3130
rect 5000 3074 5028 4558
rect 5184 4486 5212 5102
rect 5736 4826 5764 5714
rect 6104 5658 6132 5714
rect 6012 5630 6132 5658
rect 6012 5234 6040 5630
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5066 4380 5374 4389
rect 5066 4378 5072 4380
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5368 4378 5374 4380
rect 5128 4326 5130 4378
rect 5310 4326 5312 4378
rect 5066 4324 5072 4326
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5368 4324 5374 4326
rect 5066 4315 5374 4324
rect 5460 4146 5488 4558
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5368 3738 5396 4082
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5552 3466 5580 4490
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5066 3292 5374 3301
rect 5066 3290 5072 3292
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5368 3290 5374 3292
rect 5128 3238 5130 3290
rect 5310 3238 5312 3290
rect 5066 3236 5072 3238
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5368 3236 5374 3238
rect 5066 3227 5374 3236
rect 5736 3074 5764 4762
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5828 3738 5856 4150
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5920 3369 5948 3878
rect 5906 3360 5962 3369
rect 5906 3295 5962 3304
rect 4908 3058 5028 3074
rect 4896 3052 5028 3058
rect 4948 3046 5028 3052
rect 5644 3046 5764 3074
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 4896 2994 4948 3000
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4632 2650 4660 2926
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 4908 2446 4936 2994
rect 5644 2990 5672 3046
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 6104 2650 6132 3062
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4344 2100 4396 2106
rect 4344 2042 4396 2048
rect 4252 1896 4304 1902
rect 4252 1838 4304 1844
rect 4160 1556 4212 1562
rect 4160 1498 4212 1504
rect 4908 1222 4936 2382
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 5000 1970 5028 2314
rect 5066 2204 5374 2213
rect 5066 2202 5072 2204
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5368 2202 5374 2204
rect 5128 2150 5130 2202
rect 5310 2150 5312 2202
rect 5066 2148 5072 2150
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5368 2148 5374 2150
rect 5066 2139 5374 2148
rect 4988 1964 5040 1970
rect 4988 1906 5040 1912
rect 5460 1494 5488 2450
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 6012 2038 6040 2314
rect 6000 2032 6052 2038
rect 6000 1974 6052 1980
rect 5448 1488 5500 1494
rect 5448 1430 5500 1436
rect 6196 1358 6224 7278
rect 6288 2038 6316 11154
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 9994 6408 10406
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6472 8362 6500 10746
rect 6564 10674 6592 11222
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6380 6934 6408 7210
rect 6472 7206 6500 7822
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6472 5778 6500 7142
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4282 6592 4558
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6564 3466 6592 3878
rect 6656 3534 6684 9318
rect 6748 9178 6776 9454
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6840 9042 6868 11086
rect 7300 11014 7328 11154
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10606 7328 10950
rect 7484 10674 7512 11018
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10674 7696 10950
rect 7930 10704 7986 10713
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7656 10668 7708 10674
rect 7930 10639 7986 10648
rect 7656 10610 7708 10616
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7116 10062 7144 10406
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7208 9586 7236 10406
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8634 6868 8978
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6840 7970 6868 8570
rect 6748 7942 6868 7970
rect 6748 6390 6776 7942
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 7024 5370 7052 8842
rect 7484 6798 7512 10610
rect 7566 10364 7874 10373
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10299 7874 10308
rect 7566 9276 7874 9285
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9211 7874 9220
rect 7566 8188 7874 8197
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8123 7874 8132
rect 7944 7478 7972 10639
rect 8128 10062 8156 11290
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 8634 8064 9454
rect 8220 9178 8248 10678
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8312 9654 8340 9930
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8864 9586 8892 9930
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8220 8498 8248 9114
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8036 7478 8064 7754
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8206 7440 8262 7449
rect 7566 7100 7874 7109
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7035 7874 7044
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7392 6458 7420 6734
rect 7944 6458 7972 7414
rect 8206 7375 8262 7384
rect 8300 7404 8352 7410
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8036 6254 8064 6666
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 7566 6012 7874 6021
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5947 7874 5956
rect 8128 5846 8156 6734
rect 8220 6662 8248 7375
rect 8300 7346 8352 7352
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8220 5914 8248 6258
rect 8312 6254 8340 7346
rect 8404 6866 8432 9318
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8404 6458 8432 6802
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8390 6352 8446 6361
rect 8390 6287 8392 6296
rect 8444 6287 8446 6296
rect 8392 6258 8444 6264
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8220 5642 8248 5850
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6932 4078 6960 5102
rect 7024 4622 7052 5306
rect 8220 5302 8248 5578
rect 8496 5302 8524 8298
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 6798 8616 7278
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8588 5914 8616 6258
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 7566 4924 7874 4933
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4859 7874 4868
rect 8404 4622 8432 4966
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6932 3602 6960 4014
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6472 3058 6500 3402
rect 6564 3058 6592 3402
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6564 2582 6592 2994
rect 6656 2774 6684 3470
rect 6656 2746 6776 2774
rect 6748 2650 6776 2746
rect 7024 2650 7052 3470
rect 7484 3126 7512 4490
rect 7566 3836 7874 3845
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3771 7874 3780
rect 8496 3618 8524 5238
rect 8680 4593 8708 9318
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8772 8498 8800 8842
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8772 7954 8800 8298
rect 9140 7954 9168 9862
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8864 6390 8892 7686
rect 9140 6866 9168 7890
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8666 4584 8722 4593
rect 8666 4519 8722 4528
rect 8404 3590 8524 3618
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7566 2748 7874 2757
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2683 7874 2692
rect 7944 2650 7972 3402
rect 8404 3194 8432 3590
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6748 2378 6776 2586
rect 8128 2582 8156 3062
rect 8206 2952 8262 2961
rect 8206 2887 8208 2896
rect 8260 2887 8262 2896
rect 8208 2858 8260 2864
rect 8496 2582 8524 3470
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8680 2446 8708 4519
rect 8772 4282 8800 5170
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8772 3126 8800 4218
rect 8864 4078 8892 5714
rect 8956 5642 8984 6666
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4185 8984 4422
rect 8942 4176 8998 4185
rect 8942 4111 8998 4120
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8956 3482 8984 4111
rect 8864 3454 8984 3482
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8864 2774 8892 3454
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3194 8984 3334
rect 9048 3194 9076 6598
rect 9140 6390 9168 6802
rect 9232 6730 9260 12271
rect 9494 11928 9550 11937
rect 9494 11863 9550 11872
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9416 9926 9444 10610
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9324 8566 9352 8774
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9324 8090 9352 8502
rect 9416 8498 9444 9862
rect 9508 9178 9536 11863
rect 16854 11520 16910 11529
rect 16854 11455 16910 11464
rect 16578 11112 16634 11121
rect 16578 11047 16580 11056
rect 16632 11047 16634 11056
rect 16580 11018 16632 11024
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16592 10305 16620 10406
rect 16578 10296 16634 10305
rect 16578 10231 16634 10240
rect 16762 9888 16818 9897
rect 16762 9823 16818 9832
rect 16578 9480 16634 9489
rect 16578 9415 16634 9424
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 8265 9444 8434
rect 9402 8256 9458 8265
rect 9402 8191 9458 8200
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9324 7342 9352 8026
rect 9416 7546 9444 8191
rect 9508 8022 9536 9114
rect 16592 8838 16620 9415
rect 16670 9072 16726 9081
rect 16776 9042 16804 9823
rect 16670 9007 16726 9016
rect 16764 9036 16816 9042
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16578 8664 16634 8673
rect 16578 8599 16634 8608
rect 16592 8362 16620 8599
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 16578 7848 16634 7857
rect 16684 7818 16712 9007
rect 16764 8978 16816 8984
rect 16578 7783 16634 7792
rect 16672 7812 16724 7818
rect 16592 7750 16620 7783
rect 16672 7754 16724 7760
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 9404 7540 9456 7546
rect 9456 7500 9536 7528
rect 9404 7482 9456 7488
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9508 6458 9536 7500
rect 16868 6914 16896 11455
rect 19430 7032 19486 7041
rect 19430 6967 19486 6976
rect 16684 6886 16896 6914
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9126 5808 9182 5817
rect 9126 5743 9182 5752
rect 9140 5574 9168 5743
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9140 4622 9168 5510
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9232 4826 9260 5170
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9232 4146 9260 4422
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9324 3210 9352 4558
rect 9416 3738 9444 6394
rect 9508 6361 9536 6394
rect 9494 6352 9550 6361
rect 9494 6287 9550 6296
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9232 3182 9352 3210
rect 9232 3074 9260 3182
rect 9140 3046 9260 3074
rect 9312 3052 9364 3058
rect 8864 2746 9076 2774
rect 9048 2650 9076 2746
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9140 2582 9168 3046
rect 9312 2994 9364 3000
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9232 2650 9260 2926
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 7840 2440 7892 2446
rect 6826 2408 6882 2417
rect 6736 2372 6788 2378
rect 7840 2382 7892 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 6826 2343 6882 2352
rect 6736 2314 6788 2320
rect 6840 2106 6868 2343
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 7852 2038 7880 2382
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8312 2106 8340 2314
rect 8680 2106 8708 2382
rect 8300 2100 8352 2106
rect 8300 2042 8352 2048
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 9140 2038 9168 2518
rect 9324 2145 9352 2994
rect 9310 2136 9366 2145
rect 9310 2071 9312 2080
rect 9364 2071 9366 2080
rect 9312 2042 9364 2048
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 7840 2032 7892 2038
rect 7840 1974 7892 1980
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 8944 1760 8996 1766
rect 8944 1702 8996 1708
rect 7566 1660 7874 1669
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1595 7874 1604
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 4896 1216 4948 1222
rect 4896 1158 4948 1164
rect 5066 1116 5374 1125
rect 5066 1114 5072 1116
rect 5128 1114 5152 1116
rect 5208 1114 5232 1116
rect 5288 1114 5312 1116
rect 5368 1114 5374 1116
rect 5128 1062 5130 1114
rect 5310 1062 5312 1114
rect 5066 1060 5072 1062
rect 5128 1060 5152 1062
rect 5208 1060 5232 1062
rect 5288 1060 5312 1062
rect 5368 1060 5374 1062
rect 5066 1051 5374 1060
rect 8956 513 8984 1702
rect 9140 1329 9168 1838
rect 9126 1320 9182 1329
rect 9126 1255 9182 1264
rect 9508 921 9536 5578
rect 9600 4146 9628 6666
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16592 6458 16620 6559
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16578 6216 16634 6225
rect 16578 6151 16634 6160
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 13832 4010 13860 5578
rect 16592 5574 16620 6151
rect 16684 5642 16712 6886
rect 19444 6186 19472 6967
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 16578 3768 16634 3777
rect 9588 3732 9640 3738
rect 16578 3703 16634 3712
rect 9588 3674 9640 3680
rect 9600 2378 9628 3674
rect 16592 3398 16620 3703
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 9600 1737 9628 2314
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 9600 1562 9628 1663
rect 9588 1556 9640 1562
rect 9588 1498 9640 1504
rect 9494 912 9550 921
rect 9494 847 9550 856
rect 8942 504 8998 513
rect 8942 439 8998 448
<< via2 >>
rect 1950 9560 2006 9616
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 3146 9560 3202 9616
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 9218 12280 9274 12336
rect 2686 3372 2742 3428
rect 4618 9560 4674 9616
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5118 10906
rect 5118 10854 5128 10906
rect 5152 10854 5182 10906
rect 5182 10854 5194 10906
rect 5194 10854 5208 10906
rect 5232 10854 5246 10906
rect 5246 10854 5258 10906
rect 5258 10854 5288 10906
rect 5312 10854 5322 10906
rect 5322 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5118 9818
rect 5118 9766 5128 9818
rect 5152 9766 5182 9818
rect 5182 9766 5194 9818
rect 5194 9766 5208 9818
rect 5232 9766 5246 9818
rect 5246 9766 5258 9818
rect 5258 9766 5288 9818
rect 5312 9766 5322 9818
rect 5322 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5118 8730
rect 5118 8678 5128 8730
rect 5152 8678 5182 8730
rect 5182 8678 5194 8730
rect 5194 8678 5208 8730
rect 5232 8678 5246 8730
rect 5246 8678 5258 8730
rect 5258 8678 5288 8730
rect 5312 8678 5322 8730
rect 5322 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 4526 5072 4582 5128
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5118 7642
rect 5118 7590 5128 7642
rect 5152 7590 5182 7642
rect 5182 7590 5194 7642
rect 5194 7590 5208 7642
rect 5232 7590 5246 7642
rect 5246 7590 5258 7642
rect 5258 7590 5288 7642
rect 5312 7590 5322 7642
rect 5322 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5118 6554
rect 5118 6502 5128 6554
rect 5152 6502 5182 6554
rect 5182 6502 5194 6554
rect 5194 6502 5208 6554
rect 5232 6502 5246 6554
rect 5246 6502 5258 6554
rect 5258 6502 5288 6554
rect 5312 6502 5322 6554
rect 5322 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5118 5466
rect 5118 5414 5128 5466
rect 5152 5414 5182 5466
rect 5182 5414 5194 5466
rect 5194 5414 5208 5466
rect 5232 5414 5246 5466
rect 5246 5414 5258 5466
rect 5258 5414 5288 5466
rect 5312 5414 5322 5466
rect 5322 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 5446 5344 5502 5400
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5118 4378
rect 5118 4326 5128 4378
rect 5152 4326 5182 4378
rect 5182 4326 5194 4378
rect 5194 4326 5208 4378
rect 5232 4326 5246 4378
rect 5246 4326 5258 4378
rect 5258 4326 5288 4378
rect 5312 4326 5322 4378
rect 5322 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5118 3290
rect 5118 3238 5128 3290
rect 5152 3238 5182 3290
rect 5182 3238 5194 3290
rect 5194 3238 5208 3290
rect 5232 3238 5246 3290
rect 5246 3238 5258 3290
rect 5258 3238 5288 3290
rect 5312 3238 5322 3290
rect 5322 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 5906 3304 5962 3360
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5118 2202
rect 5118 2150 5128 2202
rect 5152 2150 5182 2202
rect 5182 2150 5194 2202
rect 5194 2150 5208 2202
rect 5232 2150 5246 2202
rect 5246 2150 5258 2202
rect 5258 2150 5288 2202
rect 5312 2150 5322 2202
rect 5322 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 7930 10648 7986 10704
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 8206 7384 8262 7440
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 8390 6316 8446 6352
rect 8390 6296 8392 6316
rect 8392 6296 8444 6316
rect 8444 6296 8446 6316
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 8666 4528 8722 4584
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 8206 2916 8262 2952
rect 8206 2896 8208 2916
rect 8208 2896 8260 2916
rect 8260 2896 8262 2916
rect 8942 4120 8998 4176
rect 9494 11872 9550 11928
rect 16854 11464 16910 11520
rect 16578 11076 16634 11112
rect 16578 11056 16580 11076
rect 16580 11056 16632 11076
rect 16632 11056 16634 11076
rect 16578 10240 16634 10296
rect 16762 9832 16818 9888
rect 16578 9424 16634 9480
rect 9402 8200 9458 8256
rect 16670 9016 16726 9072
rect 16578 8608 16634 8664
rect 16578 7792 16634 7848
rect 19430 6976 19486 7032
rect 9126 5752 9182 5808
rect 9494 6296 9550 6352
rect 6826 2352 6882 2408
rect 9310 2100 9366 2136
rect 9310 2080 9312 2100
rect 9312 2080 9364 2100
rect 9364 2080 9366 2100
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 5072 1114 5128 1116
rect 5152 1114 5208 1116
rect 5232 1114 5288 1116
rect 5312 1114 5368 1116
rect 5072 1062 5118 1114
rect 5118 1062 5128 1114
rect 5152 1062 5182 1114
rect 5182 1062 5194 1114
rect 5194 1062 5208 1114
rect 5232 1062 5246 1114
rect 5246 1062 5258 1114
rect 5258 1062 5288 1114
rect 5312 1062 5322 1114
rect 5322 1062 5368 1114
rect 5072 1060 5128 1062
rect 5152 1060 5208 1062
rect 5232 1060 5288 1062
rect 5312 1060 5368 1062
rect 9126 1264 9182 1320
rect 16578 6568 16634 6624
rect 16578 6160 16634 6216
rect 16578 3712 16634 3768
rect 9586 1672 9642 1728
rect 9494 856 9550 912
rect 8942 448 8998 504
<< obsm2 >>
rect 24000 0 34000 13000
<< metal3 >>
rect 9213 12338 9279 12341
rect 14000 12338 34000 12368
rect 9213 12336 34000 12338
rect 9213 12280 9218 12336
rect 9274 12280 34000 12336
rect 9213 12278 34000 12280
rect 9213 12275 9279 12278
rect 14000 12248 34000 12278
rect 9489 11930 9555 11933
rect 14000 11930 34000 11960
rect 9489 11928 34000 11930
rect 9489 11872 9494 11928
rect 9550 11872 34000 11928
rect 9489 11870 34000 11872
rect 9489 11867 9555 11870
rect 14000 11840 34000 11870
rect 14000 11520 34000 11552
rect 14000 11464 16854 11520
rect 16910 11464 34000 11520
rect 2562 11456 2878 11457
rect 2562 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2878 11456
rect 2562 11391 2878 11392
rect 7562 11456 7878 11457
rect 7562 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7878 11456
rect 14000 11432 34000 11464
rect 7562 11391 7878 11392
rect 14000 11112 34000 11144
rect 14000 11056 16578 11112
rect 16634 11056 34000 11112
rect 14000 11024 34000 11056
rect 5062 10912 5378 10913
rect 5062 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5378 10912
rect 5062 10847 5378 10848
rect 7925 10706 7991 10709
rect 14000 10706 34000 10736
rect 7925 10704 34000 10706
rect 7925 10648 7930 10704
rect 7986 10648 34000 10704
rect 7925 10646 34000 10648
rect 7925 10643 7991 10646
rect 14000 10616 34000 10646
rect 2562 10368 2878 10369
rect 2562 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2878 10368
rect 2562 10303 2878 10304
rect 7562 10368 7878 10369
rect 7562 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7878 10368
rect 7562 10303 7878 10304
rect 14000 10296 34000 10328
rect 14000 10240 16578 10296
rect 16634 10240 34000 10296
rect 14000 10208 34000 10240
rect 14000 9888 34000 9920
rect 14000 9832 16762 9888
rect 16818 9832 34000 9888
rect 5062 9824 5378 9825
rect 5062 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5378 9824
rect 14000 9800 34000 9832
rect 5062 9759 5378 9760
rect 1945 9618 2011 9621
rect 3141 9618 3207 9621
rect 4613 9618 4679 9621
rect 1945 9616 4679 9618
rect 1945 9560 1950 9616
rect 2006 9560 3146 9616
rect 3202 9560 4618 9616
rect 4674 9560 4679 9616
rect 1945 9558 4679 9560
rect 1945 9555 2011 9558
rect 3141 9555 3207 9558
rect 4613 9555 4679 9558
rect 14000 9480 34000 9512
rect 14000 9424 16578 9480
rect 16634 9424 34000 9480
rect 14000 9392 34000 9424
rect 2562 9280 2878 9281
rect 2562 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2878 9280
rect 2562 9215 2878 9216
rect 7562 9280 7878 9281
rect 7562 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7878 9280
rect 7562 9215 7878 9216
rect 14000 9072 34000 9104
rect 14000 9016 16670 9072
rect 16726 9016 34000 9072
rect 14000 8984 34000 9016
rect 5062 8736 5378 8737
rect 5062 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5378 8736
rect 5062 8671 5378 8672
rect 14000 8664 34000 8696
rect 14000 8608 16578 8664
rect 16634 8608 34000 8664
rect 14000 8576 34000 8608
rect 9397 8258 9463 8261
rect 14000 8258 34000 8288
rect 9397 8256 34000 8258
rect 9397 8200 9402 8256
rect 9458 8200 34000 8256
rect 9397 8198 34000 8200
rect 9397 8195 9463 8198
rect 2562 8192 2878 8193
rect 2562 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2878 8192
rect 2562 8127 2878 8128
rect 7562 8192 7878 8193
rect 7562 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7878 8192
rect 14000 8168 34000 8198
rect 7562 8127 7878 8128
rect 14000 7848 34000 7880
rect 14000 7792 16578 7848
rect 16634 7792 34000 7848
rect 14000 7760 34000 7792
rect 5062 7648 5378 7649
rect 5062 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5378 7648
rect 5062 7583 5378 7584
rect 8201 7442 8267 7445
rect 14000 7442 34000 7472
rect 8201 7440 34000 7442
rect 8201 7384 8206 7440
rect 8262 7384 34000 7440
rect 8201 7382 34000 7384
rect 8201 7379 8267 7382
rect 14000 7352 34000 7382
rect 2562 7104 2878 7105
rect 2562 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2878 7104
rect 2562 7039 2878 7040
rect 7562 7104 7878 7105
rect 7562 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7878 7104
rect 7562 7039 7878 7040
rect 14000 7032 34000 7064
rect 14000 6976 19430 7032
rect 19486 6976 34000 7032
rect 14000 6944 34000 6976
rect 14000 6624 34000 6656
rect 14000 6568 16578 6624
rect 16634 6568 34000 6624
rect 5062 6560 5378 6561
rect 5062 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5378 6560
rect 14000 6536 34000 6568
rect 5062 6495 5378 6496
rect 8385 6354 8451 6357
rect 9489 6354 9555 6357
rect 8385 6352 9555 6354
rect 8385 6296 8390 6352
rect 8446 6296 9494 6352
rect 9550 6296 9555 6352
rect 8385 6294 9555 6296
rect 8385 6291 8451 6294
rect 9489 6291 9555 6294
rect 14000 6216 34000 6248
rect 14000 6160 16578 6216
rect 16634 6160 34000 6216
rect 14000 6128 34000 6160
rect 2562 6016 2878 6017
rect 2562 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2878 6016
rect 2562 5951 2878 5952
rect 7562 6016 7878 6017
rect 7562 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7878 6016
rect 7562 5951 7878 5952
rect 9121 5810 9187 5813
rect 14000 5810 34000 5840
rect 9121 5808 34000 5810
rect 9121 5752 9126 5808
rect 9182 5752 34000 5808
rect 9121 5750 34000 5752
rect 9121 5747 9187 5750
rect 14000 5720 34000 5750
rect 5062 5472 5378 5473
rect 5062 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5378 5472
rect 5062 5407 5378 5408
rect 5441 5402 5507 5405
rect 14000 5402 34000 5432
rect 5441 5400 34000 5402
rect 5441 5344 5446 5400
rect 5502 5344 34000 5400
rect 5441 5342 34000 5344
rect 5441 5339 5507 5342
rect 14000 5312 34000 5342
rect 4521 5130 4587 5133
rect 4521 5128 12450 5130
rect 4521 5072 4526 5128
rect 4582 5072 12450 5128
rect 4521 5070 12450 5072
rect 4521 5067 4587 5070
rect 12390 4994 12450 5070
rect 14000 4994 34000 5024
rect 12390 4934 34000 4994
rect 7562 4928 7878 4929
rect 7562 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7878 4928
rect 14000 4904 34000 4934
rect 7562 4863 7878 4864
rect 8661 4586 8727 4589
rect 14000 4586 34000 4616
rect 8661 4584 34000 4586
rect 8661 4528 8666 4584
rect 8722 4528 34000 4584
rect 8661 4526 34000 4528
rect 8661 4523 8727 4526
rect 14000 4496 34000 4526
rect 5062 4384 5378 4385
rect 5062 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5378 4384
rect 5062 4319 5378 4320
rect 8937 4178 9003 4181
rect 14000 4178 34000 4208
rect 8937 4176 34000 4178
rect 8937 4120 8942 4176
rect 8998 4120 34000 4176
rect 8937 4118 34000 4120
rect 8937 4115 9003 4118
rect 14000 4088 34000 4118
rect 7562 3840 7878 3841
rect 7562 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7878 3840
rect 7562 3775 7878 3776
rect 14000 3768 34000 3800
rect 14000 3712 16578 3768
rect 16634 3712 34000 3768
rect 14000 3680 34000 3712
rect 2681 3430 2747 3433
rect 2484 3428 2747 3430
rect 2484 3372 2686 3428
rect 2742 3372 2747 3428
rect 2484 3370 2747 3372
rect 2681 3367 2747 3370
rect 5901 3362 5967 3365
rect 14000 3362 34000 3392
rect 5901 3360 34000 3362
rect 5901 3304 5906 3360
rect 5962 3304 34000 3360
rect 5901 3302 34000 3304
rect 5901 3299 5967 3302
rect 5062 3296 5378 3297
rect 5062 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5378 3296
rect 14000 3272 34000 3302
rect 5062 3231 5378 3232
rect 8201 2954 8267 2957
rect 14000 2954 34000 2984
rect 8201 2952 34000 2954
rect 8201 2896 8206 2952
rect 8262 2896 34000 2952
rect 8201 2894 34000 2896
rect 8201 2891 8267 2894
rect 14000 2864 34000 2894
rect 7562 2752 7878 2753
rect 7562 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7878 2752
rect 7562 2687 7878 2688
rect 14000 2546 34000 2576
rect 6870 2486 34000 2546
rect 6870 2413 6930 2486
rect 14000 2456 34000 2486
rect 6821 2408 6930 2413
rect 6821 2352 6826 2408
rect 6882 2352 6930 2408
rect 6821 2350 6930 2352
rect 6821 2347 6887 2350
rect 5062 2208 5378 2209
rect 5062 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5378 2208
rect 5062 2143 5378 2144
rect 9305 2138 9371 2141
rect 14000 2138 34000 2168
rect 9305 2136 34000 2138
rect 9305 2080 9310 2136
rect 9366 2080 34000 2136
rect 9305 2078 34000 2080
rect 9305 2075 9371 2078
rect 14000 2048 34000 2078
rect 9581 1730 9647 1733
rect 14000 1730 34000 1760
rect 9581 1728 34000 1730
rect 9581 1672 9586 1728
rect 9642 1672 34000 1728
rect 9581 1670 34000 1672
rect 9581 1667 9647 1670
rect 7562 1664 7878 1665
rect 7562 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7878 1664
rect 14000 1640 34000 1670
rect 7562 1599 7878 1600
rect 9121 1322 9187 1325
rect 14000 1322 34000 1352
rect 9121 1320 34000 1322
rect 9121 1264 9126 1320
rect 9182 1264 34000 1320
rect 9121 1262 34000 1264
rect 9121 1259 9187 1262
rect 14000 1232 34000 1262
rect 5062 1120 5378 1121
rect 5062 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5378 1120
rect 5062 1055 5378 1056
rect 9489 914 9555 917
rect 14000 914 34000 944
rect 9489 912 34000 914
rect 9489 856 9494 912
rect 9550 856 34000 912
rect 9489 854 34000 856
rect 9489 851 9555 854
rect 14000 824 34000 854
rect 8937 506 9003 509
rect 14000 506 34000 536
rect 8937 504 34000 506
rect 8937 448 8942 504
rect 8998 448 34000 504
rect 8937 446 34000 448
rect 8937 443 9003 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 5068 1116 5132 1120
rect 5068 1060 5072 1116
rect 5072 1060 5128 1116
rect 5128 1060 5132 1116
rect 5068 1056 5132 1060
rect 5148 1116 5212 1120
rect 5148 1060 5152 1116
rect 5152 1060 5208 1116
rect 5208 1060 5212 1116
rect 5148 1056 5212 1060
rect 5228 1116 5292 1120
rect 5228 1060 5232 1116
rect 5232 1060 5288 1116
rect 5288 1060 5292 1116
rect 5228 1056 5292 1060
rect 5308 1116 5372 1120
rect 5308 1060 5312 1116
rect 5312 1060 5368 1116
rect 5368 1060 5372 1116
rect 5308 1056 5372 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1040 2880 1222
rect 3560 9266 3880 11472
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1040 3880 2270
rect 5060 10912 5380 11472
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 9908 5380 10848
rect 5060 9824 5102 9908
rect 5338 9824 5380 9908
rect 5060 9760 5068 9824
rect 5372 9760 5380 9824
rect 5060 9672 5102 9760
rect 5338 9672 5380 9760
rect 5060 8736 5380 9672
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 6560 5380 7584
rect 5060 6496 5068 6560
rect 5132 6528 5148 6560
rect 5212 6528 5228 6560
rect 5292 6528 5308 6560
rect 5372 6496 5380 6560
rect 5060 6292 5102 6496
rect 5338 6292 5380 6496
rect 5060 5472 5380 6292
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3296 5380 4320
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 3148 5380 3232
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2208 5380 2912
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1120 5380 2144
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 5060 1040 5380 1056
rect 6060 10956 6380 11472
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 1040 6380 3960
rect 7560 11456 7880 11472
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 8218 7880 9216
rect 7560 8192 7602 8218
rect 7838 8192 7880 8218
rect 7560 8128 7568 8192
rect 7872 8128 7880 8192
rect 7560 7982 7602 8128
rect 7838 7982 7880 8128
rect 7560 7104 7880 7982
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 4928 7880 5952
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 4838 7880 4864
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 3840 7880 4602
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1458 7880 1600
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 7560 1040 7880 1222
rect 8560 9266 8880 11472
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 8560 1040 8880 2270
<< obsm4 >>
rect 13400 0 34000 13000
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 5102 9824 5338 9908
rect 5102 9760 5132 9824
rect 5132 9760 5148 9824
rect 5148 9760 5212 9824
rect 5212 9760 5228 9824
rect 5228 9760 5292 9824
rect 5292 9760 5308 9824
rect 5308 9760 5338 9824
rect 5102 9672 5338 9760
rect 5102 6496 5132 6528
rect 5132 6496 5148 6528
rect 5148 6496 5212 6528
rect 5212 6496 5228 6528
rect 5228 6496 5292 6528
rect 5292 6496 5308 6528
rect 5308 6496 5338 6528
rect 5102 6292 5338 6496
rect 5102 2912 5338 3148
rect 6102 10720 6338 10956
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 7602 8192 7838 8218
rect 7602 8128 7632 8192
rect 7632 8128 7648 8192
rect 7648 8128 7712 8192
rect 7712 8128 7728 8192
rect 7728 8128 7792 8192
rect 7792 8128 7808 8192
rect 7808 8128 7838 8192
rect 7602 7982 7838 8128
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 872 10956 9892 10998
rect 872 10720 6102 10956
rect 6338 10720 9892 10956
rect 872 10678 9892 10720
rect 872 9908 9892 9950
rect 872 9672 5102 9908
rect 5338 9672 9892 9908
rect 872 9630 9892 9672
rect 872 9266 9892 9308
rect 872 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 9892 9266
rect 872 8988 9892 9030
rect 872 8218 9892 8260
rect 872 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 9892 8218
rect 872 7940 9892 7982
rect 872 7576 9892 7618
rect 872 7340 6102 7576
rect 6338 7340 9892 7576
rect 872 7298 9892 7340
rect 872 6528 9892 6570
rect 872 6292 5102 6528
rect 5338 6292 9892 6528
rect 872 6250 9892 6292
rect 872 5886 9892 5928
rect 872 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 9892 5886
rect 872 5608 9892 5650
rect 872 4838 9892 4880
rect 872 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 9892 4838
rect 872 4560 9892 4602
rect 872 4196 9892 4238
rect 872 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 9892 4196
rect 872 3918 9892 3960
rect 872 3148 9892 3190
rect 872 2912 5102 3148
rect 5338 2912 9892 3148
rect 872 2870 9892 2912
rect 872 2506 9892 2548
rect 872 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 9892 2506
rect 872 2228 9892 2270
rect 872 1458 9892 1500
rect 872 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 9892 1458
rect 872 1180 9892 1222
<< obsm5 >>
rect 13400 0 34000 13000
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9568 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A_N
timestamp 1662439860
transform -1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__B
timestamp 1662439860
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A2
timestamp 1662439860
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A_N
timestamp 1662439860
transform -1 0 8924 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__C
timestamp 1662439860
transform -1 0 9568 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A0
timestamp 1662439860
transform -1 0 9384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A0
timestamp 1662439860
transform -1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1662439860
transform -1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__B
timestamp 1662439860
transform 1 0 6624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A_N
timestamp 1662439860
transform -1 0 6992 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__B
timestamp 1662439860
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1662439860
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__B
timestamp 1662439860
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A_N
timestamp 1662439860
transform 1 0 5244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__B
timestamp 1662439860
transform 1 0 4600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1662439860
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__B
timestamp 1662439860
transform -1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A_N
timestamp 1662439860
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__B
timestamp 1662439860
transform -1 0 2760 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1662439860
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__B
timestamp 1662439860
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A_N
timestamp 1662439860
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__B
timestamp 1662439860
transform -1 0 9568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1662439860
transform 1 0 3588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__B
timestamp 1662439860
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A_N
timestamp 1662439860
transform 1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__B
timestamp 1662439860
transform 1 0 2668 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1662439860
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__B
timestamp 1662439860
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A_N
timestamp 1662439860
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B
timestamp 1662439860
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1662439860
transform -1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__B
timestamp 1662439860
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A_N
timestamp 1662439860
transform -1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B
timestamp 1662439860
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1662439860
transform 1 0 8556 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B
timestamp 1662439860
transform -1 0 8096 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A_N
timestamp 1662439860
transform 1 0 8280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__B
timestamp 1662439860
transform -1 0 7452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1662439860
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B
timestamp 1662439860
transform -1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A_N
timestamp 1662439860
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__B
timestamp 1662439860
transform -1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1662439860
transform -1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B
timestamp 1662439860
transform -1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A_N
timestamp 1662439860
transform -1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B
timestamp 1662439860
transform 1 0 8004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1662439860
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B
timestamp 1662439860
transform -1 0 5520 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A_N
timestamp 1662439860
transform -1 0 5336 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B
timestamp 1662439860
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1662439860
transform 1 0 5428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B
timestamp 1662439860
transform -1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A_N
timestamp 1662439860
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B
timestamp 1662439860
transform -1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1662439860
transform 1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B
timestamp 1662439860
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A_N
timestamp 1662439860
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B
timestamp 1662439860
transform -1 0 6072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__D
timestamp 1662439860
transform -1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__RESET_B
timestamp 1662439860
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__RESET_B
timestamp 1662439860
transform -1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__RESET_B
timestamp 1662439860
transform -1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__RESET_B
timestamp 1662439860
transform 1 0 2852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__RESET_B
timestamp 1662439860
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__RESET_B
timestamp 1662439860
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__RESET_B
timestamp 1662439860
transform 1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__RESET_B
timestamp 1662439860
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__RESET_B
timestamp 1662439860
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__RESET_B
timestamp 1662439860
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__RESET_B
timestamp 1662439860
transform 1 0 8004 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__RESET_B
timestamp 1662439860
transform 1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__RESET_B
timestamp 1662439860
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__RESET_B
timestamp 1662439860
transform -1 0 7728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1662439860
transform -1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1662439860
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1662439860
transform -1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1662439860
transform -1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5704 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_64
timestamp 1662439860
transform 1 0 6808 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_80
timestamp 1662439860
transform 1 0 8280 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1662439860
transform 1 0 6072 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_68
timestamp 1662439860
transform 1 0 7176 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 7452 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 1662439860
transform 1 0 7820 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1662439860
transform 1 0 8096 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_82
timestamp 1662439860
transform 1 0 8464 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1662439860
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1662439860
transform 1 0 4968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_70
timestamp 1662439860
transform 1 0 7360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1662439860
transform 1 0 8556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_39
timestamp 1662439860
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1662439860
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_50
timestamp 1662439860
transform 1 0 5520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 1662439860
transform 1 0 6440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_76
timestamp 1662439860
transform 1 0 7912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp 1662439860
transform 1 0 9476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 1196 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1662439860
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 1196 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1662439860
transform 1 0 1196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1662439860
transform 1 0 3404 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_44
timestamp 1662439860
transform 1 0 4968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp 1662439860
transform 1 0 7912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1662439860
transform 1 0 1196 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1662439860
transform 1 0 2300 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_48
timestamp 1662439860
transform 1 0 5336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1662439860
transform 1 0 1196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1662439860
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1662439860
transform 1 0 1196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_35
timestamp 1662439860
transform 1 0 4140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1662439860
transform 1 0 1196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1662439860
transform 1 0 4416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1662439860
transform 1 0 8556 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1662439860
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1662439860
transform 1 0 1196 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_65
timestamp 1662439860
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1662439860
transform 1 0 1196 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1662439860
transform 1 0 1196 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1662439860
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_72
timestamp 1662439860
transform 1 0 7544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1662439860
transform 1 0 1196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 2300 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_24
timestamp 1662439860
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1662439860
transform 1 0 4968 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_48
timestamp 1662439860
transform 1 0 5336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_52
timestamp 1662439860
transform 1 0 5704 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_61
timestamp 1662439860
transform 1 0 6532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_66
timestamp 1662439860
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_71
timestamp 1662439860
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1662439860
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1662439860
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1662439860
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1662439860
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1662439860
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1662439860
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1662439860
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1662439860
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1662439860
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1662439860
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1662439860
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1662439860
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1662439860
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1662439860
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1662439860
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1662439860
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1662439860
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1662439860
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1662439860
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1662439860
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1662439860
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1662439860
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1662439860
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1662439860
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1662439860
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1662439860
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1662439860
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1662439860
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1662439860
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1662439860
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1662439860
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1662439860
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1662439860
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1662439860
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1662439860
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1662439860
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1662439860
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1662439860
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1662439860
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1662439860
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1662439860
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1662439860
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1662439860
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1662439860
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1662439860
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1662439860
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1662439860
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1662439860
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1662439860
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1662439860
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1662439860
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1662439860
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1662439860
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1662439860
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1662439860
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1662439860
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1662439860
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1662439860
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1662439860
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1662439860
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1662439860
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1662439860
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1662439860
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1662439860
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1662439860
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1662439860
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1662439860
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059__1
timestamp 1662439860
transform -1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060__14
timestamp 1662439860
transform -1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9384 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9384 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8648 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9476 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _066_
timestamp 1662439860
transform -1 0 9568 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6808 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _068_
timestamp 1662439860
transform 1 0 6164 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _069_
timestamp 1662439860
transform 1 0 3036 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _070_
timestamp 1662439860
transform -1 0 5244 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _071_
timestamp 1662439860
transform -1 0 8740 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _072_
timestamp 1662439860
transform 1 0 5428 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _073_
timestamp 1662439860
transform -1 0 9200 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _074_
timestamp 1662439860
transform -1 0 9384 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _075_
timestamp 1662439860
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _076_
timestamp 1662439860
transform -1 0 4232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _077_
timestamp 1662439860
transform 1 0 3680 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _078_
timestamp 1662439860
transform -1 0 4968 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _079_
timestamp 1662439860
transform 1 0 5336 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _080_
timestamp 1662439860
transform 1 0 3956 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _081_
timestamp 1662439860
transform 1 0 8096 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _082_
timestamp 1662439860
transform 1 0 7452 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _083_
timestamp 1662439860
transform 1 0 9016 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _084_
timestamp 1662439860
transform 1 0 7176 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _085_
timestamp 1662439860
transform -1 0 9200 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _086_
timestamp 1662439860
transform -1 0 8648 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _087_
timestamp 1662439860
transform 1 0 4140 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _088_
timestamp 1662439860
transform 1 0 3496 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _089_
timestamp 1662439860
transform 1 0 5152 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _090_
timestamp 1662439860
transform -1 0 6348 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _091_
timestamp 1662439860
transform -1 0 6808 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _092_
timestamp 1662439860
transform -1 0 6348 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _093__2
timestamp 1662439860
transform -1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094__3
timestamp 1662439860
transform -1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095__4
timestamp 1662439860
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096__5
timestamp 1662439860
transform -1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097__6
timestamp 1662439860
transform -1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098__7
timestamp 1662439860
transform -1 0 4600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099__8
timestamp 1662439860
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100__9
timestamp 1662439860
transform 1 0 6256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101__10
timestamp 1662439860
transform -1 0 7544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102__11
timestamp 1662439860
transform -1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103__12
timestamp 1662439860
transform -1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104__13
timestamp 1662439860
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5428 0 1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _106_
timestamp 1662439860
transform 1 0 2760 0 -1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _107_
timestamp 1662439860
transform 1 0 5060 0 1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _108_
timestamp 1662439860
transform 1 0 6072 0 1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _109_
timestamp 1662439860
transform 1 0 2760 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _110_
timestamp 1662439860
transform 1 0 2760 0 -1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _111_
timestamp 1662439860
transform 1 0 3312 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _112_
timestamp 1662439860
transform 1 0 6808 0 1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _113_
timestamp 1662439860
transform 1 0 6532 0 1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _114_
timestamp 1662439860
transform 1 0 6992 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _115_
timestamp 1662439860
transform 1 0 3312 0 -1 2176
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _116_
timestamp 1662439860
transform 1 0 3496 0 -1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _117_
timestamp 1662439860
transform 1 0 4600 0 -1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_2  _118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 6440 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _119_
timestamp 1662439860
transform 1 0 1564 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _120_
timestamp 1662439860
transform -1 0 3312 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _121_
timestamp 1662439860
transform 1 0 1472 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _122_
timestamp 1662439860
transform 1 0 1472 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _123_
timestamp 1662439860
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _124_
timestamp 1662439860
transform 1 0 3312 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _125_
timestamp 1662439860
transform 1 0 3312 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _126_
timestamp 1662439860
transform 1 0 4140 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _127_
timestamp 1662439860
transform 1 0 6164 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _128_
timestamp 1662439860
transform 1 0 6164 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _129_
timestamp 1662439860
transform 1 0 5980 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _130_
timestamp 1662439860
transform 1 0 6440 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _131_
timestamp 1662439860
transform 1 0 7636 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1662439860
transform 1 0 8832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1662439860
transform 1 0 8832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8740 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 6072 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1662439860
transform -1 0 8004 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 1662439860
transform -1 0 5152 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 1662439860
transform -1 0 5152 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 1662439860
transform 1 0 6164 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 1662439860
transform -1 0 6072 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9200 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6532 0 -1 4352
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1662439860
transform -1 0 8740 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1662439860
transform 1 0 2024 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1662439860
transform -1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1662439860
transform -1 0 4324 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1662439860
transform -1 0 6900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1662439860
transform -1 0 6072 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1662439860
transform -1 0 9016 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1662439860
transform -1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1662439860
transform -1 0 5980 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1662439860
transform -1 0 6440 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1662439860
transform 1 0 3496 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1662439860
transform -1 0 9016 0 -1 5440
box -38 -48 774 592
<< labels >>
flabel metal2 s 938 12200 994 13000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 5538 12200 5594 13000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 5998 12200 6054 13000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 6458 12200 6514 13000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 1398 12200 1454 13000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 4 nsew signal input
flabel metal2 s 1858 12200 1914 13000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 5 nsew signal input
flabel metal2 s 2318 12200 2374 13000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 6 nsew signal input
flabel metal2 s 2778 12200 2834 13000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 7 nsew signal input
flabel metal2 s 3238 12200 3294 13000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 8 nsew signal input
flabel metal2 s 3698 12200 3754 13000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 9 nsew signal input
flabel metal2 s 4158 12200 4214 13000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 10 nsew signal input
flabel metal2 s 4618 12200 4674 13000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 11 nsew signal input
flabel metal2 s 5078 12200 5134 13000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 12 nsew signal input
flabel metal3 s 14000 824 34000 944 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 13 nsew signal tristate
flabel metal3 s 14000 1640 34000 1760 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 14 nsew signal input
flabel metal3 s 14000 2048 34000 2168 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 15 nsew signal input
flabel metal3 s 14000 1232 34000 1352 0 FreeSans 480 0 0 0 one
port 16 nsew signal tristate
flabel metal3 s 14000 2456 34000 2576 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 17 nsew signal tristate
flabel metal3 s 14000 2864 34000 2984 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 18 nsew signal tristate
flabel metal3 s 14000 3272 34000 3392 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 19 nsew signal tristate
flabel metal3 s 14000 3680 34000 3800 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 20 nsew signal tristate
flabel metal3 s 14000 4088 34000 4208 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 21 nsew signal tristate
flabel metal3 s 14000 4496 34000 4616 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 22 nsew signal tristate
flabel metal3 s 14000 4904 34000 5024 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 23 nsew signal tristate
flabel metal3 s 14000 5312 34000 5432 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
flabel metal3 s 14000 5720 34000 5840 0 FreeSans 480 0 0 0 pad_gpio_in
port 25 nsew signal input
flabel metal3 s 14000 6128 34000 6248 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 26 nsew signal tristate
flabel metal3 s 14000 6536 34000 6656 0 FreeSans 480 0 0 0 pad_gpio_out
port 27 nsew signal tristate
flabel metal3 s 14000 6944 34000 7064 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 28 nsew signal tristate
flabel metal3 s 14000 7352 34000 7472 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 29 nsew signal tristate
flabel metal3 s 14000 7760 34000 7880 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 30 nsew signal tristate
flabel metal3 s 14000 8168 34000 8288 0 FreeSans 480 0 0 0 resetn
port 31 nsew signal input
flabel metal3 s 14000 8576 34000 8696 0 FreeSans 480 0 0 0 resetn_out
port 32 nsew signal tristate
flabel metal3 s 14000 8984 34000 9104 0 FreeSans 480 0 0 0 serial_clock
port 33 nsew signal input
flabel metal3 s 14000 9392 34000 9512 0 FreeSans 480 0 0 0 serial_clock_out
port 34 nsew signal tristate
flabel metal3 s 14000 9800 34000 9920 0 FreeSans 480 0 0 0 serial_data_in
port 35 nsew signal input
flabel metal3 s 14000 10208 34000 10328 0 FreeSans 480 0 0 0 serial_data_out
port 36 nsew signal tristate
flabel metal3 s 14000 10616 34000 10736 0 FreeSans 480 0 0 0 serial_load
port 37 nsew signal input
flabel metal3 s 14000 11024 34000 11144 0 FreeSans 480 0 0 0 serial_load_out
port 38 nsew signal tristate
flabel metal3 s 14000 11432 34000 11552 0 FreeSans 480 0 0 0 user_gpio_in
port 39 nsew signal tristate
flabel metal3 s 14000 11840 34000 11960 0 FreeSans 480 0 0 0 user_gpio_oeb
port 40 nsew signal input
flabel metal3 s 14000 12248 34000 12368 0 FreeSans 480 0 0 0 user_gpio_out
port 41 nsew signal input
flabel metal4 s 2560 1040 2880 11472 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 7560 1040 7880 11472 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 1180 9892 1500 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 4560 9892 4880 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 7940 9892 8260 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 3560 1040 3880 11472 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 8560 1040 8880 11472 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 2228 9892 2548 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 5608 9892 5928 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 8988 9892 9308 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 5060 1040 5380 11472 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 2870 9892 3190 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 6250 9892 6570 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 9630 9892 9950 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 6060 1040 6380 11472 0 FreeSans 1920 90 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 3918 9892 4238 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 7298 9892 7618 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 10678 9892 10998 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal3 s 14000 416 34000 536 0 FreeSans 480 0 0 0 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
