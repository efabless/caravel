magic
tech sky130A
timestamp 1638280046
<< obsli1 >>
rect 1434 2079 258450 73904
<< obsm1 >>
rect 191 684 261779 80712
<< metal2 >>
rect 193 81600 221 82200
rect 607 81600 635 82200
rect 1021 81600 1049 82200
rect 1435 81600 1463 82200
rect 1849 81600 1877 82200
rect 2263 81600 2291 82200
rect 2677 81600 2705 82200
rect 3137 81600 3165 82200
rect 3551 81600 3579 82200
rect 3965 81600 3993 82200
rect 4379 81600 4407 82200
rect 4793 81600 4821 82200
rect 5207 81600 5235 82200
rect 5621 81600 5649 82200
rect 6081 81600 6109 82200
rect 6495 81600 6523 82200
rect 6909 81600 6937 82200
rect 7323 81600 7351 82200
rect 7737 81600 7765 82200
rect 8151 81600 8179 82200
rect 8565 81600 8593 82200
rect 9025 81600 9053 82200
rect 9439 81600 9467 82200
rect 9853 81600 9881 82200
rect 10267 81600 10295 82200
rect 10681 81600 10709 82200
rect 11095 81600 11123 82200
rect 11509 81600 11537 82200
rect 11969 81600 11997 82200
rect 12383 81600 12411 82200
rect 12797 81600 12825 82200
rect 13211 81600 13239 82200
rect 13625 81600 13653 82200
rect 14039 81600 14067 82200
rect 14453 81600 14481 82200
rect 14913 81600 14941 82200
rect 15327 81600 15355 82200
rect 15741 81600 15769 82200
rect 16155 81600 16183 82200
rect 16569 81600 16597 82200
rect 16983 81600 17011 82200
rect 17397 81600 17425 82200
rect 17857 81600 17885 82200
rect 18271 81600 18299 82200
rect 18685 81600 18713 82200
rect 19099 81600 19127 82200
rect 19513 81600 19541 82200
rect 19927 81600 19955 82200
rect 20341 81600 20369 82200
rect 20801 81600 20829 82200
rect 21215 81600 21243 82200
rect 21629 81600 21657 82200
rect 22043 81600 22071 82200
rect 22457 81600 22485 82200
rect 22871 81600 22899 82200
rect 23285 81600 23313 82200
rect 23745 81600 23773 82200
rect 24159 81600 24187 82200
rect 24573 81600 24601 82200
rect 24987 81600 25015 82200
rect 25401 81600 25429 82200
rect 25815 81600 25843 82200
rect 26229 81600 26257 82200
rect 26689 81600 26717 82200
rect 27103 81600 27131 82200
rect 27517 81600 27545 82200
rect 27931 81600 27959 82200
rect 28345 81600 28373 82200
rect 28759 81600 28787 82200
rect 29173 81600 29201 82200
rect 29633 81600 29661 82200
rect 30047 81600 30075 82200
rect 30461 81600 30489 82200
rect 30875 81600 30903 82200
rect 31289 81600 31317 82200
rect 31703 81600 31731 82200
rect 32117 81600 32145 82200
rect 32577 81600 32605 82200
rect 32991 81600 33019 82200
rect 33405 81600 33433 82200
rect 33819 81600 33847 82200
rect 34233 81600 34261 82200
rect 34647 81600 34675 82200
rect 35061 81600 35089 82200
rect 35521 81600 35549 82200
rect 35935 81600 35963 82200
rect 36349 81600 36377 82200
rect 36763 81600 36791 82200
rect 37177 81600 37205 82200
rect 37591 81600 37619 82200
rect 38005 81600 38033 82200
rect 38465 81600 38493 82200
rect 38879 81600 38907 82200
rect 39293 81600 39321 82200
rect 39707 81600 39735 82200
rect 40121 81600 40149 82200
rect 40535 81600 40563 82200
rect 40949 81600 40977 82200
rect 41409 81600 41437 82200
rect 41823 81600 41851 82200
rect 42237 81600 42265 82200
rect 42651 81600 42679 82200
rect 43065 81600 43093 82200
rect 43479 81600 43507 82200
rect 43893 81600 43921 82200
rect 44353 81600 44381 82200
rect 44767 81600 44795 82200
rect 45181 81600 45209 82200
rect 45595 81600 45623 82200
rect 46009 81600 46037 82200
rect 46423 81600 46451 82200
rect 46837 81600 46865 82200
rect 47297 81600 47325 82200
rect 47711 81600 47739 82200
rect 48125 81600 48153 82200
rect 48539 81600 48567 82200
rect 48953 81600 48981 82200
rect 49367 81600 49395 82200
rect 49781 81600 49809 82200
rect 50241 81600 50269 82200
rect 50655 81600 50683 82200
rect 51069 81600 51097 82200
rect 51483 81600 51511 82200
rect 51897 81600 51925 82200
rect 52311 81600 52339 82200
rect 52725 81600 52753 82200
rect 53185 81600 53213 82200
rect 53599 81600 53627 82200
rect 54013 81600 54041 82200
rect 54427 81600 54455 82200
rect 54841 81600 54869 82200
rect 55255 81600 55283 82200
rect 55669 81600 55697 82200
rect 56129 81600 56157 82200
rect 56543 81600 56571 82200
rect 56957 81600 56985 82200
rect 57371 81600 57399 82200
rect 57785 81600 57813 82200
rect 58199 81600 58227 82200
rect 58613 81600 58641 82200
rect 59073 81600 59101 82200
rect 59487 81600 59515 82200
rect 59901 81600 59929 82200
rect 60315 81600 60343 82200
rect 60729 81600 60757 82200
rect 61143 81600 61171 82200
rect 61557 81600 61585 82200
rect 62017 81600 62045 82200
rect 62431 81600 62459 82200
rect 62845 81600 62873 82200
rect 63259 81600 63287 82200
rect 63673 81600 63701 82200
rect 64087 81600 64115 82200
rect 64501 81600 64529 82200
rect 64961 81600 64989 82200
rect 65375 81600 65403 82200
rect 65789 81600 65817 82200
rect 66203 81600 66231 82200
rect 66617 81600 66645 82200
rect 67031 81600 67059 82200
rect 67445 81600 67473 82200
rect 67905 81600 67933 82200
rect 68319 81600 68347 82200
rect 68733 81600 68761 82200
rect 69147 81600 69175 82200
rect 69561 81600 69589 82200
rect 69975 81600 70003 82200
rect 70389 81600 70417 82200
rect 70849 81600 70877 82200
rect 71263 81600 71291 82200
rect 71677 81600 71705 82200
rect 72091 81600 72119 82200
rect 72505 81600 72533 82200
rect 72919 81600 72947 82200
rect 73333 81600 73361 82200
rect 73793 81600 73821 82200
rect 74207 81600 74235 82200
rect 74621 81600 74649 82200
rect 75035 81600 75063 82200
rect 75449 81600 75477 82200
rect 75863 81600 75891 82200
rect 76277 81600 76305 82200
rect 76737 81600 76765 82200
rect 77151 81600 77179 82200
rect 77565 81600 77593 82200
rect 77979 81600 78007 82200
rect 78393 81600 78421 82200
rect 78807 81600 78835 82200
rect 79221 81600 79249 82200
rect 79681 81600 79709 82200
rect 80095 81600 80123 82200
rect 80509 81600 80537 82200
rect 80923 81600 80951 82200
rect 81337 81600 81365 82200
rect 81751 81600 81779 82200
rect 82165 81600 82193 82200
rect 82625 81600 82653 82200
rect 83039 81600 83067 82200
rect 83453 81600 83481 82200
rect 83867 81600 83895 82200
rect 84281 81600 84309 82200
rect 84695 81600 84723 82200
rect 85109 81600 85137 82200
rect 85569 81600 85597 82200
rect 85983 81600 86011 82200
rect 86397 81600 86425 82200
rect 86811 81600 86839 82200
rect 87225 81600 87253 82200
rect 87639 81600 87667 82200
rect 88053 81600 88081 82200
rect 88513 81600 88541 82200
rect 88927 81600 88955 82200
rect 89341 81600 89369 82200
rect 89755 81600 89783 82200
rect 90169 81600 90197 82200
rect 90583 81600 90611 82200
rect 90997 81600 91025 82200
rect 91457 81600 91485 82200
rect 91871 81600 91899 82200
rect 92285 81600 92313 82200
rect 92699 81600 92727 82200
rect 93113 81600 93141 82200
rect 93527 81600 93555 82200
rect 93941 81600 93969 82200
rect 94401 81600 94429 82200
rect 94815 81600 94843 82200
rect 95229 81600 95257 82200
rect 95643 81600 95671 82200
rect 96057 81600 96085 82200
rect 96471 81600 96499 82200
rect 96885 81600 96913 82200
rect 97345 81600 97373 82200
rect 97759 81600 97787 82200
rect 98173 81600 98201 82200
rect 98587 81600 98615 82200
rect 99001 81600 99029 82200
rect 99415 81600 99443 82200
rect 99829 81600 99857 82200
rect 100289 81600 100317 82200
rect 100703 81600 100731 82200
rect 101117 81600 101145 82200
rect 101531 81600 101559 82200
rect 101945 81600 101973 82200
rect 102359 81600 102387 82200
rect 102773 81600 102801 82200
rect 103233 81600 103261 82200
rect 103647 81600 103675 82200
rect 104061 81600 104089 82200
rect 104475 81600 104503 82200
rect 104889 81600 104917 82200
rect 105303 81600 105331 82200
rect 105717 81600 105745 82200
rect 106177 81600 106205 82200
rect 106591 81600 106619 82200
rect 107005 81600 107033 82200
rect 107419 81600 107447 82200
rect 107833 81600 107861 82200
rect 108247 81600 108275 82200
rect 108661 81600 108689 82200
rect 109121 81600 109149 82200
rect 109535 81600 109563 82200
rect 109949 81600 109977 82200
rect 110363 81600 110391 82200
rect 110777 81600 110805 82200
rect 111191 81600 111219 82200
rect 111605 81600 111633 82200
rect 112065 81600 112093 82200
rect 112479 81600 112507 82200
rect 112893 81600 112921 82200
rect 113307 81600 113335 82200
rect 113721 81600 113749 82200
rect 114135 81600 114163 82200
rect 114549 81600 114577 82200
rect 115009 81600 115037 82200
rect 115423 81600 115451 82200
rect 115837 81600 115865 82200
rect 116251 81600 116279 82200
rect 116665 81600 116693 82200
rect 117079 81600 117107 82200
rect 117493 81600 117521 82200
rect 117953 81600 117981 82200
rect 118367 81600 118395 82200
rect 118781 81600 118809 82200
rect 119195 81600 119223 82200
rect 119609 81600 119637 82200
rect 120023 81600 120051 82200
rect 120437 81600 120465 82200
rect 120897 81600 120925 82200
rect 121311 81600 121339 82200
rect 121725 81600 121753 82200
rect 122139 81600 122167 82200
rect 122553 81600 122581 82200
rect 122967 81600 122995 82200
rect 123381 81600 123409 82200
rect 123841 81600 123869 82200
rect 124255 81600 124283 82200
rect 124669 81600 124697 82200
rect 125083 81600 125111 82200
rect 125497 81600 125525 82200
rect 125911 81600 125939 82200
rect 126325 81600 126353 82200
rect 126785 81600 126813 82200
rect 127199 81600 127227 82200
rect 127613 81600 127641 82200
rect 128027 81600 128055 82200
rect 128441 81600 128469 82200
rect 128855 81600 128883 82200
rect 129269 81600 129297 82200
rect 129729 81600 129757 82200
rect 130143 81600 130171 82200
rect 130557 81600 130585 82200
rect 130971 81600 130999 82200
rect 131385 81600 131413 82200
rect 131799 81600 131827 82200
rect 132213 81600 132241 82200
rect 132673 81600 132701 82200
rect 133087 81600 133115 82200
rect 133501 81600 133529 82200
rect 133915 81600 133943 82200
rect 134329 81600 134357 82200
rect 134743 81600 134771 82200
rect 135157 81600 135185 82200
rect 135617 81600 135645 82200
rect 136031 81600 136059 82200
rect 136445 81600 136473 82200
rect 136859 81600 136887 82200
rect 137273 81600 137301 82200
rect 137687 81600 137715 82200
rect 138101 81600 138129 82200
rect 138561 81600 138589 82200
rect 138975 81600 139003 82200
rect 139389 81600 139417 82200
rect 139803 81600 139831 82200
rect 140217 81600 140245 82200
rect 140631 81600 140659 82200
rect 141045 81600 141073 82200
rect 141505 81600 141533 82200
rect 141919 81600 141947 82200
rect 142333 81600 142361 82200
rect 142747 81600 142775 82200
rect 143161 81600 143189 82200
rect 143575 81600 143603 82200
rect 143989 81600 144017 82200
rect 144449 81600 144477 82200
rect 144863 81600 144891 82200
rect 145277 81600 145305 82200
rect 145691 81600 145719 82200
rect 146105 81600 146133 82200
rect 146519 81600 146547 82200
rect 146933 81600 146961 82200
rect 147393 81600 147421 82200
rect 147807 81600 147835 82200
rect 148221 81600 148249 82200
rect 148635 81600 148663 82200
rect 149049 81600 149077 82200
rect 149463 81600 149491 82200
rect 149877 81600 149905 82200
rect 150337 81600 150365 82200
rect 150751 81600 150779 82200
rect 151165 81600 151193 82200
rect 151579 81600 151607 82200
rect 151993 81600 152021 82200
rect 152407 81600 152435 82200
rect 152821 81600 152849 82200
rect 153281 81600 153309 82200
rect 153695 81600 153723 82200
rect 154109 81600 154137 82200
rect 154523 81600 154551 82200
rect 154937 81600 154965 82200
rect 155351 81600 155379 82200
rect 155765 81600 155793 82200
rect 156225 81600 156253 82200
rect 156639 81600 156667 82200
rect 157053 81600 157081 82200
rect 157467 81600 157495 82200
rect 157881 81600 157909 82200
rect 158295 81600 158323 82200
rect 158709 81600 158737 82200
rect 159169 81600 159197 82200
rect 159583 81600 159611 82200
rect 159997 81600 160025 82200
rect 160411 81600 160439 82200
rect 160825 81600 160853 82200
rect 161239 81600 161267 82200
rect 161653 81600 161681 82200
rect 162113 81600 162141 82200
rect 162527 81600 162555 82200
rect 162941 81600 162969 82200
rect 163355 81600 163383 82200
rect 163769 81600 163797 82200
rect 164183 81600 164211 82200
rect 164597 81600 164625 82200
rect 165057 81600 165085 82200
rect 165471 81600 165499 82200
rect 165885 81600 165913 82200
rect 166299 81600 166327 82200
rect 166713 81600 166741 82200
rect 167127 81600 167155 82200
rect 167541 81600 167569 82200
rect 168001 81600 168029 82200
rect 168415 81600 168443 82200
rect 168829 81600 168857 82200
rect 169243 81600 169271 82200
rect 169657 81600 169685 82200
rect 170071 81600 170099 82200
rect 170485 81600 170513 82200
rect 170945 81600 170973 82200
rect 171359 81600 171387 82200
rect 171773 81600 171801 82200
rect 172187 81600 172215 82200
rect 172601 81600 172629 82200
rect 173015 81600 173043 82200
rect 173429 81600 173457 82200
rect 173889 81600 173917 82200
rect 174303 81600 174331 82200
rect 174717 81600 174745 82200
rect 175131 81600 175159 82200
rect 175545 81600 175573 82200
rect 175959 81600 175987 82200
rect 176373 81600 176401 82200
rect 176833 81600 176861 82200
rect 177247 81600 177275 82200
rect 177661 81600 177689 82200
rect 178075 81600 178103 82200
rect 178489 81600 178517 82200
rect 178903 81600 178931 82200
rect 179317 81600 179345 82200
rect 179777 81600 179805 82200
rect 180191 81600 180219 82200
rect 180605 81600 180633 82200
rect 181019 81600 181047 82200
rect 181433 81600 181461 82200
rect 181847 81600 181875 82200
rect 182261 81600 182289 82200
rect 182721 81600 182749 82200
rect 183135 81600 183163 82200
rect 183549 81600 183577 82200
rect 183963 81600 183991 82200
rect 184377 81600 184405 82200
rect 184791 81600 184819 82200
rect 185205 81600 185233 82200
rect 185665 81600 185693 82200
rect 186079 81600 186107 82200
rect 186493 81600 186521 82200
rect 186907 81600 186935 82200
rect 187321 81600 187349 82200
rect 187735 81600 187763 82200
rect 188149 81600 188177 82200
rect 188609 81600 188637 82200
rect 189023 81600 189051 82200
rect 189437 81600 189465 82200
rect 189851 81600 189879 82200
rect 190265 81600 190293 82200
rect 190679 81600 190707 82200
rect 191093 81600 191121 82200
rect 191553 81600 191581 82200
rect 191967 81600 191995 82200
rect 192381 81600 192409 82200
rect 192795 81600 192823 82200
rect 193209 81600 193237 82200
rect 193623 81600 193651 82200
rect 194037 81600 194065 82200
rect 194497 81600 194525 82200
rect 194911 81600 194939 82200
rect 195325 81600 195353 82200
rect 195739 81600 195767 82200
rect 196153 81600 196181 82200
rect 196567 81600 196595 82200
rect 196981 81600 197009 82200
rect 197441 81600 197469 82200
rect 197855 81600 197883 82200
rect 198269 81600 198297 82200
rect 198683 81600 198711 82200
rect 199097 81600 199125 82200
rect 199511 81600 199539 82200
rect 199925 81600 199953 82200
rect 200385 81600 200413 82200
rect 200799 81600 200827 82200
rect 201213 81600 201241 82200
rect 201627 81600 201655 82200
rect 202041 81600 202069 82200
rect 202455 81600 202483 82200
rect 202869 81600 202897 82200
rect 203329 81600 203357 82200
rect 203743 81600 203771 82200
rect 204157 81600 204185 82200
rect 204571 81600 204599 82200
rect 204985 81600 205013 82200
rect 205399 81600 205427 82200
rect 205813 81600 205841 82200
rect 206273 81600 206301 82200
rect 206687 81600 206715 82200
rect 207101 81600 207129 82200
rect 207515 81600 207543 82200
rect 207929 81600 207957 82200
rect 208343 81600 208371 82200
rect 208757 81600 208785 82200
rect 209217 81600 209245 82200
rect 209631 81600 209659 82200
rect 210045 81600 210073 82200
rect 210459 81600 210487 82200
rect 210873 81600 210901 82200
rect 211287 81600 211315 82200
rect 211701 81600 211729 82200
rect 212161 81600 212189 82200
rect 212575 81600 212603 82200
rect 212989 81600 213017 82200
rect 213403 81600 213431 82200
rect 213817 81600 213845 82200
rect 214231 81600 214259 82200
rect 214645 81600 214673 82200
rect 215105 81600 215133 82200
rect 215519 81600 215547 82200
rect 215933 81600 215961 82200
rect 216347 81600 216375 82200
rect 216761 81600 216789 82200
rect 217175 81600 217203 82200
rect 217589 81600 217617 82200
rect 218049 81600 218077 82200
rect 218463 81600 218491 82200
rect 218877 81600 218905 82200
rect 219291 81600 219319 82200
rect 219705 81600 219733 82200
rect 220119 81600 220147 82200
rect 220533 81600 220561 82200
rect 220993 81600 221021 82200
rect 221407 81600 221435 82200
rect 221821 81600 221849 82200
rect 222235 81600 222263 82200
rect 222649 81600 222677 82200
rect 223063 81600 223091 82200
rect 223477 81600 223505 82200
rect 223937 81600 223965 82200
rect 224351 81600 224379 82200
rect 224765 81600 224793 82200
rect 225179 81600 225207 82200
rect 225593 81600 225621 82200
rect 226007 81600 226035 82200
rect 226421 81600 226449 82200
rect 226881 81600 226909 82200
rect 227295 81600 227323 82200
rect 227709 81600 227737 82200
rect 228123 81600 228151 82200
rect 228537 81600 228565 82200
rect 228951 81600 228979 82200
rect 229365 81600 229393 82200
rect 229825 81600 229853 82200
rect 230239 81600 230267 82200
rect 230653 81600 230681 82200
rect 231067 81600 231095 82200
rect 231481 81600 231509 82200
rect 231895 81600 231923 82200
rect 232309 81600 232337 82200
rect 232769 81600 232797 82200
rect 233183 81600 233211 82200
rect 233597 81600 233625 82200
rect 234011 81600 234039 82200
rect 234425 81600 234453 82200
rect 234839 81600 234867 82200
rect 235253 81600 235281 82200
rect 235713 81600 235741 82200
rect 236127 81600 236155 82200
rect 236541 81600 236569 82200
rect 236955 81600 236983 82200
rect 237369 81600 237397 82200
rect 237783 81600 237811 82200
rect 238197 81600 238225 82200
rect 238657 81600 238685 82200
rect 239071 81600 239099 82200
rect 239485 81600 239513 82200
rect 239899 81600 239927 82200
rect 240313 81600 240341 82200
rect 240727 81600 240755 82200
rect 241141 81600 241169 82200
rect 241601 81600 241629 82200
rect 242015 81600 242043 82200
rect 242429 81600 242457 82200
rect 242843 81600 242871 82200
rect 243257 81600 243285 82200
rect 243671 81600 243699 82200
rect 244085 81600 244113 82200
rect 244545 81600 244573 82200
rect 244959 81600 244987 82200
rect 245373 81600 245401 82200
rect 245787 81600 245815 82200
rect 246201 81600 246229 82200
rect 246615 81600 246643 82200
rect 247029 81600 247057 82200
rect 247489 81600 247517 82200
rect 247903 81600 247931 82200
rect 248317 81600 248345 82200
rect 248731 81600 248759 82200
rect 249145 81600 249173 82200
rect 249559 81600 249587 82200
rect 249973 81600 250001 82200
rect 250433 81600 250461 82200
rect 250847 81600 250875 82200
rect 251261 81600 251289 82200
rect 251675 81600 251703 82200
rect 252089 81600 252117 82200
rect 252503 81600 252531 82200
rect 252917 81600 252945 82200
rect 253377 81600 253405 82200
rect 253791 81600 253819 82200
rect 254205 81600 254233 82200
rect 254619 81600 254647 82200
rect 255033 81600 255061 82200
rect 255447 81600 255475 82200
rect 255861 81600 255889 82200
rect 256321 81600 256349 82200
rect 256735 81600 256763 82200
rect 257149 81600 257177 82200
rect 257563 81600 257591 82200
rect 257977 81600 258005 82200
rect 258391 81600 258419 82200
rect 258805 81600 258833 82200
rect 259265 81600 259293 82200
rect 259679 81600 259707 82200
rect 260093 81600 260121 82200
rect 260507 81600 260535 82200
rect 260921 81600 260949 82200
rect 261335 81600 261363 82200
rect 261749 81600 261777 82200
rect 16385 -200 16413 400
rect 49137 -200 49165 400
rect 81889 -200 81917 400
rect 114641 -200 114669 400
rect 147393 -200 147421 400
rect 180145 -200 180173 400
rect 212897 -200 212925 400
rect 245649 -200 245677 400
<< obsm2 >>
rect 249 81572 579 81641
rect 663 81572 993 81641
rect 1077 81572 1407 81641
rect 1491 81572 1821 81641
rect 1905 81572 2235 81641
rect 2319 81572 2649 81641
rect 2733 81572 3109 81641
rect 3193 81572 3523 81641
rect 3607 81572 3937 81641
rect 4021 81572 4351 81641
rect 4435 81572 4765 81641
rect 4849 81572 5179 81641
rect 5263 81572 5593 81641
rect 5677 81572 6053 81641
rect 6137 81572 6467 81641
rect 6551 81572 6881 81641
rect 6965 81572 7295 81641
rect 7379 81572 7709 81641
rect 7793 81572 8123 81641
rect 8207 81572 8537 81641
rect 8621 81572 8997 81641
rect 9081 81572 9411 81641
rect 9495 81572 9825 81641
rect 9909 81572 10239 81641
rect 10323 81572 10653 81641
rect 10737 81572 11067 81641
rect 11151 81572 11481 81641
rect 11565 81572 11941 81641
rect 12025 81572 12355 81641
rect 12439 81572 12769 81641
rect 12853 81572 13183 81641
rect 13267 81572 13597 81641
rect 13681 81572 14011 81641
rect 14095 81572 14425 81641
rect 14509 81572 14885 81641
rect 14969 81572 15299 81641
rect 15383 81572 15713 81641
rect 15797 81572 16127 81641
rect 16211 81572 16541 81641
rect 16625 81572 16955 81641
rect 17039 81572 17369 81641
rect 17453 81572 17829 81641
rect 17913 81572 18243 81641
rect 18327 81572 18657 81641
rect 18741 81572 19071 81641
rect 19155 81572 19485 81641
rect 19569 81572 19899 81641
rect 19983 81572 20313 81641
rect 20397 81572 20773 81641
rect 20857 81572 21187 81641
rect 21271 81572 21601 81641
rect 21685 81572 22015 81641
rect 22099 81572 22429 81641
rect 22513 81572 22843 81641
rect 22927 81572 23257 81641
rect 23341 81572 23717 81641
rect 23801 81572 24131 81641
rect 24215 81572 24545 81641
rect 24629 81572 24959 81641
rect 25043 81572 25373 81641
rect 25457 81572 25787 81641
rect 25871 81572 26201 81641
rect 26285 81572 26661 81641
rect 26745 81572 27075 81641
rect 27159 81572 27489 81641
rect 27573 81572 27903 81641
rect 27987 81572 28317 81641
rect 28401 81572 28731 81641
rect 28815 81572 29145 81641
rect 29229 81572 29605 81641
rect 29689 81572 30019 81641
rect 30103 81572 30433 81641
rect 30517 81572 30847 81641
rect 30931 81572 31261 81641
rect 31345 81572 31675 81641
rect 31759 81572 32089 81641
rect 32173 81572 32549 81641
rect 32633 81572 32963 81641
rect 33047 81572 33377 81641
rect 33461 81572 33791 81641
rect 33875 81572 34205 81641
rect 34289 81572 34619 81641
rect 34703 81572 35033 81641
rect 35117 81572 35493 81641
rect 35577 81572 35907 81641
rect 35991 81572 36321 81641
rect 36405 81572 36735 81641
rect 36819 81572 37149 81641
rect 37233 81572 37563 81641
rect 37647 81572 37977 81641
rect 38061 81572 38437 81641
rect 38521 81572 38851 81641
rect 38935 81572 39265 81641
rect 39349 81572 39679 81641
rect 39763 81572 40093 81641
rect 40177 81572 40507 81641
rect 40591 81572 40921 81641
rect 41005 81572 41381 81641
rect 41465 81572 41795 81641
rect 41879 81572 42209 81641
rect 42293 81572 42623 81641
rect 42707 81572 43037 81641
rect 43121 81572 43451 81641
rect 43535 81572 43865 81641
rect 43949 81572 44325 81641
rect 44409 81572 44739 81641
rect 44823 81572 45153 81641
rect 45237 81572 45567 81641
rect 45651 81572 45981 81641
rect 46065 81572 46395 81641
rect 46479 81572 46809 81641
rect 46893 81572 47269 81641
rect 47353 81572 47683 81641
rect 47767 81572 48097 81641
rect 48181 81572 48511 81641
rect 48595 81572 48925 81641
rect 49009 81572 49339 81641
rect 49423 81572 49753 81641
rect 49837 81572 50213 81641
rect 50297 81572 50627 81641
rect 50711 81572 51041 81641
rect 51125 81572 51455 81641
rect 51539 81572 51869 81641
rect 51953 81572 52283 81641
rect 52367 81572 52697 81641
rect 52781 81572 53157 81641
rect 53241 81572 53571 81641
rect 53655 81572 53985 81641
rect 54069 81572 54399 81641
rect 54483 81572 54813 81641
rect 54897 81572 55227 81641
rect 55311 81572 55641 81641
rect 55725 81572 56101 81641
rect 56185 81572 56515 81641
rect 56599 81572 56929 81641
rect 57013 81572 57343 81641
rect 57427 81572 57757 81641
rect 57841 81572 58171 81641
rect 58255 81572 58585 81641
rect 58669 81572 59045 81641
rect 59129 81572 59459 81641
rect 59543 81572 59873 81641
rect 59957 81572 60287 81641
rect 60371 81572 60701 81641
rect 60785 81572 61115 81641
rect 61199 81572 61529 81641
rect 61613 81572 61989 81641
rect 62073 81572 62403 81641
rect 62487 81572 62817 81641
rect 62901 81572 63231 81641
rect 63315 81572 63645 81641
rect 63729 81572 64059 81641
rect 64143 81572 64473 81641
rect 64557 81572 64933 81641
rect 65017 81572 65347 81641
rect 65431 81572 65761 81641
rect 65845 81572 66175 81641
rect 66259 81572 66589 81641
rect 66673 81572 67003 81641
rect 67087 81572 67417 81641
rect 67501 81572 67877 81641
rect 67961 81572 68291 81641
rect 68375 81572 68705 81641
rect 68789 81572 69119 81641
rect 69203 81572 69533 81641
rect 69617 81572 69947 81641
rect 70031 81572 70361 81641
rect 70445 81572 70821 81641
rect 70905 81572 71235 81641
rect 71319 81572 71649 81641
rect 71733 81572 72063 81641
rect 72147 81572 72477 81641
rect 72561 81572 72891 81641
rect 72975 81572 73305 81641
rect 73389 81572 73765 81641
rect 73849 81572 74179 81641
rect 74263 81572 74593 81641
rect 74677 81572 75007 81641
rect 75091 81572 75421 81641
rect 75505 81572 75835 81641
rect 75919 81572 76249 81641
rect 76333 81572 76709 81641
rect 76793 81572 77123 81641
rect 77207 81572 77537 81641
rect 77621 81572 77951 81641
rect 78035 81572 78365 81641
rect 78449 81572 78779 81641
rect 78863 81572 79193 81641
rect 79277 81572 79653 81641
rect 79737 81572 80067 81641
rect 80151 81572 80481 81641
rect 80565 81572 80895 81641
rect 80979 81572 81309 81641
rect 81393 81572 81723 81641
rect 81807 81572 82137 81641
rect 82221 81572 82597 81641
rect 82681 81572 83011 81641
rect 83095 81572 83425 81641
rect 83509 81572 83839 81641
rect 83923 81572 84253 81641
rect 84337 81572 84667 81641
rect 84751 81572 85081 81641
rect 85165 81572 85541 81641
rect 85625 81572 85955 81641
rect 86039 81572 86369 81641
rect 86453 81572 86783 81641
rect 86867 81572 87197 81641
rect 87281 81572 87611 81641
rect 87695 81572 88025 81641
rect 88109 81572 88485 81641
rect 88569 81572 88899 81641
rect 88983 81572 89313 81641
rect 89397 81572 89727 81641
rect 89811 81572 90141 81641
rect 90225 81572 90555 81641
rect 90639 81572 90969 81641
rect 91053 81572 91429 81641
rect 91513 81572 91843 81641
rect 91927 81572 92257 81641
rect 92341 81572 92671 81641
rect 92755 81572 93085 81641
rect 93169 81572 93499 81641
rect 93583 81572 93913 81641
rect 93997 81572 94373 81641
rect 94457 81572 94787 81641
rect 94871 81572 95201 81641
rect 95285 81572 95615 81641
rect 95699 81572 96029 81641
rect 96113 81572 96443 81641
rect 96527 81572 96857 81641
rect 96941 81572 97317 81641
rect 97401 81572 97731 81641
rect 97815 81572 98145 81641
rect 98229 81572 98559 81641
rect 98643 81572 98973 81641
rect 99057 81572 99387 81641
rect 99471 81572 99801 81641
rect 99885 81572 100261 81641
rect 100345 81572 100675 81641
rect 100759 81572 101089 81641
rect 101173 81572 101503 81641
rect 101587 81572 101917 81641
rect 102001 81572 102331 81641
rect 102415 81572 102745 81641
rect 102829 81572 103205 81641
rect 103289 81572 103619 81641
rect 103703 81572 104033 81641
rect 104117 81572 104447 81641
rect 104531 81572 104861 81641
rect 104945 81572 105275 81641
rect 105359 81572 105689 81641
rect 105773 81572 106149 81641
rect 106233 81572 106563 81641
rect 106647 81572 106977 81641
rect 107061 81572 107391 81641
rect 107475 81572 107805 81641
rect 107889 81572 108219 81641
rect 108303 81572 108633 81641
rect 108717 81572 109093 81641
rect 109177 81572 109507 81641
rect 109591 81572 109921 81641
rect 110005 81572 110335 81641
rect 110419 81572 110749 81641
rect 110833 81572 111163 81641
rect 111247 81572 111577 81641
rect 111661 81572 112037 81641
rect 112121 81572 112451 81641
rect 112535 81572 112865 81641
rect 112949 81572 113279 81641
rect 113363 81572 113693 81641
rect 113777 81572 114107 81641
rect 114191 81572 114521 81641
rect 114605 81572 114981 81641
rect 115065 81572 115395 81641
rect 115479 81572 115809 81641
rect 115893 81572 116223 81641
rect 116307 81572 116637 81641
rect 116721 81572 117051 81641
rect 117135 81572 117465 81641
rect 117549 81572 117925 81641
rect 118009 81572 118339 81641
rect 118423 81572 118753 81641
rect 118837 81572 119167 81641
rect 119251 81572 119581 81641
rect 119665 81572 119995 81641
rect 120079 81572 120409 81641
rect 120493 81572 120869 81641
rect 120953 81572 121283 81641
rect 121367 81572 121697 81641
rect 121781 81572 122111 81641
rect 122195 81572 122525 81641
rect 122609 81572 122939 81641
rect 123023 81572 123353 81641
rect 123437 81572 123813 81641
rect 123897 81572 124227 81641
rect 124311 81572 124641 81641
rect 124725 81572 125055 81641
rect 125139 81572 125469 81641
rect 125553 81572 125883 81641
rect 125967 81572 126297 81641
rect 126381 81572 126757 81641
rect 126841 81572 127171 81641
rect 127255 81572 127585 81641
rect 127669 81572 127999 81641
rect 128083 81572 128413 81641
rect 128497 81572 128827 81641
rect 128911 81572 129241 81641
rect 129325 81572 129701 81641
rect 129785 81572 130115 81641
rect 130199 81572 130529 81641
rect 130613 81572 130943 81641
rect 131027 81572 131357 81641
rect 131441 81572 131771 81641
rect 131855 81572 132185 81641
rect 132269 81572 132645 81641
rect 132729 81572 133059 81641
rect 133143 81572 133473 81641
rect 133557 81572 133887 81641
rect 133971 81572 134301 81641
rect 134385 81572 134715 81641
rect 134799 81572 135129 81641
rect 135213 81572 135589 81641
rect 135673 81572 136003 81641
rect 136087 81572 136417 81641
rect 136501 81572 136831 81641
rect 136915 81572 137245 81641
rect 137329 81572 137659 81641
rect 137743 81572 138073 81641
rect 138157 81572 138533 81641
rect 138617 81572 138947 81641
rect 139031 81572 139361 81641
rect 139445 81572 139775 81641
rect 139859 81572 140189 81641
rect 140273 81572 140603 81641
rect 140687 81572 141017 81641
rect 141101 81572 141477 81641
rect 141561 81572 141891 81641
rect 141975 81572 142305 81641
rect 142389 81572 142719 81641
rect 142803 81572 143133 81641
rect 143217 81572 143547 81641
rect 143631 81572 143961 81641
rect 144045 81572 144421 81641
rect 144505 81572 144835 81641
rect 144919 81572 145249 81641
rect 145333 81572 145663 81641
rect 145747 81572 146077 81641
rect 146161 81572 146491 81641
rect 146575 81572 146905 81641
rect 146989 81572 147365 81641
rect 147449 81572 147779 81641
rect 147863 81572 148193 81641
rect 148277 81572 148607 81641
rect 148691 81572 149021 81641
rect 149105 81572 149435 81641
rect 149519 81572 149849 81641
rect 149933 81572 150309 81641
rect 150393 81572 150723 81641
rect 150807 81572 151137 81641
rect 151221 81572 151551 81641
rect 151635 81572 151965 81641
rect 152049 81572 152379 81641
rect 152463 81572 152793 81641
rect 152877 81572 153253 81641
rect 153337 81572 153667 81641
rect 153751 81572 154081 81641
rect 154165 81572 154495 81641
rect 154579 81572 154909 81641
rect 154993 81572 155323 81641
rect 155407 81572 155737 81641
rect 155821 81572 156197 81641
rect 156281 81572 156611 81641
rect 156695 81572 157025 81641
rect 157109 81572 157439 81641
rect 157523 81572 157853 81641
rect 157937 81572 158267 81641
rect 158351 81572 158681 81641
rect 158765 81572 159141 81641
rect 159225 81572 159555 81641
rect 159639 81572 159969 81641
rect 160053 81572 160383 81641
rect 160467 81572 160797 81641
rect 160881 81572 161211 81641
rect 161295 81572 161625 81641
rect 161709 81572 162085 81641
rect 162169 81572 162499 81641
rect 162583 81572 162913 81641
rect 162997 81572 163327 81641
rect 163411 81572 163741 81641
rect 163825 81572 164155 81641
rect 164239 81572 164569 81641
rect 164653 81572 165029 81641
rect 165113 81572 165443 81641
rect 165527 81572 165857 81641
rect 165941 81572 166271 81641
rect 166355 81572 166685 81641
rect 166769 81572 167099 81641
rect 167183 81572 167513 81641
rect 167597 81572 167973 81641
rect 168057 81572 168387 81641
rect 168471 81572 168801 81641
rect 168885 81572 169215 81641
rect 169299 81572 169629 81641
rect 169713 81572 170043 81641
rect 170127 81572 170457 81641
rect 170541 81572 170917 81641
rect 171001 81572 171331 81641
rect 171415 81572 171745 81641
rect 171829 81572 172159 81641
rect 172243 81572 172573 81641
rect 172657 81572 172987 81641
rect 173071 81572 173401 81641
rect 173485 81572 173861 81641
rect 173945 81572 174275 81641
rect 174359 81572 174689 81641
rect 174773 81572 175103 81641
rect 175187 81572 175517 81641
rect 175601 81572 175931 81641
rect 176015 81572 176345 81641
rect 176429 81572 176805 81641
rect 176889 81572 177219 81641
rect 177303 81572 177633 81641
rect 177717 81572 178047 81641
rect 178131 81572 178461 81641
rect 178545 81572 178875 81641
rect 178959 81572 179289 81641
rect 179373 81572 179749 81641
rect 179833 81572 180163 81641
rect 180247 81572 180577 81641
rect 180661 81572 180991 81641
rect 181075 81572 181405 81641
rect 181489 81572 181819 81641
rect 181903 81572 182233 81641
rect 182317 81572 182693 81641
rect 182777 81572 183107 81641
rect 183191 81572 183521 81641
rect 183605 81572 183935 81641
rect 184019 81572 184349 81641
rect 184433 81572 184763 81641
rect 184847 81572 185177 81641
rect 185261 81572 185637 81641
rect 185721 81572 186051 81641
rect 186135 81572 186465 81641
rect 186549 81572 186879 81641
rect 186963 81572 187293 81641
rect 187377 81572 187707 81641
rect 187791 81572 188121 81641
rect 188205 81572 188581 81641
rect 188665 81572 188995 81641
rect 189079 81572 189409 81641
rect 189493 81572 189823 81641
rect 189907 81572 190237 81641
rect 190321 81572 190651 81641
rect 190735 81572 191065 81641
rect 191149 81572 191525 81641
rect 191609 81572 191939 81641
rect 192023 81572 192353 81641
rect 192437 81572 192767 81641
rect 192851 81572 193181 81641
rect 193265 81572 193595 81641
rect 193679 81572 194009 81641
rect 194093 81572 194469 81641
rect 194553 81572 194883 81641
rect 194967 81572 195297 81641
rect 195381 81572 195711 81641
rect 195795 81572 196125 81641
rect 196209 81572 196539 81641
rect 196623 81572 196953 81641
rect 197037 81572 197413 81641
rect 197497 81572 197827 81641
rect 197911 81572 198241 81641
rect 198325 81572 198655 81641
rect 198739 81572 199069 81641
rect 199153 81572 199483 81641
rect 199567 81572 199897 81641
rect 199981 81572 200357 81641
rect 200441 81572 200771 81641
rect 200855 81572 201185 81641
rect 201269 81572 201599 81641
rect 201683 81572 202013 81641
rect 202097 81572 202427 81641
rect 202511 81572 202841 81641
rect 202925 81572 203301 81641
rect 203385 81572 203715 81641
rect 203799 81572 204129 81641
rect 204213 81572 204543 81641
rect 204627 81572 204957 81641
rect 205041 81572 205371 81641
rect 205455 81572 205785 81641
rect 205869 81572 206245 81641
rect 206329 81572 206659 81641
rect 206743 81572 207073 81641
rect 207157 81572 207487 81641
rect 207571 81572 207901 81641
rect 207985 81572 208315 81641
rect 208399 81572 208729 81641
rect 208813 81572 209189 81641
rect 209273 81572 209603 81641
rect 209687 81572 210017 81641
rect 210101 81572 210431 81641
rect 210515 81572 210845 81641
rect 210929 81572 211259 81641
rect 211343 81572 211673 81641
rect 211757 81572 212133 81641
rect 212217 81572 212547 81641
rect 212631 81572 212961 81641
rect 213045 81572 213375 81641
rect 213459 81572 213789 81641
rect 213873 81572 214203 81641
rect 214287 81572 214617 81641
rect 214701 81572 215077 81641
rect 215161 81572 215491 81641
rect 215575 81572 215905 81641
rect 215989 81572 216319 81641
rect 216403 81572 216733 81641
rect 216817 81572 217147 81641
rect 217231 81572 217561 81641
rect 217645 81572 218021 81641
rect 218105 81572 218435 81641
rect 218519 81572 218849 81641
rect 218933 81572 219263 81641
rect 219347 81572 219677 81641
rect 219761 81572 220091 81641
rect 220175 81572 220505 81641
rect 220589 81572 220965 81641
rect 221049 81572 221379 81641
rect 221463 81572 221793 81641
rect 221877 81572 222207 81641
rect 222291 81572 222621 81641
rect 222705 81572 223035 81641
rect 223119 81572 223449 81641
rect 223533 81572 223909 81641
rect 223993 81572 224323 81641
rect 224407 81572 224737 81641
rect 224821 81572 225151 81641
rect 225235 81572 225565 81641
rect 225649 81572 225979 81641
rect 226063 81572 226393 81641
rect 226477 81572 226853 81641
rect 226937 81572 227267 81641
rect 227351 81572 227681 81641
rect 227765 81572 228095 81641
rect 228179 81572 228509 81641
rect 228593 81572 228923 81641
rect 229007 81572 229337 81641
rect 229421 81572 229797 81641
rect 229881 81572 230211 81641
rect 230295 81572 230625 81641
rect 230709 81572 231039 81641
rect 231123 81572 231453 81641
rect 231537 81572 231867 81641
rect 231951 81572 232281 81641
rect 232365 81572 232741 81641
rect 232825 81572 233155 81641
rect 233239 81572 233569 81641
rect 233653 81572 233983 81641
rect 234067 81572 234397 81641
rect 234481 81572 234811 81641
rect 234895 81572 235225 81641
rect 235309 81572 235685 81641
rect 235769 81572 236099 81641
rect 236183 81572 236513 81641
rect 236597 81572 236927 81641
rect 237011 81572 237341 81641
rect 237425 81572 237755 81641
rect 237839 81572 238169 81641
rect 238253 81572 238629 81641
rect 238713 81572 239043 81641
rect 239127 81572 239457 81641
rect 239541 81572 239871 81641
rect 239955 81572 240285 81641
rect 240369 81572 240699 81641
rect 240783 81572 241113 81641
rect 241197 81572 241573 81641
rect 241657 81572 241987 81641
rect 242071 81572 242401 81641
rect 242485 81572 242815 81641
rect 242899 81572 243229 81641
rect 243313 81572 243643 81641
rect 243727 81572 244057 81641
rect 244141 81572 244517 81641
rect 244601 81572 244931 81641
rect 245015 81572 245345 81641
rect 245429 81572 245759 81641
rect 245843 81572 246173 81641
rect 246257 81572 246587 81641
rect 246671 81572 247001 81641
rect 247085 81572 247461 81641
rect 247545 81572 247875 81641
rect 247959 81572 248289 81641
rect 248373 81572 248703 81641
rect 248787 81572 249117 81641
rect 249201 81572 249531 81641
rect 249615 81572 249945 81641
rect 250029 81572 250405 81641
rect 250489 81572 250819 81641
rect 250903 81572 251233 81641
rect 251317 81572 251647 81641
rect 251731 81572 252061 81641
rect 252145 81572 252475 81641
rect 252559 81572 252889 81641
rect 252973 81572 253349 81641
rect 253433 81572 253763 81641
rect 253847 81572 254177 81641
rect 254261 81572 254591 81641
rect 254675 81572 255005 81641
rect 255089 81572 255419 81641
rect 255503 81572 255833 81641
rect 255917 81572 256293 81641
rect 256377 81572 256707 81641
rect 256791 81572 257121 81641
rect 257205 81572 257535 81641
rect 257619 81572 257949 81641
rect 258033 81572 258363 81641
rect 258447 81572 258777 81641
rect 258861 81572 259237 81641
rect 259321 81572 259651 81641
rect 259735 81572 260065 81641
rect 260149 81572 260479 81641
rect 260563 81572 260893 81641
rect 260977 81572 261307 81641
rect 261391 81572 261721 81641
rect 194 428 261776 81572
rect 194 355 16357 428
rect 16441 355 49109 428
rect 49193 355 81861 428
rect 81945 355 114613 428
rect 114697 355 147365 428
rect 147449 355 180117 428
rect 180201 355 212869 428
rect 212953 355 245621 428
rect 245705 355 261776 428
<< metal3 >>
rect 261600 81536 262200 81596
rect 261600 80788 262200 80848
rect 261600 80040 262200 80100
rect 261600 79292 262200 79352
rect 261600 78544 262200 78604
rect 261600 77796 262200 77856
rect 261600 77048 262200 77108
rect 261600 76300 262200 76360
rect 261600 75552 262200 75612
rect 261600 74804 262200 74864
rect 261600 74056 262200 74116
rect 261600 73308 262200 73368
rect 261600 72560 262200 72620
rect 261600 71812 262200 71872
rect 261600 71064 262200 71124
rect 261600 70248 262200 70308
rect 261600 69500 262200 69560
rect 261600 68752 262200 68812
rect 261600 68004 262200 68064
rect 261600 67256 262200 67316
rect 261600 66508 262200 66568
rect 261600 65760 262200 65820
rect 261600 65012 262200 65072
rect 261600 64264 262200 64324
rect 261600 63516 262200 63576
rect 261600 62768 262200 62828
rect 261600 62020 262200 62080
rect 261600 61272 262200 61332
rect 261600 60524 262200 60584
rect 261600 59776 262200 59836
rect 261600 59028 262200 59088
rect 261600 58212 262200 58272
rect 261600 57464 262200 57524
rect 261600 56716 262200 56776
rect 261600 55968 262200 56028
rect 261600 55220 262200 55280
rect 261600 54472 262200 54532
rect 261600 53724 262200 53784
rect 261600 52976 262200 53036
rect 261600 52228 262200 52288
rect 261600 51480 262200 51540
rect 261600 50732 262200 50792
rect 261600 49984 262200 50044
rect 261600 49236 262200 49296
rect 261600 48488 262200 48548
rect 261600 47740 262200 47800
rect 261600 46924 262200 46984
rect 261600 46176 262200 46236
rect 261600 45428 262200 45488
rect 261600 44680 262200 44740
rect 261600 43932 262200 43992
rect 261600 43184 262200 43244
rect 261600 42436 262200 42496
rect 261600 41688 262200 41748
rect 261600 40940 262200 41000
rect 261600 40192 262200 40252
rect 261600 39444 262200 39504
rect 261600 38696 262200 38756
rect 261600 37948 262200 38008
rect 261600 37200 262200 37260
rect 261600 36452 262200 36512
rect 261600 35704 262200 35764
rect 261600 34888 262200 34948
rect 261600 34140 262200 34200
rect 261600 33392 262200 33452
rect 261600 32644 262200 32704
rect 261600 31896 262200 31956
rect 261600 31148 262200 31208
rect 261600 30400 262200 30460
rect 261600 29652 262200 29712
rect 261600 28904 262200 28964
rect 261600 28156 262200 28216
rect 261600 27408 262200 27468
rect 261600 26660 262200 26720
rect 261600 25912 262200 25972
rect 261600 25164 262200 25224
rect 261600 24416 262200 24476
rect 261600 23600 262200 23660
rect 261600 22852 262200 22912
rect 261600 22104 262200 22164
rect 261600 21356 262200 21416
rect 261600 20608 262200 20668
rect 261600 19860 262200 19920
rect 261600 19112 262200 19172
rect 261600 18364 262200 18424
rect 261600 17616 262200 17676
rect 261600 16868 262200 16928
rect 261600 16120 262200 16180
rect 261600 15372 262200 15432
rect 261600 14624 262200 14684
rect 261600 13876 262200 13936
rect 261600 13128 262200 13188
rect 261600 12380 262200 12440
rect 261600 11564 262200 11624
rect 261600 10816 262200 10876
rect 261600 10068 262200 10128
rect 261600 9320 262200 9380
rect 261600 8572 262200 8632
rect 261600 7824 262200 7884
rect 261600 7076 262200 7136
rect 261600 6328 262200 6388
rect 261600 5580 262200 5640
rect 261600 4832 262200 4892
rect 261600 4084 262200 4144
rect 261600 3336 262200 3396
rect 261600 2588 262200 2648
rect 261600 1840 262200 1900
rect 261600 1092 262200 1152
rect 261600 344 262200 404
<< obsm3 >>
rect 1334 81496 261560 81582
rect 1334 80888 261600 81496
rect 1334 80748 261560 80888
rect 1334 80140 261600 80748
rect 1334 80000 261560 80140
rect 1334 79392 261600 80000
rect 1334 79252 261560 79392
rect 1334 78644 261600 79252
rect 1334 78504 261560 78644
rect 1334 77896 261600 78504
rect 1334 77756 261560 77896
rect 1334 77148 261600 77756
rect 1334 77008 261560 77148
rect 1334 76400 261600 77008
rect 1334 76260 261560 76400
rect 1334 75652 261600 76260
rect 1334 75512 261560 75652
rect 1334 74904 261600 75512
rect 1334 74764 261560 74904
rect 1334 74156 261600 74764
rect 1334 74016 261560 74156
rect 1334 73408 261600 74016
rect 1334 73268 261560 73408
rect 1334 72660 261600 73268
rect 1334 72520 261560 72660
rect 1334 71912 261600 72520
rect 1334 71772 261560 71912
rect 1334 71164 261600 71772
rect 1334 71024 261560 71164
rect 1334 70348 261600 71024
rect 1334 70208 261560 70348
rect 1334 69600 261600 70208
rect 1334 69460 261560 69600
rect 1334 68852 261600 69460
rect 1334 68712 261560 68852
rect 1334 68104 261600 68712
rect 1334 67964 261560 68104
rect 1334 67356 261600 67964
rect 1334 67216 261560 67356
rect 1334 66608 261600 67216
rect 1334 66468 261560 66608
rect 1334 65860 261600 66468
rect 1334 65720 261560 65860
rect 1334 65112 261600 65720
rect 1334 64972 261560 65112
rect 1334 64364 261600 64972
rect 1334 64224 261560 64364
rect 1334 63616 261600 64224
rect 1334 63476 261560 63616
rect 1334 62868 261600 63476
rect 1334 62728 261560 62868
rect 1334 62120 261600 62728
rect 1334 61980 261560 62120
rect 1334 61372 261600 61980
rect 1334 61232 261560 61372
rect 1334 60624 261600 61232
rect 1334 60484 261560 60624
rect 1334 59876 261600 60484
rect 1334 59736 261560 59876
rect 1334 59128 261600 59736
rect 1334 58988 261560 59128
rect 1334 58312 261600 58988
rect 1334 58172 261560 58312
rect 1334 57564 261600 58172
rect 1334 57424 261560 57564
rect 1334 56816 261600 57424
rect 1334 56676 261560 56816
rect 1334 56068 261600 56676
rect 1334 55928 261560 56068
rect 1334 55320 261600 55928
rect 1334 55180 261560 55320
rect 1334 54572 261600 55180
rect 1334 54432 261560 54572
rect 1334 53824 261600 54432
rect 1334 53684 261560 53824
rect 1334 53076 261600 53684
rect 1334 52936 261560 53076
rect 1334 52328 261600 52936
rect 1334 52188 261560 52328
rect 1334 51580 261600 52188
rect 1334 51440 261560 51580
rect 1334 50832 261600 51440
rect 1334 50692 261560 50832
rect 1334 50084 261600 50692
rect 1334 49944 261560 50084
rect 1334 49336 261600 49944
rect 1334 49196 261560 49336
rect 1334 48588 261600 49196
rect 1334 48448 261560 48588
rect 1334 47840 261600 48448
rect 1334 47700 261560 47840
rect 1334 47024 261600 47700
rect 1334 46884 261560 47024
rect 1334 46276 261600 46884
rect 1334 46136 261560 46276
rect 1334 45528 261600 46136
rect 1334 45388 261560 45528
rect 1334 44780 261600 45388
rect 1334 44640 261560 44780
rect 1334 44032 261600 44640
rect 1334 43892 261560 44032
rect 1334 43284 261600 43892
rect 1334 43144 261560 43284
rect 1334 42536 261600 43144
rect 1334 42396 261560 42536
rect 1334 41788 261600 42396
rect 1334 41648 261560 41788
rect 1334 41040 261600 41648
rect 1334 40900 261560 41040
rect 1334 40292 261600 40900
rect 1334 40152 261560 40292
rect 1334 39544 261600 40152
rect 1334 39404 261560 39544
rect 1334 38796 261600 39404
rect 1334 38656 261560 38796
rect 1334 38048 261600 38656
rect 1334 37908 261560 38048
rect 1334 37300 261600 37908
rect 1334 37160 261560 37300
rect 1334 36552 261600 37160
rect 1334 36412 261560 36552
rect 1334 35804 261600 36412
rect 1334 35664 261560 35804
rect 1334 34988 261600 35664
rect 1334 34848 261560 34988
rect 1334 34240 261600 34848
rect 1334 34100 261560 34240
rect 1334 33492 261600 34100
rect 1334 33352 261560 33492
rect 1334 32744 261600 33352
rect 1334 32604 261560 32744
rect 1334 31996 261600 32604
rect 1334 31856 261560 31996
rect 1334 31248 261600 31856
rect 1334 31108 261560 31248
rect 1334 30500 261600 31108
rect 1334 30360 261560 30500
rect 1334 29752 261600 30360
rect 1334 29612 261560 29752
rect 1334 29004 261600 29612
rect 1334 28864 261560 29004
rect 1334 28256 261600 28864
rect 1334 28116 261560 28256
rect 1334 27508 261600 28116
rect 1334 27368 261560 27508
rect 1334 26760 261600 27368
rect 1334 26620 261560 26760
rect 1334 26012 261600 26620
rect 1334 25872 261560 26012
rect 1334 25264 261600 25872
rect 1334 25124 261560 25264
rect 1334 24516 261600 25124
rect 1334 24376 261560 24516
rect 1334 23700 261600 24376
rect 1334 23560 261560 23700
rect 1334 22952 261600 23560
rect 1334 22812 261560 22952
rect 1334 22204 261600 22812
rect 1334 22064 261560 22204
rect 1334 21456 261600 22064
rect 1334 21316 261560 21456
rect 1334 20708 261600 21316
rect 1334 20568 261560 20708
rect 1334 19960 261600 20568
rect 1334 19820 261560 19960
rect 1334 19212 261600 19820
rect 1334 19072 261560 19212
rect 1334 18464 261600 19072
rect 1334 18324 261560 18464
rect 1334 17716 261600 18324
rect 1334 17576 261560 17716
rect 1334 16968 261600 17576
rect 1334 16828 261560 16968
rect 1334 16220 261600 16828
rect 1334 16080 261560 16220
rect 1334 15472 261600 16080
rect 1334 15332 261560 15472
rect 1334 14724 261600 15332
rect 1334 14584 261560 14724
rect 1334 13976 261600 14584
rect 1334 13836 261560 13976
rect 1334 13228 261600 13836
rect 1334 13088 261560 13228
rect 1334 12480 261600 13088
rect 1334 12340 261560 12480
rect 1334 11664 261600 12340
rect 1334 11524 261560 11664
rect 1334 10916 261600 11524
rect 1334 10776 261560 10916
rect 1334 10168 261600 10776
rect 1334 10028 261560 10168
rect 1334 9420 261600 10028
rect 1334 9280 261560 9420
rect 1334 8672 261600 9280
rect 1334 8532 261560 8672
rect 1334 7924 261600 8532
rect 1334 7784 261560 7924
rect 1334 7176 261600 7784
rect 1334 7036 261560 7176
rect 1334 6428 261600 7036
rect 1334 6288 261560 6428
rect 1334 5680 261600 6288
rect 1334 5540 261560 5680
rect 1334 4932 261600 5540
rect 1334 4792 261560 4932
rect 1334 4184 261600 4792
rect 1334 4044 261560 4184
rect 1334 3436 261600 4044
rect 1334 3296 261560 3436
rect 1334 2688 261600 3296
rect 1334 2548 261560 2688
rect 1334 1940 261600 2548
rect 1334 1800 261560 1940
rect 1334 1192 261600 1800
rect 1334 1052 261560 1192
rect 1334 444 261600 1052
rect 1334 357 261560 444
<< obsm4 >>
rect 502 697 259460 74906
<< metal5 >>
rect 552 78428 261418 78748
rect 552 71928 1100 72248
rect 54900 71928 60100 72248
rect 258900 71928 261418 72248
rect 552 65428 1100 65748
rect 54900 65428 60100 65748
rect 258900 65428 261418 65748
rect 552 58928 1100 59248
rect 54900 58928 60100 59248
rect 258900 58928 261418 59248
rect 552 52428 1100 52748
rect 54900 52428 60100 52748
rect 258900 52428 261418 52748
rect 552 45928 1100 46248
rect 54900 45928 60100 46248
rect 258900 45928 261418 46248
rect 552 39428 1100 39748
rect 54900 39428 60100 39748
rect 258900 39428 261418 39748
rect 552 32928 1100 33248
rect 54900 32928 60100 33248
rect 258900 32928 261418 33248
rect 552 26428 1100 26748
rect 54900 26428 60100 26748
rect 258900 26428 261418 26748
rect 552 19928 1100 20248
rect 54900 19928 60100 20248
rect 258900 19928 261418 20248
rect 552 13428 1100 13748
rect 54900 13428 60100 13748
rect 258900 13428 261418 13748
rect 552 6928 1100 7248
rect 54900 6928 60100 7248
rect 258900 6928 261418 7248
<< obsm5 >>
rect 502 72408 259460 74906
rect 1260 71768 54740 72408
rect 60260 71768 258740 72408
rect 502 65908 259460 71768
rect 1260 65268 54740 65908
rect 60260 65268 258740 65908
rect 502 59408 259460 65268
rect 1260 58768 54740 59408
rect 60260 58768 258740 59408
rect 502 52908 259460 58768
rect 1260 52268 54740 52908
rect 60260 52268 258740 52908
rect 502 46408 259460 52268
rect 1260 45768 54740 46408
rect 60260 45768 258740 46408
rect 502 39908 259460 45768
rect 1260 39268 54740 39908
rect 60260 39268 258740 39908
rect 502 33408 259460 39268
rect 1260 32768 54740 33408
rect 60260 32768 258740 33408
rect 502 26908 259460 32768
rect 1260 26268 54740 26908
rect 60260 26268 258740 26908
rect 502 20408 259460 26268
rect 1260 19768 54740 20408
rect 60260 19768 258740 20408
rect 502 13908 259460 19768
rect 1260 13268 54740 13908
rect 60260 13268 258740 13908
rect 502 7408 259460 13268
rect 1260 6768 54740 7408
rect 60260 6768 258740 7408
rect 502 1078 259460 6768
<< labels >>
rlabel metal5 s 552 13428 1100 13748 6 VGND
port 1 nsew ground input
rlabel metal5 s 54900 13428 60100 13748 6 VGND
port 1 nsew ground input
rlabel metal5 s 258900 13428 261418 13748 6 VGND
port 1 nsew ground input
rlabel metal5 s 552 26428 1100 26748 6 VGND
port 1 nsew ground input
rlabel metal5 s 54900 26428 60100 26748 6 VGND
port 1 nsew ground input
rlabel metal5 s 258900 26428 261418 26748 6 VGND
port 1 nsew ground input
rlabel metal5 s 552 39428 1100 39748 6 VGND
port 1 nsew ground input
rlabel metal5 s 54900 39428 60100 39748 6 VGND
port 1 nsew ground input
rlabel metal5 s 258900 39428 261418 39748 6 VGND
port 1 nsew ground input
rlabel metal5 s 552 52428 1100 52748 6 VGND
port 1 nsew ground input
rlabel metal5 s 54900 52428 60100 52748 6 VGND
port 1 nsew ground input
rlabel metal5 s 258900 52428 261418 52748 6 VGND
port 1 nsew ground input
rlabel metal5 s 552 65428 1100 65748 6 VGND
port 1 nsew ground input
rlabel metal5 s 54900 65428 60100 65748 6 VGND
port 1 nsew ground input
rlabel metal5 s 258900 65428 261418 65748 6 VGND
port 1 nsew ground input
rlabel metal5 s 552 78428 261418 78748 6 VGND
port 1 nsew ground input
rlabel metal5 s 552 6928 1100 7248 6 VPWR
port 2 nsew power input
rlabel metal5 s 54900 6928 60100 7248 6 VPWR
port 2 nsew power input
rlabel metal5 s 258900 6928 261418 7248 6 VPWR
port 2 nsew power input
rlabel metal5 s 552 19928 1100 20248 6 VPWR
port 2 nsew power input
rlabel metal5 s 54900 19928 60100 20248 6 VPWR
port 2 nsew power input
rlabel metal5 s 258900 19928 261418 20248 6 VPWR
port 2 nsew power input
rlabel metal5 s 552 32928 1100 33248 6 VPWR
port 2 nsew power input
rlabel metal5 s 54900 32928 60100 33248 6 VPWR
port 2 nsew power input
rlabel metal5 s 258900 32928 261418 33248 6 VPWR
port 2 nsew power input
rlabel metal5 s 552 45928 1100 46248 6 VPWR
port 2 nsew power input
rlabel metal5 s 54900 45928 60100 46248 6 VPWR
port 2 nsew power input
rlabel metal5 s 258900 45928 261418 46248 6 VPWR
port 2 nsew power input
rlabel metal5 s 552 58928 1100 59248 6 VPWR
port 2 nsew power input
rlabel metal5 s 54900 58928 60100 59248 6 VPWR
port 2 nsew power input
rlabel metal5 s 258900 58928 261418 59248 6 VPWR
port 2 nsew power input
rlabel metal5 s 552 71928 1100 72248 6 VPWR
port 2 nsew power input
rlabel metal5 s 54900 71928 60100 72248 6 VPWR
port 2 nsew power input
rlabel metal5 s 258900 71928 261418 72248 6 VPWR
port 2 nsew power input
rlabel metal2 s 147393 -200 147421 400 6 core_clk
port 3 nsew signal input
rlabel metal2 s 49137 -200 49165 400 6 core_rstn
port 4 nsew signal input
rlabel metal3 s 261600 31896 262200 31956 6 debug_in
port 5 nsew signal input
rlabel metal3 s 261600 32644 262200 32704 6 debug_mode
port 6 nsew signal output
rlabel metal3 s 261600 33392 262200 33452 6 debug_oeb
port 7 nsew signal output
rlabel metal3 s 261600 34140 262200 34200 6 debug_out
port 8 nsew signal output
rlabel metal3 s 261600 72560 262200 72620 6 flash_clk
port 9 nsew signal output
rlabel metal3 s 261600 71812 262200 71872 6 flash_csb
port 10 nsew signal output
rlabel metal3 s 261600 73308 262200 73368 6 flash_io0_di
port 11 nsew signal input
rlabel metal3 s 261600 74056 262200 74116 6 flash_io0_do
port 12 nsew signal output
rlabel metal3 s 261600 74804 262200 74864 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal3 s 261600 75552 262200 75612 6 flash_io1_di
port 14 nsew signal input
rlabel metal3 s 261600 76300 262200 76360 6 flash_io1_do
port 15 nsew signal output
rlabel metal3 s 261600 77048 262200 77108 6 flash_io1_oeb
port 16 nsew signal output
rlabel metal3 s 261600 77796 262200 77856 6 flash_io2_di
port 17 nsew signal input
rlabel metal3 s 261600 78544 262200 78604 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 261600 79292 262200 79352 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal3 s 261600 80040 262200 80100 6 flash_io3_di
port 20 nsew signal input
rlabel metal3 s 261600 80788 262200 80848 6 flash_io3_do
port 21 nsew signal output
rlabel metal3 s 261600 81536 262200 81596 6 flash_io3_oeb
port 22 nsew signal output
rlabel metal2 s 16385 -200 16413 400 6 gpio_in_pad
port 23 nsew signal input
rlabel metal2 s 81889 -200 81917 400 6 gpio_inenb_pad
port 24 nsew signal output
rlabel metal2 s 114641 -200 114669 400 6 gpio_mode0_pad
port 25 nsew signal output
rlabel metal2 s 180145 -200 180173 400 6 gpio_mode1_pad
port 26 nsew signal output
rlabel metal2 s 212897 -200 212925 400 6 gpio_out_pad
port 27 nsew signal output
rlabel metal2 s 245649 -200 245677 400 6 gpio_outenb_pad
port 28 nsew signal output
rlabel metal3 s 261600 45428 262200 45488 6 hk_ack_i
port 29 nsew signal input
rlabel metal3 s 261600 46924 262200 46984 6 hk_cyc_o
port 30 nsew signal output
rlabel metal3 s 261600 47740 262200 47800 6 hk_dat_i[0]
port 31 nsew signal input
rlabel metal3 s 261600 55220 262200 55280 6 hk_dat_i[10]
port 32 nsew signal input
rlabel metal3 s 261600 55968 262200 56028 6 hk_dat_i[11]
port 33 nsew signal input
rlabel metal3 s 261600 56716 262200 56776 6 hk_dat_i[12]
port 34 nsew signal input
rlabel metal3 s 261600 57464 262200 57524 6 hk_dat_i[13]
port 35 nsew signal input
rlabel metal3 s 261600 58212 262200 58272 6 hk_dat_i[14]
port 36 nsew signal input
rlabel metal3 s 261600 59028 262200 59088 6 hk_dat_i[15]
port 37 nsew signal input
rlabel metal3 s 261600 59776 262200 59836 6 hk_dat_i[16]
port 38 nsew signal input
rlabel metal3 s 261600 60524 262200 60584 6 hk_dat_i[17]
port 39 nsew signal input
rlabel metal3 s 261600 61272 262200 61332 6 hk_dat_i[18]
port 40 nsew signal input
rlabel metal3 s 261600 62020 262200 62080 6 hk_dat_i[19]
port 41 nsew signal input
rlabel metal3 s 261600 48488 262200 48548 6 hk_dat_i[1]
port 42 nsew signal input
rlabel metal3 s 261600 62768 262200 62828 6 hk_dat_i[20]
port 43 nsew signal input
rlabel metal3 s 261600 63516 262200 63576 6 hk_dat_i[21]
port 44 nsew signal input
rlabel metal3 s 261600 64264 262200 64324 6 hk_dat_i[22]
port 45 nsew signal input
rlabel metal3 s 261600 65012 262200 65072 6 hk_dat_i[23]
port 46 nsew signal input
rlabel metal3 s 261600 65760 262200 65820 6 hk_dat_i[24]
port 47 nsew signal input
rlabel metal3 s 261600 66508 262200 66568 6 hk_dat_i[25]
port 48 nsew signal input
rlabel metal3 s 261600 67256 262200 67316 6 hk_dat_i[26]
port 49 nsew signal input
rlabel metal3 s 261600 68004 262200 68064 6 hk_dat_i[27]
port 50 nsew signal input
rlabel metal3 s 261600 68752 262200 68812 6 hk_dat_i[28]
port 51 nsew signal input
rlabel metal3 s 261600 69500 262200 69560 6 hk_dat_i[29]
port 52 nsew signal input
rlabel metal3 s 261600 49236 262200 49296 6 hk_dat_i[2]
port 53 nsew signal input
rlabel metal3 s 261600 70248 262200 70308 6 hk_dat_i[30]
port 54 nsew signal input
rlabel metal3 s 261600 71064 262200 71124 6 hk_dat_i[31]
port 55 nsew signal input
rlabel metal3 s 261600 49984 262200 50044 6 hk_dat_i[3]
port 56 nsew signal input
rlabel metal3 s 261600 50732 262200 50792 6 hk_dat_i[4]
port 57 nsew signal input
rlabel metal3 s 261600 51480 262200 51540 6 hk_dat_i[5]
port 58 nsew signal input
rlabel metal3 s 261600 52228 262200 52288 6 hk_dat_i[6]
port 59 nsew signal input
rlabel metal3 s 261600 52976 262200 53036 6 hk_dat_i[7]
port 60 nsew signal input
rlabel metal3 s 261600 53724 262200 53784 6 hk_dat_i[8]
port 61 nsew signal input
rlabel metal3 s 261600 54472 262200 54532 6 hk_dat_i[9]
port 62 nsew signal input
rlabel metal3 s 261600 46176 262200 46236 6 hk_stb_o
port 63 nsew signal output
rlabel metal2 s 260921 81600 260949 82200 6 irq[0]
port 64 nsew signal input
rlabel metal2 s 261335 81600 261363 82200 6 irq[1]
port 65 nsew signal input
rlabel metal2 s 261749 81600 261777 82200 6 irq[2]
port 66 nsew signal input
rlabel metal3 s 261600 37200 262200 37260 6 irq[3]
port 67 nsew signal input
rlabel metal3 s 261600 36452 262200 36512 6 irq[4]
port 68 nsew signal input
rlabel metal3 s 261600 35704 262200 35764 6 irq[5]
port 69 nsew signal input
rlabel metal2 s 193 81600 221 82200 6 la_iena[0]
port 70 nsew signal output
rlabel metal2 s 168415 81600 168443 82200 6 la_iena[100]
port 71 nsew signal output
rlabel metal2 s 170071 81600 170099 82200 6 la_iena[101]
port 72 nsew signal output
rlabel metal2 s 171773 81600 171801 82200 6 la_iena[102]
port 73 nsew signal output
rlabel metal2 s 173429 81600 173457 82200 6 la_iena[103]
port 74 nsew signal output
rlabel metal2 s 175131 81600 175159 82200 6 la_iena[104]
port 75 nsew signal output
rlabel metal2 s 176833 81600 176861 82200 6 la_iena[105]
port 76 nsew signal output
rlabel metal2 s 178489 81600 178517 82200 6 la_iena[106]
port 77 nsew signal output
rlabel metal2 s 180191 81600 180219 82200 6 la_iena[107]
port 78 nsew signal output
rlabel metal2 s 181847 81600 181875 82200 6 la_iena[108]
port 79 nsew signal output
rlabel metal2 s 183549 81600 183577 82200 6 la_iena[109]
port 80 nsew signal output
rlabel metal2 s 16983 81600 17011 82200 6 la_iena[10]
port 81 nsew signal output
rlabel metal2 s 185205 81600 185233 82200 6 la_iena[110]
port 82 nsew signal output
rlabel metal2 s 186907 81600 186935 82200 6 la_iena[111]
port 83 nsew signal output
rlabel metal2 s 188609 81600 188637 82200 6 la_iena[112]
port 84 nsew signal output
rlabel metal2 s 190265 81600 190293 82200 6 la_iena[113]
port 85 nsew signal output
rlabel metal2 s 191967 81600 191995 82200 6 la_iena[114]
port 86 nsew signal output
rlabel metal2 s 193623 81600 193651 82200 6 la_iena[115]
port 87 nsew signal output
rlabel metal2 s 195325 81600 195353 82200 6 la_iena[116]
port 88 nsew signal output
rlabel metal2 s 196981 81600 197009 82200 6 la_iena[117]
port 89 nsew signal output
rlabel metal2 s 198683 81600 198711 82200 6 la_iena[118]
port 90 nsew signal output
rlabel metal2 s 200385 81600 200413 82200 6 la_iena[119]
port 91 nsew signal output
rlabel metal2 s 18685 81600 18713 82200 6 la_iena[11]
port 92 nsew signal output
rlabel metal2 s 202041 81600 202069 82200 6 la_iena[120]
port 93 nsew signal output
rlabel metal2 s 203743 81600 203771 82200 6 la_iena[121]
port 94 nsew signal output
rlabel metal2 s 205399 81600 205427 82200 6 la_iena[122]
port 95 nsew signal output
rlabel metal2 s 207101 81600 207129 82200 6 la_iena[123]
port 96 nsew signal output
rlabel metal2 s 208757 81600 208785 82200 6 la_iena[124]
port 97 nsew signal output
rlabel metal2 s 210459 81600 210487 82200 6 la_iena[125]
port 98 nsew signal output
rlabel metal2 s 212161 81600 212189 82200 6 la_iena[126]
port 99 nsew signal output
rlabel metal2 s 213817 81600 213845 82200 6 la_iena[127]
port 100 nsew signal output
rlabel metal2 s 20341 81600 20369 82200 6 la_iena[12]
port 101 nsew signal output
rlabel metal2 s 22043 81600 22071 82200 6 la_iena[13]
port 102 nsew signal output
rlabel metal2 s 23745 81600 23773 82200 6 la_iena[14]
port 103 nsew signal output
rlabel metal2 s 25401 81600 25429 82200 6 la_iena[15]
port 104 nsew signal output
rlabel metal2 s 27103 81600 27131 82200 6 la_iena[16]
port 105 nsew signal output
rlabel metal2 s 28759 81600 28787 82200 6 la_iena[17]
port 106 nsew signal output
rlabel metal2 s 30461 81600 30489 82200 6 la_iena[18]
port 107 nsew signal output
rlabel metal2 s 32117 81600 32145 82200 6 la_iena[19]
port 108 nsew signal output
rlabel metal2 s 1849 81600 1877 82200 6 la_iena[1]
port 109 nsew signal output
rlabel metal2 s 33819 81600 33847 82200 6 la_iena[20]
port 110 nsew signal output
rlabel metal2 s 35521 81600 35549 82200 6 la_iena[21]
port 111 nsew signal output
rlabel metal2 s 37177 81600 37205 82200 6 la_iena[22]
port 112 nsew signal output
rlabel metal2 s 38879 81600 38907 82200 6 la_iena[23]
port 113 nsew signal output
rlabel metal2 s 40535 81600 40563 82200 6 la_iena[24]
port 114 nsew signal output
rlabel metal2 s 42237 81600 42265 82200 6 la_iena[25]
port 115 nsew signal output
rlabel metal2 s 43893 81600 43921 82200 6 la_iena[26]
port 116 nsew signal output
rlabel metal2 s 45595 81600 45623 82200 6 la_iena[27]
port 117 nsew signal output
rlabel metal2 s 47297 81600 47325 82200 6 la_iena[28]
port 118 nsew signal output
rlabel metal2 s 48953 81600 48981 82200 6 la_iena[29]
port 119 nsew signal output
rlabel metal2 s 3551 81600 3579 82200 6 la_iena[2]
port 120 nsew signal output
rlabel metal2 s 50655 81600 50683 82200 6 la_iena[30]
port 121 nsew signal output
rlabel metal2 s 52311 81600 52339 82200 6 la_iena[31]
port 122 nsew signal output
rlabel metal2 s 54013 81600 54041 82200 6 la_iena[32]
port 123 nsew signal output
rlabel metal2 s 55669 81600 55697 82200 6 la_iena[33]
port 124 nsew signal output
rlabel metal2 s 57371 81600 57399 82200 6 la_iena[34]
port 125 nsew signal output
rlabel metal2 s 59073 81600 59101 82200 6 la_iena[35]
port 126 nsew signal output
rlabel metal2 s 60729 81600 60757 82200 6 la_iena[36]
port 127 nsew signal output
rlabel metal2 s 62431 81600 62459 82200 6 la_iena[37]
port 128 nsew signal output
rlabel metal2 s 64087 81600 64115 82200 6 la_iena[38]
port 129 nsew signal output
rlabel metal2 s 65789 81600 65817 82200 6 la_iena[39]
port 130 nsew signal output
rlabel metal2 s 5207 81600 5235 82200 6 la_iena[3]
port 131 nsew signal output
rlabel metal2 s 67445 81600 67473 82200 6 la_iena[40]
port 132 nsew signal output
rlabel metal2 s 69147 81600 69175 82200 6 la_iena[41]
port 133 nsew signal output
rlabel metal2 s 70849 81600 70877 82200 6 la_iena[42]
port 134 nsew signal output
rlabel metal2 s 72505 81600 72533 82200 6 la_iena[43]
port 135 nsew signal output
rlabel metal2 s 74207 81600 74235 82200 6 la_iena[44]
port 136 nsew signal output
rlabel metal2 s 75863 81600 75891 82200 6 la_iena[45]
port 137 nsew signal output
rlabel metal2 s 77565 81600 77593 82200 6 la_iena[46]
port 138 nsew signal output
rlabel metal2 s 79221 81600 79249 82200 6 la_iena[47]
port 139 nsew signal output
rlabel metal2 s 80923 81600 80951 82200 6 la_iena[48]
port 140 nsew signal output
rlabel metal2 s 82625 81600 82653 82200 6 la_iena[49]
port 141 nsew signal output
rlabel metal2 s 6909 81600 6937 82200 6 la_iena[4]
port 142 nsew signal output
rlabel metal2 s 84281 81600 84309 82200 6 la_iena[50]
port 143 nsew signal output
rlabel metal2 s 85983 81600 86011 82200 6 la_iena[51]
port 144 nsew signal output
rlabel metal2 s 87639 81600 87667 82200 6 la_iena[52]
port 145 nsew signal output
rlabel metal2 s 89341 81600 89369 82200 6 la_iena[53]
port 146 nsew signal output
rlabel metal2 s 90997 81600 91025 82200 6 la_iena[54]
port 147 nsew signal output
rlabel metal2 s 92699 81600 92727 82200 6 la_iena[55]
port 148 nsew signal output
rlabel metal2 s 94401 81600 94429 82200 6 la_iena[56]
port 149 nsew signal output
rlabel metal2 s 96057 81600 96085 82200 6 la_iena[57]
port 150 nsew signal output
rlabel metal2 s 97759 81600 97787 82200 6 la_iena[58]
port 151 nsew signal output
rlabel metal2 s 99415 81600 99443 82200 6 la_iena[59]
port 152 nsew signal output
rlabel metal2 s 8565 81600 8593 82200 6 la_iena[5]
port 153 nsew signal output
rlabel metal2 s 101117 81600 101145 82200 6 la_iena[60]
port 154 nsew signal output
rlabel metal2 s 102773 81600 102801 82200 6 la_iena[61]
port 155 nsew signal output
rlabel metal2 s 104475 81600 104503 82200 6 la_iena[62]
port 156 nsew signal output
rlabel metal2 s 106177 81600 106205 82200 6 la_iena[63]
port 157 nsew signal output
rlabel metal2 s 107833 81600 107861 82200 6 la_iena[64]
port 158 nsew signal output
rlabel metal2 s 109535 81600 109563 82200 6 la_iena[65]
port 159 nsew signal output
rlabel metal2 s 111191 81600 111219 82200 6 la_iena[66]
port 160 nsew signal output
rlabel metal2 s 112893 81600 112921 82200 6 la_iena[67]
port 161 nsew signal output
rlabel metal2 s 114549 81600 114577 82200 6 la_iena[68]
port 162 nsew signal output
rlabel metal2 s 116251 81600 116279 82200 6 la_iena[69]
port 163 nsew signal output
rlabel metal2 s 10267 81600 10295 82200 6 la_iena[6]
port 164 nsew signal output
rlabel metal2 s 117953 81600 117981 82200 6 la_iena[70]
port 165 nsew signal output
rlabel metal2 s 119609 81600 119637 82200 6 la_iena[71]
port 166 nsew signal output
rlabel metal2 s 121311 81600 121339 82200 6 la_iena[72]
port 167 nsew signal output
rlabel metal2 s 122967 81600 122995 82200 6 la_iena[73]
port 168 nsew signal output
rlabel metal2 s 124669 81600 124697 82200 6 la_iena[74]
port 169 nsew signal output
rlabel metal2 s 126325 81600 126353 82200 6 la_iena[75]
port 170 nsew signal output
rlabel metal2 s 128027 81600 128055 82200 6 la_iena[76]
port 171 nsew signal output
rlabel metal2 s 129729 81600 129757 82200 6 la_iena[77]
port 172 nsew signal output
rlabel metal2 s 131385 81600 131413 82200 6 la_iena[78]
port 173 nsew signal output
rlabel metal2 s 133087 81600 133115 82200 6 la_iena[79]
port 174 nsew signal output
rlabel metal2 s 11969 81600 11997 82200 6 la_iena[7]
port 175 nsew signal output
rlabel metal2 s 134743 81600 134771 82200 6 la_iena[80]
port 176 nsew signal output
rlabel metal2 s 136445 81600 136473 82200 6 la_iena[81]
port 177 nsew signal output
rlabel metal2 s 138101 81600 138129 82200 6 la_iena[82]
port 178 nsew signal output
rlabel metal2 s 139803 81600 139831 82200 6 la_iena[83]
port 179 nsew signal output
rlabel metal2 s 141505 81600 141533 82200 6 la_iena[84]
port 180 nsew signal output
rlabel metal2 s 143161 81600 143189 82200 6 la_iena[85]
port 181 nsew signal output
rlabel metal2 s 144863 81600 144891 82200 6 la_iena[86]
port 182 nsew signal output
rlabel metal2 s 146519 81600 146547 82200 6 la_iena[87]
port 183 nsew signal output
rlabel metal2 s 148221 81600 148249 82200 6 la_iena[88]
port 184 nsew signal output
rlabel metal2 s 149877 81600 149905 82200 6 la_iena[89]
port 185 nsew signal output
rlabel metal2 s 13625 81600 13653 82200 6 la_iena[8]
port 186 nsew signal output
rlabel metal2 s 151579 81600 151607 82200 6 la_iena[90]
port 187 nsew signal output
rlabel metal2 s 153281 81600 153309 82200 6 la_iena[91]
port 188 nsew signal output
rlabel metal2 s 154937 81600 154965 82200 6 la_iena[92]
port 189 nsew signal output
rlabel metal2 s 156639 81600 156667 82200 6 la_iena[93]
port 190 nsew signal output
rlabel metal2 s 158295 81600 158323 82200 6 la_iena[94]
port 191 nsew signal output
rlabel metal2 s 159997 81600 160025 82200 6 la_iena[95]
port 192 nsew signal output
rlabel metal2 s 161653 81600 161681 82200 6 la_iena[96]
port 193 nsew signal output
rlabel metal2 s 163355 81600 163383 82200 6 la_iena[97]
port 194 nsew signal output
rlabel metal2 s 165057 81600 165085 82200 6 la_iena[98]
port 195 nsew signal output
rlabel metal2 s 166713 81600 166741 82200 6 la_iena[99]
port 196 nsew signal output
rlabel metal2 s 15327 81600 15355 82200 6 la_iena[9]
port 197 nsew signal output
rlabel metal2 s 607 81600 635 82200 6 la_input[0]
port 198 nsew signal input
rlabel metal2 s 168829 81600 168857 82200 6 la_input[100]
port 199 nsew signal input
rlabel metal2 s 170485 81600 170513 82200 6 la_input[101]
port 200 nsew signal input
rlabel metal2 s 172187 81600 172215 82200 6 la_input[102]
port 201 nsew signal input
rlabel metal2 s 173889 81600 173917 82200 6 la_input[103]
port 202 nsew signal input
rlabel metal2 s 175545 81600 175573 82200 6 la_input[104]
port 203 nsew signal input
rlabel metal2 s 177247 81600 177275 82200 6 la_input[105]
port 204 nsew signal input
rlabel metal2 s 178903 81600 178931 82200 6 la_input[106]
port 205 nsew signal input
rlabel metal2 s 180605 81600 180633 82200 6 la_input[107]
port 206 nsew signal input
rlabel metal2 s 182261 81600 182289 82200 6 la_input[108]
port 207 nsew signal input
rlabel metal2 s 183963 81600 183991 82200 6 la_input[109]
port 208 nsew signal input
rlabel metal2 s 17397 81600 17425 82200 6 la_input[10]
port 209 nsew signal input
rlabel metal2 s 185665 81600 185693 82200 6 la_input[110]
port 210 nsew signal input
rlabel metal2 s 187321 81600 187349 82200 6 la_input[111]
port 211 nsew signal input
rlabel metal2 s 189023 81600 189051 82200 6 la_input[112]
port 212 nsew signal input
rlabel metal2 s 190679 81600 190707 82200 6 la_input[113]
port 213 nsew signal input
rlabel metal2 s 192381 81600 192409 82200 6 la_input[114]
port 214 nsew signal input
rlabel metal2 s 194037 81600 194065 82200 6 la_input[115]
port 215 nsew signal input
rlabel metal2 s 195739 81600 195767 82200 6 la_input[116]
port 216 nsew signal input
rlabel metal2 s 197441 81600 197469 82200 6 la_input[117]
port 217 nsew signal input
rlabel metal2 s 199097 81600 199125 82200 6 la_input[118]
port 218 nsew signal input
rlabel metal2 s 200799 81600 200827 82200 6 la_input[119]
port 219 nsew signal input
rlabel metal2 s 19099 81600 19127 82200 6 la_input[11]
port 220 nsew signal input
rlabel metal2 s 202455 81600 202483 82200 6 la_input[120]
port 221 nsew signal input
rlabel metal2 s 204157 81600 204185 82200 6 la_input[121]
port 222 nsew signal input
rlabel metal2 s 205813 81600 205841 82200 6 la_input[122]
port 223 nsew signal input
rlabel metal2 s 207515 81600 207543 82200 6 la_input[123]
port 224 nsew signal input
rlabel metal2 s 209217 81600 209245 82200 6 la_input[124]
port 225 nsew signal input
rlabel metal2 s 210873 81600 210901 82200 6 la_input[125]
port 226 nsew signal input
rlabel metal2 s 212575 81600 212603 82200 6 la_input[126]
port 227 nsew signal input
rlabel metal2 s 214231 81600 214259 82200 6 la_input[127]
port 228 nsew signal input
rlabel metal2 s 20801 81600 20829 82200 6 la_input[12]
port 229 nsew signal input
rlabel metal2 s 22457 81600 22485 82200 6 la_input[13]
port 230 nsew signal input
rlabel metal2 s 24159 81600 24187 82200 6 la_input[14]
port 231 nsew signal input
rlabel metal2 s 25815 81600 25843 82200 6 la_input[15]
port 232 nsew signal input
rlabel metal2 s 27517 81600 27545 82200 6 la_input[16]
port 233 nsew signal input
rlabel metal2 s 29173 81600 29201 82200 6 la_input[17]
port 234 nsew signal input
rlabel metal2 s 30875 81600 30903 82200 6 la_input[18]
port 235 nsew signal input
rlabel metal2 s 32577 81600 32605 82200 6 la_input[19]
port 236 nsew signal input
rlabel metal2 s 2263 81600 2291 82200 6 la_input[1]
port 237 nsew signal input
rlabel metal2 s 34233 81600 34261 82200 6 la_input[20]
port 238 nsew signal input
rlabel metal2 s 35935 81600 35963 82200 6 la_input[21]
port 239 nsew signal input
rlabel metal2 s 37591 81600 37619 82200 6 la_input[22]
port 240 nsew signal input
rlabel metal2 s 39293 81600 39321 82200 6 la_input[23]
port 241 nsew signal input
rlabel metal2 s 40949 81600 40977 82200 6 la_input[24]
port 242 nsew signal input
rlabel metal2 s 42651 81600 42679 82200 6 la_input[25]
port 243 nsew signal input
rlabel metal2 s 44353 81600 44381 82200 6 la_input[26]
port 244 nsew signal input
rlabel metal2 s 46009 81600 46037 82200 6 la_input[27]
port 245 nsew signal input
rlabel metal2 s 47711 81600 47739 82200 6 la_input[28]
port 246 nsew signal input
rlabel metal2 s 49367 81600 49395 82200 6 la_input[29]
port 247 nsew signal input
rlabel metal2 s 3965 81600 3993 82200 6 la_input[2]
port 248 nsew signal input
rlabel metal2 s 51069 81600 51097 82200 6 la_input[30]
port 249 nsew signal input
rlabel metal2 s 52725 81600 52753 82200 6 la_input[31]
port 250 nsew signal input
rlabel metal2 s 54427 81600 54455 82200 6 la_input[32]
port 251 nsew signal input
rlabel metal2 s 56129 81600 56157 82200 6 la_input[33]
port 252 nsew signal input
rlabel metal2 s 57785 81600 57813 82200 6 la_input[34]
port 253 nsew signal input
rlabel metal2 s 59487 81600 59515 82200 6 la_input[35]
port 254 nsew signal input
rlabel metal2 s 61143 81600 61171 82200 6 la_input[36]
port 255 nsew signal input
rlabel metal2 s 62845 81600 62873 82200 6 la_input[37]
port 256 nsew signal input
rlabel metal2 s 64501 81600 64529 82200 6 la_input[38]
port 257 nsew signal input
rlabel metal2 s 66203 81600 66231 82200 6 la_input[39]
port 258 nsew signal input
rlabel metal2 s 5621 81600 5649 82200 6 la_input[3]
port 259 nsew signal input
rlabel metal2 s 67905 81600 67933 82200 6 la_input[40]
port 260 nsew signal input
rlabel metal2 s 69561 81600 69589 82200 6 la_input[41]
port 261 nsew signal input
rlabel metal2 s 71263 81600 71291 82200 6 la_input[42]
port 262 nsew signal input
rlabel metal2 s 72919 81600 72947 82200 6 la_input[43]
port 263 nsew signal input
rlabel metal2 s 74621 81600 74649 82200 6 la_input[44]
port 264 nsew signal input
rlabel metal2 s 76277 81600 76305 82200 6 la_input[45]
port 265 nsew signal input
rlabel metal2 s 77979 81600 78007 82200 6 la_input[46]
port 266 nsew signal input
rlabel metal2 s 79681 81600 79709 82200 6 la_input[47]
port 267 nsew signal input
rlabel metal2 s 81337 81600 81365 82200 6 la_input[48]
port 268 nsew signal input
rlabel metal2 s 83039 81600 83067 82200 6 la_input[49]
port 269 nsew signal input
rlabel metal2 s 7323 81600 7351 82200 6 la_input[4]
port 270 nsew signal input
rlabel metal2 s 84695 81600 84723 82200 6 la_input[50]
port 271 nsew signal input
rlabel metal2 s 86397 81600 86425 82200 6 la_input[51]
port 272 nsew signal input
rlabel metal2 s 88053 81600 88081 82200 6 la_input[52]
port 273 nsew signal input
rlabel metal2 s 89755 81600 89783 82200 6 la_input[53]
port 274 nsew signal input
rlabel metal2 s 91457 81600 91485 82200 6 la_input[54]
port 275 nsew signal input
rlabel metal2 s 93113 81600 93141 82200 6 la_input[55]
port 276 nsew signal input
rlabel metal2 s 94815 81600 94843 82200 6 la_input[56]
port 277 nsew signal input
rlabel metal2 s 96471 81600 96499 82200 6 la_input[57]
port 278 nsew signal input
rlabel metal2 s 98173 81600 98201 82200 6 la_input[58]
port 279 nsew signal input
rlabel metal2 s 99829 81600 99857 82200 6 la_input[59]
port 280 nsew signal input
rlabel metal2 s 9025 81600 9053 82200 6 la_input[5]
port 281 nsew signal input
rlabel metal2 s 101531 81600 101559 82200 6 la_input[60]
port 282 nsew signal input
rlabel metal2 s 103233 81600 103261 82200 6 la_input[61]
port 283 nsew signal input
rlabel metal2 s 104889 81600 104917 82200 6 la_input[62]
port 284 nsew signal input
rlabel metal2 s 106591 81600 106619 82200 6 la_input[63]
port 285 nsew signal input
rlabel metal2 s 108247 81600 108275 82200 6 la_input[64]
port 286 nsew signal input
rlabel metal2 s 109949 81600 109977 82200 6 la_input[65]
port 287 nsew signal input
rlabel metal2 s 111605 81600 111633 82200 6 la_input[66]
port 288 nsew signal input
rlabel metal2 s 113307 81600 113335 82200 6 la_input[67]
port 289 nsew signal input
rlabel metal2 s 115009 81600 115037 82200 6 la_input[68]
port 290 nsew signal input
rlabel metal2 s 116665 81600 116693 82200 6 la_input[69]
port 291 nsew signal input
rlabel metal2 s 10681 81600 10709 82200 6 la_input[6]
port 292 nsew signal input
rlabel metal2 s 118367 81600 118395 82200 6 la_input[70]
port 293 nsew signal input
rlabel metal2 s 120023 81600 120051 82200 6 la_input[71]
port 294 nsew signal input
rlabel metal2 s 121725 81600 121753 82200 6 la_input[72]
port 295 nsew signal input
rlabel metal2 s 123381 81600 123409 82200 6 la_input[73]
port 296 nsew signal input
rlabel metal2 s 125083 81600 125111 82200 6 la_input[74]
port 297 nsew signal input
rlabel metal2 s 126785 81600 126813 82200 6 la_input[75]
port 298 nsew signal input
rlabel metal2 s 128441 81600 128469 82200 6 la_input[76]
port 299 nsew signal input
rlabel metal2 s 130143 81600 130171 82200 6 la_input[77]
port 300 nsew signal input
rlabel metal2 s 131799 81600 131827 82200 6 la_input[78]
port 301 nsew signal input
rlabel metal2 s 133501 81600 133529 82200 6 la_input[79]
port 302 nsew signal input
rlabel metal2 s 12383 81600 12411 82200 6 la_input[7]
port 303 nsew signal input
rlabel metal2 s 135157 81600 135185 82200 6 la_input[80]
port 304 nsew signal input
rlabel metal2 s 136859 81600 136887 82200 6 la_input[81]
port 305 nsew signal input
rlabel metal2 s 138561 81600 138589 82200 6 la_input[82]
port 306 nsew signal input
rlabel metal2 s 140217 81600 140245 82200 6 la_input[83]
port 307 nsew signal input
rlabel metal2 s 141919 81600 141947 82200 6 la_input[84]
port 308 nsew signal input
rlabel metal2 s 143575 81600 143603 82200 6 la_input[85]
port 309 nsew signal input
rlabel metal2 s 145277 81600 145305 82200 6 la_input[86]
port 310 nsew signal input
rlabel metal2 s 146933 81600 146961 82200 6 la_input[87]
port 311 nsew signal input
rlabel metal2 s 148635 81600 148663 82200 6 la_input[88]
port 312 nsew signal input
rlabel metal2 s 150337 81600 150365 82200 6 la_input[89]
port 313 nsew signal input
rlabel metal2 s 14039 81600 14067 82200 6 la_input[8]
port 314 nsew signal input
rlabel metal2 s 151993 81600 152021 82200 6 la_input[90]
port 315 nsew signal input
rlabel metal2 s 153695 81600 153723 82200 6 la_input[91]
port 316 nsew signal input
rlabel metal2 s 155351 81600 155379 82200 6 la_input[92]
port 317 nsew signal input
rlabel metal2 s 157053 81600 157081 82200 6 la_input[93]
port 318 nsew signal input
rlabel metal2 s 158709 81600 158737 82200 6 la_input[94]
port 319 nsew signal input
rlabel metal2 s 160411 81600 160439 82200 6 la_input[95]
port 320 nsew signal input
rlabel metal2 s 162113 81600 162141 82200 6 la_input[96]
port 321 nsew signal input
rlabel metal2 s 163769 81600 163797 82200 6 la_input[97]
port 322 nsew signal input
rlabel metal2 s 165471 81600 165499 82200 6 la_input[98]
port 323 nsew signal input
rlabel metal2 s 167127 81600 167155 82200 6 la_input[99]
port 324 nsew signal input
rlabel metal2 s 15741 81600 15769 82200 6 la_input[9]
port 325 nsew signal input
rlabel metal2 s 1021 81600 1049 82200 6 la_oenb[0]
port 326 nsew signal output
rlabel metal2 s 169243 81600 169271 82200 6 la_oenb[100]
port 327 nsew signal output
rlabel metal2 s 170945 81600 170973 82200 6 la_oenb[101]
port 328 nsew signal output
rlabel metal2 s 172601 81600 172629 82200 6 la_oenb[102]
port 329 nsew signal output
rlabel metal2 s 174303 81600 174331 82200 6 la_oenb[103]
port 330 nsew signal output
rlabel metal2 s 175959 81600 175987 82200 6 la_oenb[104]
port 331 nsew signal output
rlabel metal2 s 177661 81600 177689 82200 6 la_oenb[105]
port 332 nsew signal output
rlabel metal2 s 179317 81600 179345 82200 6 la_oenb[106]
port 333 nsew signal output
rlabel metal2 s 181019 81600 181047 82200 6 la_oenb[107]
port 334 nsew signal output
rlabel metal2 s 182721 81600 182749 82200 6 la_oenb[108]
port 335 nsew signal output
rlabel metal2 s 184377 81600 184405 82200 6 la_oenb[109]
port 336 nsew signal output
rlabel metal2 s 17857 81600 17885 82200 6 la_oenb[10]
port 337 nsew signal output
rlabel metal2 s 186079 81600 186107 82200 6 la_oenb[110]
port 338 nsew signal output
rlabel metal2 s 187735 81600 187763 82200 6 la_oenb[111]
port 339 nsew signal output
rlabel metal2 s 189437 81600 189465 82200 6 la_oenb[112]
port 340 nsew signal output
rlabel metal2 s 191093 81600 191121 82200 6 la_oenb[113]
port 341 nsew signal output
rlabel metal2 s 192795 81600 192823 82200 6 la_oenb[114]
port 342 nsew signal output
rlabel metal2 s 194497 81600 194525 82200 6 la_oenb[115]
port 343 nsew signal output
rlabel metal2 s 196153 81600 196181 82200 6 la_oenb[116]
port 344 nsew signal output
rlabel metal2 s 197855 81600 197883 82200 6 la_oenb[117]
port 345 nsew signal output
rlabel metal2 s 199511 81600 199539 82200 6 la_oenb[118]
port 346 nsew signal output
rlabel metal2 s 201213 81600 201241 82200 6 la_oenb[119]
port 347 nsew signal output
rlabel metal2 s 19513 81600 19541 82200 6 la_oenb[11]
port 348 nsew signal output
rlabel metal2 s 202869 81600 202897 82200 6 la_oenb[120]
port 349 nsew signal output
rlabel metal2 s 204571 81600 204599 82200 6 la_oenb[121]
port 350 nsew signal output
rlabel metal2 s 206273 81600 206301 82200 6 la_oenb[122]
port 351 nsew signal output
rlabel metal2 s 207929 81600 207957 82200 6 la_oenb[123]
port 352 nsew signal output
rlabel metal2 s 209631 81600 209659 82200 6 la_oenb[124]
port 353 nsew signal output
rlabel metal2 s 211287 81600 211315 82200 6 la_oenb[125]
port 354 nsew signal output
rlabel metal2 s 212989 81600 213017 82200 6 la_oenb[126]
port 355 nsew signal output
rlabel metal2 s 214645 81600 214673 82200 6 la_oenb[127]
port 356 nsew signal output
rlabel metal2 s 21215 81600 21243 82200 6 la_oenb[12]
port 357 nsew signal output
rlabel metal2 s 22871 81600 22899 82200 6 la_oenb[13]
port 358 nsew signal output
rlabel metal2 s 24573 81600 24601 82200 6 la_oenb[14]
port 359 nsew signal output
rlabel metal2 s 26229 81600 26257 82200 6 la_oenb[15]
port 360 nsew signal output
rlabel metal2 s 27931 81600 27959 82200 6 la_oenb[16]
port 361 nsew signal output
rlabel metal2 s 29633 81600 29661 82200 6 la_oenb[17]
port 362 nsew signal output
rlabel metal2 s 31289 81600 31317 82200 6 la_oenb[18]
port 363 nsew signal output
rlabel metal2 s 32991 81600 33019 82200 6 la_oenb[19]
port 364 nsew signal output
rlabel metal2 s 2677 81600 2705 82200 6 la_oenb[1]
port 365 nsew signal output
rlabel metal2 s 34647 81600 34675 82200 6 la_oenb[20]
port 366 nsew signal output
rlabel metal2 s 36349 81600 36377 82200 6 la_oenb[21]
port 367 nsew signal output
rlabel metal2 s 38005 81600 38033 82200 6 la_oenb[22]
port 368 nsew signal output
rlabel metal2 s 39707 81600 39735 82200 6 la_oenb[23]
port 369 nsew signal output
rlabel metal2 s 41409 81600 41437 82200 6 la_oenb[24]
port 370 nsew signal output
rlabel metal2 s 43065 81600 43093 82200 6 la_oenb[25]
port 371 nsew signal output
rlabel metal2 s 44767 81600 44795 82200 6 la_oenb[26]
port 372 nsew signal output
rlabel metal2 s 46423 81600 46451 82200 6 la_oenb[27]
port 373 nsew signal output
rlabel metal2 s 48125 81600 48153 82200 6 la_oenb[28]
port 374 nsew signal output
rlabel metal2 s 49781 81600 49809 82200 6 la_oenb[29]
port 375 nsew signal output
rlabel metal2 s 4379 81600 4407 82200 6 la_oenb[2]
port 376 nsew signal output
rlabel metal2 s 51483 81600 51511 82200 6 la_oenb[30]
port 377 nsew signal output
rlabel metal2 s 53185 81600 53213 82200 6 la_oenb[31]
port 378 nsew signal output
rlabel metal2 s 54841 81600 54869 82200 6 la_oenb[32]
port 379 nsew signal output
rlabel metal2 s 56543 81600 56571 82200 6 la_oenb[33]
port 380 nsew signal output
rlabel metal2 s 58199 81600 58227 82200 6 la_oenb[34]
port 381 nsew signal output
rlabel metal2 s 59901 81600 59929 82200 6 la_oenb[35]
port 382 nsew signal output
rlabel metal2 s 61557 81600 61585 82200 6 la_oenb[36]
port 383 nsew signal output
rlabel metal2 s 63259 81600 63287 82200 6 la_oenb[37]
port 384 nsew signal output
rlabel metal2 s 64961 81600 64989 82200 6 la_oenb[38]
port 385 nsew signal output
rlabel metal2 s 66617 81600 66645 82200 6 la_oenb[39]
port 386 nsew signal output
rlabel metal2 s 6081 81600 6109 82200 6 la_oenb[3]
port 387 nsew signal output
rlabel metal2 s 68319 81600 68347 82200 6 la_oenb[40]
port 388 nsew signal output
rlabel metal2 s 69975 81600 70003 82200 6 la_oenb[41]
port 389 nsew signal output
rlabel metal2 s 71677 81600 71705 82200 6 la_oenb[42]
port 390 nsew signal output
rlabel metal2 s 73333 81600 73361 82200 6 la_oenb[43]
port 391 nsew signal output
rlabel metal2 s 75035 81600 75063 82200 6 la_oenb[44]
port 392 nsew signal output
rlabel metal2 s 76737 81600 76765 82200 6 la_oenb[45]
port 393 nsew signal output
rlabel metal2 s 78393 81600 78421 82200 6 la_oenb[46]
port 394 nsew signal output
rlabel metal2 s 80095 81600 80123 82200 6 la_oenb[47]
port 395 nsew signal output
rlabel metal2 s 81751 81600 81779 82200 6 la_oenb[48]
port 396 nsew signal output
rlabel metal2 s 83453 81600 83481 82200 6 la_oenb[49]
port 397 nsew signal output
rlabel metal2 s 7737 81600 7765 82200 6 la_oenb[4]
port 398 nsew signal output
rlabel metal2 s 85109 81600 85137 82200 6 la_oenb[50]
port 399 nsew signal output
rlabel metal2 s 86811 81600 86839 82200 6 la_oenb[51]
port 400 nsew signal output
rlabel metal2 s 88513 81600 88541 82200 6 la_oenb[52]
port 401 nsew signal output
rlabel metal2 s 90169 81600 90197 82200 6 la_oenb[53]
port 402 nsew signal output
rlabel metal2 s 91871 81600 91899 82200 6 la_oenb[54]
port 403 nsew signal output
rlabel metal2 s 93527 81600 93555 82200 6 la_oenb[55]
port 404 nsew signal output
rlabel metal2 s 95229 81600 95257 82200 6 la_oenb[56]
port 405 nsew signal output
rlabel metal2 s 96885 81600 96913 82200 6 la_oenb[57]
port 406 nsew signal output
rlabel metal2 s 98587 81600 98615 82200 6 la_oenb[58]
port 407 nsew signal output
rlabel metal2 s 100289 81600 100317 82200 6 la_oenb[59]
port 408 nsew signal output
rlabel metal2 s 9439 81600 9467 82200 6 la_oenb[5]
port 409 nsew signal output
rlabel metal2 s 101945 81600 101973 82200 6 la_oenb[60]
port 410 nsew signal output
rlabel metal2 s 103647 81600 103675 82200 6 la_oenb[61]
port 411 nsew signal output
rlabel metal2 s 105303 81600 105331 82200 6 la_oenb[62]
port 412 nsew signal output
rlabel metal2 s 107005 81600 107033 82200 6 la_oenb[63]
port 413 nsew signal output
rlabel metal2 s 108661 81600 108689 82200 6 la_oenb[64]
port 414 nsew signal output
rlabel metal2 s 110363 81600 110391 82200 6 la_oenb[65]
port 415 nsew signal output
rlabel metal2 s 112065 81600 112093 82200 6 la_oenb[66]
port 416 nsew signal output
rlabel metal2 s 113721 81600 113749 82200 6 la_oenb[67]
port 417 nsew signal output
rlabel metal2 s 115423 81600 115451 82200 6 la_oenb[68]
port 418 nsew signal output
rlabel metal2 s 117079 81600 117107 82200 6 la_oenb[69]
port 419 nsew signal output
rlabel metal2 s 11095 81600 11123 82200 6 la_oenb[6]
port 420 nsew signal output
rlabel metal2 s 118781 81600 118809 82200 6 la_oenb[70]
port 421 nsew signal output
rlabel metal2 s 120437 81600 120465 82200 6 la_oenb[71]
port 422 nsew signal output
rlabel metal2 s 122139 81600 122167 82200 6 la_oenb[72]
port 423 nsew signal output
rlabel metal2 s 123841 81600 123869 82200 6 la_oenb[73]
port 424 nsew signal output
rlabel metal2 s 125497 81600 125525 82200 6 la_oenb[74]
port 425 nsew signal output
rlabel metal2 s 127199 81600 127227 82200 6 la_oenb[75]
port 426 nsew signal output
rlabel metal2 s 128855 81600 128883 82200 6 la_oenb[76]
port 427 nsew signal output
rlabel metal2 s 130557 81600 130585 82200 6 la_oenb[77]
port 428 nsew signal output
rlabel metal2 s 132213 81600 132241 82200 6 la_oenb[78]
port 429 nsew signal output
rlabel metal2 s 133915 81600 133943 82200 6 la_oenb[79]
port 430 nsew signal output
rlabel metal2 s 12797 81600 12825 82200 6 la_oenb[7]
port 431 nsew signal output
rlabel metal2 s 135617 81600 135645 82200 6 la_oenb[80]
port 432 nsew signal output
rlabel metal2 s 137273 81600 137301 82200 6 la_oenb[81]
port 433 nsew signal output
rlabel metal2 s 138975 81600 139003 82200 6 la_oenb[82]
port 434 nsew signal output
rlabel metal2 s 140631 81600 140659 82200 6 la_oenb[83]
port 435 nsew signal output
rlabel metal2 s 142333 81600 142361 82200 6 la_oenb[84]
port 436 nsew signal output
rlabel metal2 s 143989 81600 144017 82200 6 la_oenb[85]
port 437 nsew signal output
rlabel metal2 s 145691 81600 145719 82200 6 la_oenb[86]
port 438 nsew signal output
rlabel metal2 s 147393 81600 147421 82200 6 la_oenb[87]
port 439 nsew signal output
rlabel metal2 s 149049 81600 149077 82200 6 la_oenb[88]
port 440 nsew signal output
rlabel metal2 s 150751 81600 150779 82200 6 la_oenb[89]
port 441 nsew signal output
rlabel metal2 s 14453 81600 14481 82200 6 la_oenb[8]
port 442 nsew signal output
rlabel metal2 s 152407 81600 152435 82200 6 la_oenb[90]
port 443 nsew signal output
rlabel metal2 s 154109 81600 154137 82200 6 la_oenb[91]
port 444 nsew signal output
rlabel metal2 s 155765 81600 155793 82200 6 la_oenb[92]
port 445 nsew signal output
rlabel metal2 s 157467 81600 157495 82200 6 la_oenb[93]
port 446 nsew signal output
rlabel metal2 s 159169 81600 159197 82200 6 la_oenb[94]
port 447 nsew signal output
rlabel metal2 s 160825 81600 160853 82200 6 la_oenb[95]
port 448 nsew signal output
rlabel metal2 s 162527 81600 162555 82200 6 la_oenb[96]
port 449 nsew signal output
rlabel metal2 s 164183 81600 164211 82200 6 la_oenb[97]
port 450 nsew signal output
rlabel metal2 s 165885 81600 165913 82200 6 la_oenb[98]
port 451 nsew signal output
rlabel metal2 s 167541 81600 167569 82200 6 la_oenb[99]
port 452 nsew signal output
rlabel metal2 s 16155 81600 16183 82200 6 la_oenb[9]
port 453 nsew signal output
rlabel metal2 s 1435 81600 1463 82200 6 la_output[0]
port 454 nsew signal output
rlabel metal2 s 169657 81600 169685 82200 6 la_output[100]
port 455 nsew signal output
rlabel metal2 s 171359 81600 171387 82200 6 la_output[101]
port 456 nsew signal output
rlabel metal2 s 173015 81600 173043 82200 6 la_output[102]
port 457 nsew signal output
rlabel metal2 s 174717 81600 174745 82200 6 la_output[103]
port 458 nsew signal output
rlabel metal2 s 176373 81600 176401 82200 6 la_output[104]
port 459 nsew signal output
rlabel metal2 s 178075 81600 178103 82200 6 la_output[105]
port 460 nsew signal output
rlabel metal2 s 179777 81600 179805 82200 6 la_output[106]
port 461 nsew signal output
rlabel metal2 s 181433 81600 181461 82200 6 la_output[107]
port 462 nsew signal output
rlabel metal2 s 183135 81600 183163 82200 6 la_output[108]
port 463 nsew signal output
rlabel metal2 s 184791 81600 184819 82200 6 la_output[109]
port 464 nsew signal output
rlabel metal2 s 18271 81600 18299 82200 6 la_output[10]
port 465 nsew signal output
rlabel metal2 s 186493 81600 186521 82200 6 la_output[110]
port 466 nsew signal output
rlabel metal2 s 188149 81600 188177 82200 6 la_output[111]
port 467 nsew signal output
rlabel metal2 s 189851 81600 189879 82200 6 la_output[112]
port 468 nsew signal output
rlabel metal2 s 191553 81600 191581 82200 6 la_output[113]
port 469 nsew signal output
rlabel metal2 s 193209 81600 193237 82200 6 la_output[114]
port 470 nsew signal output
rlabel metal2 s 194911 81600 194939 82200 6 la_output[115]
port 471 nsew signal output
rlabel metal2 s 196567 81600 196595 82200 6 la_output[116]
port 472 nsew signal output
rlabel metal2 s 198269 81600 198297 82200 6 la_output[117]
port 473 nsew signal output
rlabel metal2 s 199925 81600 199953 82200 6 la_output[118]
port 474 nsew signal output
rlabel metal2 s 201627 81600 201655 82200 6 la_output[119]
port 475 nsew signal output
rlabel metal2 s 19927 81600 19955 82200 6 la_output[11]
port 476 nsew signal output
rlabel metal2 s 203329 81600 203357 82200 6 la_output[120]
port 477 nsew signal output
rlabel metal2 s 204985 81600 205013 82200 6 la_output[121]
port 478 nsew signal output
rlabel metal2 s 206687 81600 206715 82200 6 la_output[122]
port 479 nsew signal output
rlabel metal2 s 208343 81600 208371 82200 6 la_output[123]
port 480 nsew signal output
rlabel metal2 s 210045 81600 210073 82200 6 la_output[124]
port 481 nsew signal output
rlabel metal2 s 211701 81600 211729 82200 6 la_output[125]
port 482 nsew signal output
rlabel metal2 s 213403 81600 213431 82200 6 la_output[126]
port 483 nsew signal output
rlabel metal2 s 215105 81600 215133 82200 6 la_output[127]
port 484 nsew signal output
rlabel metal2 s 21629 81600 21657 82200 6 la_output[12]
port 485 nsew signal output
rlabel metal2 s 23285 81600 23313 82200 6 la_output[13]
port 486 nsew signal output
rlabel metal2 s 24987 81600 25015 82200 6 la_output[14]
port 487 nsew signal output
rlabel metal2 s 26689 81600 26717 82200 6 la_output[15]
port 488 nsew signal output
rlabel metal2 s 28345 81600 28373 82200 6 la_output[16]
port 489 nsew signal output
rlabel metal2 s 30047 81600 30075 82200 6 la_output[17]
port 490 nsew signal output
rlabel metal2 s 31703 81600 31731 82200 6 la_output[18]
port 491 nsew signal output
rlabel metal2 s 33405 81600 33433 82200 6 la_output[19]
port 492 nsew signal output
rlabel metal2 s 3137 81600 3165 82200 6 la_output[1]
port 493 nsew signal output
rlabel metal2 s 35061 81600 35089 82200 6 la_output[20]
port 494 nsew signal output
rlabel metal2 s 36763 81600 36791 82200 6 la_output[21]
port 495 nsew signal output
rlabel metal2 s 38465 81600 38493 82200 6 la_output[22]
port 496 nsew signal output
rlabel metal2 s 40121 81600 40149 82200 6 la_output[23]
port 497 nsew signal output
rlabel metal2 s 41823 81600 41851 82200 6 la_output[24]
port 498 nsew signal output
rlabel metal2 s 43479 81600 43507 82200 6 la_output[25]
port 499 nsew signal output
rlabel metal2 s 45181 81600 45209 82200 6 la_output[26]
port 500 nsew signal output
rlabel metal2 s 46837 81600 46865 82200 6 la_output[27]
port 501 nsew signal output
rlabel metal2 s 48539 81600 48567 82200 6 la_output[28]
port 502 nsew signal output
rlabel metal2 s 50241 81600 50269 82200 6 la_output[29]
port 503 nsew signal output
rlabel metal2 s 4793 81600 4821 82200 6 la_output[2]
port 504 nsew signal output
rlabel metal2 s 51897 81600 51925 82200 6 la_output[30]
port 505 nsew signal output
rlabel metal2 s 53599 81600 53627 82200 6 la_output[31]
port 506 nsew signal output
rlabel metal2 s 55255 81600 55283 82200 6 la_output[32]
port 507 nsew signal output
rlabel metal2 s 56957 81600 56985 82200 6 la_output[33]
port 508 nsew signal output
rlabel metal2 s 58613 81600 58641 82200 6 la_output[34]
port 509 nsew signal output
rlabel metal2 s 60315 81600 60343 82200 6 la_output[35]
port 510 nsew signal output
rlabel metal2 s 62017 81600 62045 82200 6 la_output[36]
port 511 nsew signal output
rlabel metal2 s 63673 81600 63701 82200 6 la_output[37]
port 512 nsew signal output
rlabel metal2 s 65375 81600 65403 82200 6 la_output[38]
port 513 nsew signal output
rlabel metal2 s 67031 81600 67059 82200 6 la_output[39]
port 514 nsew signal output
rlabel metal2 s 6495 81600 6523 82200 6 la_output[3]
port 515 nsew signal output
rlabel metal2 s 68733 81600 68761 82200 6 la_output[40]
port 516 nsew signal output
rlabel metal2 s 70389 81600 70417 82200 6 la_output[41]
port 517 nsew signal output
rlabel metal2 s 72091 81600 72119 82200 6 la_output[42]
port 518 nsew signal output
rlabel metal2 s 73793 81600 73821 82200 6 la_output[43]
port 519 nsew signal output
rlabel metal2 s 75449 81600 75477 82200 6 la_output[44]
port 520 nsew signal output
rlabel metal2 s 77151 81600 77179 82200 6 la_output[45]
port 521 nsew signal output
rlabel metal2 s 78807 81600 78835 82200 6 la_output[46]
port 522 nsew signal output
rlabel metal2 s 80509 81600 80537 82200 6 la_output[47]
port 523 nsew signal output
rlabel metal2 s 82165 81600 82193 82200 6 la_output[48]
port 524 nsew signal output
rlabel metal2 s 83867 81600 83895 82200 6 la_output[49]
port 525 nsew signal output
rlabel metal2 s 8151 81600 8179 82200 6 la_output[4]
port 526 nsew signal output
rlabel metal2 s 85569 81600 85597 82200 6 la_output[50]
port 527 nsew signal output
rlabel metal2 s 87225 81600 87253 82200 6 la_output[51]
port 528 nsew signal output
rlabel metal2 s 88927 81600 88955 82200 6 la_output[52]
port 529 nsew signal output
rlabel metal2 s 90583 81600 90611 82200 6 la_output[53]
port 530 nsew signal output
rlabel metal2 s 92285 81600 92313 82200 6 la_output[54]
port 531 nsew signal output
rlabel metal2 s 93941 81600 93969 82200 6 la_output[55]
port 532 nsew signal output
rlabel metal2 s 95643 81600 95671 82200 6 la_output[56]
port 533 nsew signal output
rlabel metal2 s 97345 81600 97373 82200 6 la_output[57]
port 534 nsew signal output
rlabel metal2 s 99001 81600 99029 82200 6 la_output[58]
port 535 nsew signal output
rlabel metal2 s 100703 81600 100731 82200 6 la_output[59]
port 536 nsew signal output
rlabel metal2 s 9853 81600 9881 82200 6 la_output[5]
port 537 nsew signal output
rlabel metal2 s 102359 81600 102387 82200 6 la_output[60]
port 538 nsew signal output
rlabel metal2 s 104061 81600 104089 82200 6 la_output[61]
port 539 nsew signal output
rlabel metal2 s 105717 81600 105745 82200 6 la_output[62]
port 540 nsew signal output
rlabel metal2 s 107419 81600 107447 82200 6 la_output[63]
port 541 nsew signal output
rlabel metal2 s 109121 81600 109149 82200 6 la_output[64]
port 542 nsew signal output
rlabel metal2 s 110777 81600 110805 82200 6 la_output[65]
port 543 nsew signal output
rlabel metal2 s 112479 81600 112507 82200 6 la_output[66]
port 544 nsew signal output
rlabel metal2 s 114135 81600 114163 82200 6 la_output[67]
port 545 nsew signal output
rlabel metal2 s 115837 81600 115865 82200 6 la_output[68]
port 546 nsew signal output
rlabel metal2 s 117493 81600 117521 82200 6 la_output[69]
port 547 nsew signal output
rlabel metal2 s 11509 81600 11537 82200 6 la_output[6]
port 548 nsew signal output
rlabel metal2 s 119195 81600 119223 82200 6 la_output[70]
port 549 nsew signal output
rlabel metal2 s 120897 81600 120925 82200 6 la_output[71]
port 550 nsew signal output
rlabel metal2 s 122553 81600 122581 82200 6 la_output[72]
port 551 nsew signal output
rlabel metal2 s 124255 81600 124283 82200 6 la_output[73]
port 552 nsew signal output
rlabel metal2 s 125911 81600 125939 82200 6 la_output[74]
port 553 nsew signal output
rlabel metal2 s 127613 81600 127641 82200 6 la_output[75]
port 554 nsew signal output
rlabel metal2 s 129269 81600 129297 82200 6 la_output[76]
port 555 nsew signal output
rlabel metal2 s 130971 81600 130999 82200 6 la_output[77]
port 556 nsew signal output
rlabel metal2 s 132673 81600 132701 82200 6 la_output[78]
port 557 nsew signal output
rlabel metal2 s 134329 81600 134357 82200 6 la_output[79]
port 558 nsew signal output
rlabel metal2 s 13211 81600 13239 82200 6 la_output[7]
port 559 nsew signal output
rlabel metal2 s 136031 81600 136059 82200 6 la_output[80]
port 560 nsew signal output
rlabel metal2 s 137687 81600 137715 82200 6 la_output[81]
port 561 nsew signal output
rlabel metal2 s 139389 81600 139417 82200 6 la_output[82]
port 562 nsew signal output
rlabel metal2 s 141045 81600 141073 82200 6 la_output[83]
port 563 nsew signal output
rlabel metal2 s 142747 81600 142775 82200 6 la_output[84]
port 564 nsew signal output
rlabel metal2 s 144449 81600 144477 82200 6 la_output[85]
port 565 nsew signal output
rlabel metal2 s 146105 81600 146133 82200 6 la_output[86]
port 566 nsew signal output
rlabel metal2 s 147807 81600 147835 82200 6 la_output[87]
port 567 nsew signal output
rlabel metal2 s 149463 81600 149491 82200 6 la_output[88]
port 568 nsew signal output
rlabel metal2 s 151165 81600 151193 82200 6 la_output[89]
port 569 nsew signal output
rlabel metal2 s 14913 81600 14941 82200 6 la_output[8]
port 570 nsew signal output
rlabel metal2 s 152821 81600 152849 82200 6 la_output[90]
port 571 nsew signal output
rlabel metal2 s 154523 81600 154551 82200 6 la_output[91]
port 572 nsew signal output
rlabel metal2 s 156225 81600 156253 82200 6 la_output[92]
port 573 nsew signal output
rlabel metal2 s 157881 81600 157909 82200 6 la_output[93]
port 574 nsew signal output
rlabel metal2 s 159583 81600 159611 82200 6 la_output[94]
port 575 nsew signal output
rlabel metal2 s 161239 81600 161267 82200 6 la_output[95]
port 576 nsew signal output
rlabel metal2 s 162941 81600 162969 82200 6 la_output[96]
port 577 nsew signal output
rlabel metal2 s 164597 81600 164625 82200 6 la_output[97]
port 578 nsew signal output
rlabel metal2 s 166299 81600 166327 82200 6 la_output[98]
port 579 nsew signal output
rlabel metal2 s 168001 81600 168029 82200 6 la_output[99]
port 580 nsew signal output
rlabel metal2 s 16569 81600 16597 82200 6 la_output[9]
port 581 nsew signal output
rlabel metal2 s 215519 81600 215547 82200 6 mprj_ack_i
port 582 nsew signal input
rlabel metal2 s 217589 81600 217617 82200 6 mprj_adr_o[0]
port 583 nsew signal output
rlabel metal2 s 231895 81600 231923 82200 6 mprj_adr_o[10]
port 584 nsew signal output
rlabel metal2 s 233183 81600 233211 82200 6 mprj_adr_o[11]
port 585 nsew signal output
rlabel metal2 s 234425 81600 234453 82200 6 mprj_adr_o[12]
port 586 nsew signal output
rlabel metal2 s 235713 81600 235741 82200 6 mprj_adr_o[13]
port 587 nsew signal output
rlabel metal2 s 236955 81600 236983 82200 6 mprj_adr_o[14]
port 588 nsew signal output
rlabel metal2 s 238197 81600 238225 82200 6 mprj_adr_o[15]
port 589 nsew signal output
rlabel metal2 s 239485 81600 239513 82200 6 mprj_adr_o[16]
port 590 nsew signal output
rlabel metal2 s 240727 81600 240755 82200 6 mprj_adr_o[17]
port 591 nsew signal output
rlabel metal2 s 242015 81600 242043 82200 6 mprj_adr_o[18]
port 592 nsew signal output
rlabel metal2 s 243257 81600 243285 82200 6 mprj_adr_o[19]
port 593 nsew signal output
rlabel metal2 s 219291 81600 219319 82200 6 mprj_adr_o[1]
port 594 nsew signal output
rlabel metal2 s 244545 81600 244573 82200 6 mprj_adr_o[20]
port 595 nsew signal output
rlabel metal2 s 245787 81600 245815 82200 6 mprj_adr_o[21]
port 596 nsew signal output
rlabel metal2 s 247029 81600 247057 82200 6 mprj_adr_o[22]
port 597 nsew signal output
rlabel metal2 s 248317 81600 248345 82200 6 mprj_adr_o[23]
port 598 nsew signal output
rlabel metal2 s 249559 81600 249587 82200 6 mprj_adr_o[24]
port 599 nsew signal output
rlabel metal2 s 250847 81600 250875 82200 6 mprj_adr_o[25]
port 600 nsew signal output
rlabel metal2 s 252089 81600 252117 82200 6 mprj_adr_o[26]
port 601 nsew signal output
rlabel metal2 s 253377 81600 253405 82200 6 mprj_adr_o[27]
port 602 nsew signal output
rlabel metal2 s 254619 81600 254647 82200 6 mprj_adr_o[28]
port 603 nsew signal output
rlabel metal2 s 255861 81600 255889 82200 6 mprj_adr_o[29]
port 604 nsew signal output
rlabel metal2 s 220993 81600 221021 82200 6 mprj_adr_o[2]
port 605 nsew signal output
rlabel metal2 s 257149 81600 257177 82200 6 mprj_adr_o[30]
port 606 nsew signal output
rlabel metal2 s 258391 81600 258419 82200 6 mprj_adr_o[31]
port 607 nsew signal output
rlabel metal2 s 222649 81600 222677 82200 6 mprj_adr_o[3]
port 608 nsew signal output
rlabel metal2 s 224351 81600 224379 82200 6 mprj_adr_o[4]
port 609 nsew signal output
rlabel metal2 s 225593 81600 225621 82200 6 mprj_adr_o[5]
port 610 nsew signal output
rlabel metal2 s 226881 81600 226909 82200 6 mprj_adr_o[6]
port 611 nsew signal output
rlabel metal2 s 228123 81600 228151 82200 6 mprj_adr_o[7]
port 612 nsew signal output
rlabel metal2 s 229365 81600 229393 82200 6 mprj_adr_o[8]
port 613 nsew signal output
rlabel metal2 s 230653 81600 230681 82200 6 mprj_adr_o[9]
port 614 nsew signal output
rlabel metal2 s 215933 81600 215961 82200 6 mprj_cyc_o
port 615 nsew signal output
rlabel metal2 s 218049 81600 218077 82200 6 mprj_dat_i[0]
port 616 nsew signal input
rlabel metal2 s 232309 81600 232337 82200 6 mprj_dat_i[10]
port 617 nsew signal input
rlabel metal2 s 233597 81600 233625 82200 6 mprj_dat_i[11]
port 618 nsew signal input
rlabel metal2 s 234839 81600 234867 82200 6 mprj_dat_i[12]
port 619 nsew signal input
rlabel metal2 s 236127 81600 236155 82200 6 mprj_dat_i[13]
port 620 nsew signal input
rlabel metal2 s 237369 81600 237397 82200 6 mprj_dat_i[14]
port 621 nsew signal input
rlabel metal2 s 238657 81600 238685 82200 6 mprj_dat_i[15]
port 622 nsew signal input
rlabel metal2 s 239899 81600 239927 82200 6 mprj_dat_i[16]
port 623 nsew signal input
rlabel metal2 s 241141 81600 241169 82200 6 mprj_dat_i[17]
port 624 nsew signal input
rlabel metal2 s 242429 81600 242457 82200 6 mprj_dat_i[18]
port 625 nsew signal input
rlabel metal2 s 243671 81600 243699 82200 6 mprj_dat_i[19]
port 626 nsew signal input
rlabel metal2 s 219705 81600 219733 82200 6 mprj_dat_i[1]
port 627 nsew signal input
rlabel metal2 s 244959 81600 244987 82200 6 mprj_dat_i[20]
port 628 nsew signal input
rlabel metal2 s 246201 81600 246229 82200 6 mprj_dat_i[21]
port 629 nsew signal input
rlabel metal2 s 247489 81600 247517 82200 6 mprj_dat_i[22]
port 630 nsew signal input
rlabel metal2 s 248731 81600 248759 82200 6 mprj_dat_i[23]
port 631 nsew signal input
rlabel metal2 s 249973 81600 250001 82200 6 mprj_dat_i[24]
port 632 nsew signal input
rlabel metal2 s 251261 81600 251289 82200 6 mprj_dat_i[25]
port 633 nsew signal input
rlabel metal2 s 252503 81600 252531 82200 6 mprj_dat_i[26]
port 634 nsew signal input
rlabel metal2 s 253791 81600 253819 82200 6 mprj_dat_i[27]
port 635 nsew signal input
rlabel metal2 s 255033 81600 255061 82200 6 mprj_dat_i[28]
port 636 nsew signal input
rlabel metal2 s 256321 81600 256349 82200 6 mprj_dat_i[29]
port 637 nsew signal input
rlabel metal2 s 221407 81600 221435 82200 6 mprj_dat_i[2]
port 638 nsew signal input
rlabel metal2 s 257563 81600 257591 82200 6 mprj_dat_i[30]
port 639 nsew signal input
rlabel metal2 s 258805 81600 258833 82200 6 mprj_dat_i[31]
port 640 nsew signal input
rlabel metal2 s 223063 81600 223091 82200 6 mprj_dat_i[3]
port 641 nsew signal input
rlabel metal2 s 224765 81600 224793 82200 6 mprj_dat_i[4]
port 642 nsew signal input
rlabel metal2 s 226007 81600 226035 82200 6 mprj_dat_i[5]
port 643 nsew signal input
rlabel metal2 s 227295 81600 227323 82200 6 mprj_dat_i[6]
port 644 nsew signal input
rlabel metal2 s 228537 81600 228565 82200 6 mprj_dat_i[7]
port 645 nsew signal input
rlabel metal2 s 229825 81600 229853 82200 6 mprj_dat_i[8]
port 646 nsew signal input
rlabel metal2 s 231067 81600 231095 82200 6 mprj_dat_i[9]
port 647 nsew signal input
rlabel metal2 s 218463 81600 218491 82200 6 mprj_dat_o[0]
port 648 nsew signal output
rlabel metal2 s 232769 81600 232797 82200 6 mprj_dat_o[10]
port 649 nsew signal output
rlabel metal2 s 234011 81600 234039 82200 6 mprj_dat_o[11]
port 650 nsew signal output
rlabel metal2 s 235253 81600 235281 82200 6 mprj_dat_o[12]
port 651 nsew signal output
rlabel metal2 s 236541 81600 236569 82200 6 mprj_dat_o[13]
port 652 nsew signal output
rlabel metal2 s 237783 81600 237811 82200 6 mprj_dat_o[14]
port 653 nsew signal output
rlabel metal2 s 239071 81600 239099 82200 6 mprj_dat_o[15]
port 654 nsew signal output
rlabel metal2 s 240313 81600 240341 82200 6 mprj_dat_o[16]
port 655 nsew signal output
rlabel metal2 s 241601 81600 241629 82200 6 mprj_dat_o[17]
port 656 nsew signal output
rlabel metal2 s 242843 81600 242871 82200 6 mprj_dat_o[18]
port 657 nsew signal output
rlabel metal2 s 244085 81600 244113 82200 6 mprj_dat_o[19]
port 658 nsew signal output
rlabel metal2 s 220119 81600 220147 82200 6 mprj_dat_o[1]
port 659 nsew signal output
rlabel metal2 s 245373 81600 245401 82200 6 mprj_dat_o[20]
port 660 nsew signal output
rlabel metal2 s 246615 81600 246643 82200 6 mprj_dat_o[21]
port 661 nsew signal output
rlabel metal2 s 247903 81600 247931 82200 6 mprj_dat_o[22]
port 662 nsew signal output
rlabel metal2 s 249145 81600 249173 82200 6 mprj_dat_o[23]
port 663 nsew signal output
rlabel metal2 s 250433 81600 250461 82200 6 mprj_dat_o[24]
port 664 nsew signal output
rlabel metal2 s 251675 81600 251703 82200 6 mprj_dat_o[25]
port 665 nsew signal output
rlabel metal2 s 252917 81600 252945 82200 6 mprj_dat_o[26]
port 666 nsew signal output
rlabel metal2 s 254205 81600 254233 82200 6 mprj_dat_o[27]
port 667 nsew signal output
rlabel metal2 s 255447 81600 255475 82200 6 mprj_dat_o[28]
port 668 nsew signal output
rlabel metal2 s 256735 81600 256763 82200 6 mprj_dat_o[29]
port 669 nsew signal output
rlabel metal2 s 221821 81600 221849 82200 6 mprj_dat_o[2]
port 670 nsew signal output
rlabel metal2 s 257977 81600 258005 82200 6 mprj_dat_o[30]
port 671 nsew signal output
rlabel metal2 s 259265 81600 259293 82200 6 mprj_dat_o[31]
port 672 nsew signal output
rlabel metal2 s 223477 81600 223505 82200 6 mprj_dat_o[3]
port 673 nsew signal output
rlabel metal2 s 225179 81600 225207 82200 6 mprj_dat_o[4]
port 674 nsew signal output
rlabel metal2 s 226421 81600 226449 82200 6 mprj_dat_o[5]
port 675 nsew signal output
rlabel metal2 s 227709 81600 227737 82200 6 mprj_dat_o[6]
port 676 nsew signal output
rlabel metal2 s 228951 81600 228979 82200 6 mprj_dat_o[7]
port 677 nsew signal output
rlabel metal2 s 230239 81600 230267 82200 6 mprj_dat_o[8]
port 678 nsew signal output
rlabel metal2 s 231481 81600 231509 82200 6 mprj_dat_o[9]
port 679 nsew signal output
rlabel metal2 s 218877 81600 218905 82200 6 mprj_sel_o[0]
port 680 nsew signal output
rlabel metal2 s 220533 81600 220561 82200 6 mprj_sel_o[1]
port 681 nsew signal output
rlabel metal2 s 222235 81600 222263 82200 6 mprj_sel_o[2]
port 682 nsew signal output
rlabel metal2 s 223937 81600 223965 82200 6 mprj_sel_o[3]
port 683 nsew signal output
rlabel metal2 s 216347 81600 216375 82200 6 mprj_stb_o
port 684 nsew signal output
rlabel metal2 s 216761 81600 216789 82200 6 mprj_wb_iena
port 685 nsew signal output
rlabel metal2 s 217175 81600 217203 82200 6 mprj_we_o
port 686 nsew signal output
rlabel metal3 s 261600 44680 262200 44740 6 qspi_enabled
port 687 nsew signal output
rlabel metal3 s 261600 41688 262200 41748 6 ser_rx
port 688 nsew signal input
rlabel metal3 s 261600 42436 262200 42496 6 ser_tx
port 689 nsew signal output
rlabel metal3 s 261600 40192 262200 40252 6 spi_csb
port 690 nsew signal output
rlabel metal3 s 261600 43184 262200 43244 6 spi_enabled
port 691 nsew signal output
rlabel metal3 s 261600 39444 262200 39504 6 spi_sck
port 692 nsew signal output
rlabel metal3 s 261600 40940 262200 41000 6 spi_sdi
port 693 nsew signal input
rlabel metal3 s 261600 38696 262200 38756 6 spi_sdo
port 694 nsew signal output
rlabel metal3 s 261600 37948 262200 38008 6 spi_sdoenb
port 695 nsew signal output
rlabel metal3 s 261600 1092 262200 1152 6 sram_ro_addr[0]
port 696 nsew signal input
rlabel metal3 s 261600 1840 262200 1900 6 sram_ro_addr[1]
port 697 nsew signal input
rlabel metal3 s 261600 2588 262200 2648 6 sram_ro_addr[2]
port 698 nsew signal input
rlabel metal3 s 261600 3336 262200 3396 6 sram_ro_addr[3]
port 699 nsew signal input
rlabel metal3 s 261600 4084 262200 4144 6 sram_ro_addr[4]
port 700 nsew signal input
rlabel metal3 s 261600 4832 262200 4892 6 sram_ro_addr[5]
port 701 nsew signal input
rlabel metal3 s 261600 5580 262200 5640 6 sram_ro_addr[6]
port 702 nsew signal input
rlabel metal3 s 261600 6328 262200 6388 6 sram_ro_addr[7]
port 703 nsew signal input
rlabel metal3 s 261600 7076 262200 7136 6 sram_ro_clk
port 704 nsew signal input
rlabel metal3 s 261600 344 262200 404 6 sram_ro_csb
port 705 nsew signal input
rlabel metal3 s 261600 7824 262200 7884 6 sram_ro_data[0]
port 706 nsew signal output
rlabel metal3 s 261600 15372 262200 15432 6 sram_ro_data[10]
port 707 nsew signal output
rlabel metal3 s 261600 16120 262200 16180 6 sram_ro_data[11]
port 708 nsew signal output
rlabel metal3 s 261600 16868 262200 16928 6 sram_ro_data[12]
port 709 nsew signal output
rlabel metal3 s 261600 17616 262200 17676 6 sram_ro_data[13]
port 710 nsew signal output
rlabel metal3 s 261600 18364 262200 18424 6 sram_ro_data[14]
port 711 nsew signal output
rlabel metal3 s 261600 19112 262200 19172 6 sram_ro_data[15]
port 712 nsew signal output
rlabel metal3 s 261600 19860 262200 19920 6 sram_ro_data[16]
port 713 nsew signal output
rlabel metal3 s 261600 20608 262200 20668 6 sram_ro_data[17]
port 714 nsew signal output
rlabel metal3 s 261600 21356 262200 21416 6 sram_ro_data[18]
port 715 nsew signal output
rlabel metal3 s 261600 22104 262200 22164 6 sram_ro_data[19]
port 716 nsew signal output
rlabel metal3 s 261600 8572 262200 8632 6 sram_ro_data[1]
port 717 nsew signal output
rlabel metal3 s 261600 22852 262200 22912 6 sram_ro_data[20]
port 718 nsew signal output
rlabel metal3 s 261600 23600 262200 23660 6 sram_ro_data[21]
port 719 nsew signal output
rlabel metal3 s 261600 24416 262200 24476 6 sram_ro_data[22]
port 720 nsew signal output
rlabel metal3 s 261600 25164 262200 25224 6 sram_ro_data[23]
port 721 nsew signal output
rlabel metal3 s 261600 25912 262200 25972 6 sram_ro_data[24]
port 722 nsew signal output
rlabel metal3 s 261600 26660 262200 26720 6 sram_ro_data[25]
port 723 nsew signal output
rlabel metal3 s 261600 27408 262200 27468 6 sram_ro_data[26]
port 724 nsew signal output
rlabel metal3 s 261600 28156 262200 28216 6 sram_ro_data[27]
port 725 nsew signal output
rlabel metal3 s 261600 28904 262200 28964 6 sram_ro_data[28]
port 726 nsew signal output
rlabel metal3 s 261600 29652 262200 29712 6 sram_ro_data[29]
port 727 nsew signal output
rlabel metal3 s 261600 9320 262200 9380 6 sram_ro_data[2]
port 728 nsew signal output
rlabel metal3 s 261600 30400 262200 30460 6 sram_ro_data[30]
port 729 nsew signal output
rlabel metal3 s 261600 31148 262200 31208 6 sram_ro_data[31]
port 730 nsew signal output
rlabel metal3 s 261600 10068 262200 10128 6 sram_ro_data[3]
port 731 nsew signal output
rlabel metal3 s 261600 10816 262200 10876 6 sram_ro_data[4]
port 732 nsew signal output
rlabel metal3 s 261600 11564 262200 11624 6 sram_ro_data[5]
port 733 nsew signal output
rlabel metal3 s 261600 12380 262200 12440 6 sram_ro_data[6]
port 734 nsew signal output
rlabel metal3 s 261600 13128 262200 13188 6 sram_ro_data[7]
port 735 nsew signal output
rlabel metal3 s 261600 13876 262200 13936 6 sram_ro_data[8]
port 736 nsew signal output
rlabel metal3 s 261600 14624 262200 14684 6 sram_ro_data[9]
port 737 nsew signal output
rlabel metal3 s 261600 34888 262200 34948 6 trap
port 738 nsew signal output
rlabel metal3 s 261600 43932 262200 43992 6 uart_enabled
port 739 nsew signal output
rlabel metal2 s 259679 81600 259707 82200 6 user_irq_ena[0]
port 740 nsew signal output
rlabel metal2 s 260093 81600 260121 82200 6 user_irq_ena[1]
port 741 nsew signal output
rlabel metal2 s 260507 81600 260535 82200 6 user_irq_ena[2]
port 742 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 262000 82000
string LEFview TRUE
<< end >>
