module caravel_logo ();
endmodule
