magic
tech sky130A
magscale 1 2
timestamp 1650313688
<< checkpaint >>
rect -378 4132 11142 12732
rect -102 372 11142 4132
rect 1738 -220 11142 372
<< isosubstrate >>
rect 1090 1552 2656 4518
<< viali >>
rect 1685 11305 1719 11339
rect 3893 11305 3927 11339
rect 4077 11305 4111 11339
rect 6193 11305 6227 11339
rect 6377 11305 6411 11339
rect 7205 11305 7239 11339
rect 7389 11305 7423 11339
rect 9321 11305 9355 11339
rect 1777 11237 1811 11271
rect 4445 11237 4479 11271
rect 5733 11237 5767 11271
rect 5917 11237 5951 11271
rect 7941 11237 7975 11271
rect 8309 11237 8343 11271
rect 2973 11169 3007 11203
rect 2145 11101 2179 11135
rect 2237 11101 2271 11135
rect 2881 11101 2915 11135
rect 3157 11101 3191 11135
rect 4261 11101 4295 11135
rect 4905 11101 4939 11135
rect 5641 11101 5675 11135
rect 7481 11101 7515 11135
rect 7757 11101 7791 11135
rect 8033 11101 8067 11135
rect 8493 11101 8527 11135
rect 9137 11101 9171 11135
rect 2513 11033 2547 11067
rect 2697 11033 2731 11067
rect 4537 11033 4571 11067
rect 4721 11033 4755 11067
rect 4997 11033 5031 11067
rect 5181 11033 5215 11067
rect 5365 11033 5399 11067
rect 6561 11033 6595 11067
rect 7021 11033 7055 11067
rect 7573 11033 7607 11067
rect 8861 11033 8895 11067
rect 9045 11033 9079 11067
rect 9413 11033 9447 11067
rect 2053 10965 2087 10999
rect 2421 10965 2455 10999
rect 3341 10965 3375 10999
rect 3617 10965 3651 10999
rect 5457 10965 5491 10999
rect 8217 10965 8251 10999
rect 1409 10761 1443 10795
rect 5181 10761 5215 10795
rect 8217 10761 8251 10795
rect 8585 10761 8619 10795
rect 1593 10625 1627 10659
rect 1869 10625 1903 10659
rect 3709 10625 3743 10659
rect 4445 10625 4479 10659
rect 5457 10625 5491 10659
rect 6193 10625 6227 10659
rect 6929 10625 6963 10659
rect 7205 10625 7239 10659
rect 7481 10625 7515 10659
rect 7757 10625 7791 10659
rect 8033 10625 8067 10659
rect 8401 10625 8435 10659
rect 2237 10557 2271 10591
rect 4905 10557 4939 10591
rect 5917 10557 5951 10591
rect 8769 10557 8803 10591
rect 9505 10557 9539 10591
rect 1777 10489 1811 10523
rect 7573 10489 7607 10523
rect 9137 10489 9171 10523
rect 4273 10421 4307 10455
rect 4721 10421 4755 10455
rect 5733 10421 5767 10455
rect 6285 10421 6319 10455
rect 6653 10421 6687 10455
rect 7021 10421 7055 10455
rect 7389 10421 7423 10455
rect 7941 10421 7975 10455
rect 9229 10421 9263 10455
rect 2881 10217 2915 10251
rect 3249 10217 3283 10251
rect 3893 10217 3927 10251
rect 4721 10217 4755 10251
rect 1317 10013 1351 10047
rect 1961 10013 1995 10047
rect 2053 10013 2087 10047
rect 3341 10013 3375 10047
rect 3617 10013 3651 10047
rect 6101 10013 6135 10047
rect 6469 10013 6503 10047
rect 7941 10013 7975 10047
rect 9413 10013 9447 10047
rect 6009 9945 6043 9979
rect 8505 9945 8539 9979
rect 2697 9877 2731 9911
rect 4077 9877 4111 9911
rect 8769 9877 8803 9911
rect 1317 9673 1351 9707
rect 6745 9673 6779 9707
rect 2789 9605 2823 9639
rect 6193 9605 6227 9639
rect 6561 9605 6595 9639
rect 3249 9537 3283 9571
rect 5365 9537 5399 9571
rect 6377 9537 6411 9571
rect 6837 9537 6871 9571
rect 6929 9537 6963 9571
rect 8769 9537 8803 9571
rect 3065 9469 3099 9503
rect 3525 9469 3559 9503
rect 3893 9469 3927 9503
rect 7297 9469 7331 9503
rect 3433 9333 3467 9367
rect 5929 9333 5963 9367
rect 9333 9333 9367 9367
rect 3065 9129 3099 9163
rect 3985 9129 4019 9163
rect 4169 9129 4203 9163
rect 4537 9129 4571 9163
rect 5733 9129 5767 9163
rect 5181 9061 5215 9095
rect 8493 9061 8527 9095
rect 6193 8993 6227 9027
rect 1317 8925 1351 8959
rect 1961 8925 1995 8959
rect 2053 8925 2087 8959
rect 3433 8925 3467 8959
rect 3801 8925 3835 8959
rect 3893 8925 3927 8959
rect 4353 8925 4387 8959
rect 4629 8925 4663 8959
rect 5089 8925 5123 8959
rect 5549 8925 5583 8959
rect 8309 8925 8343 8959
rect 9321 8925 9355 8959
rect 2789 8857 2823 8891
rect 2973 8857 3007 8891
rect 5365 8857 5399 8891
rect 6009 8857 6043 8891
rect 6469 8857 6503 8891
rect 8125 8857 8159 8891
rect 2697 8789 2731 8823
rect 3341 8789 3375 8823
rect 3617 8789 3651 8823
rect 4905 8789 4939 8823
rect 5917 8789 5951 8823
rect 7941 8789 7975 8823
rect 8769 8789 8803 8823
rect 1777 8585 1811 8619
rect 6285 8585 6319 8619
rect 6837 8585 6871 8619
rect 7205 8585 7239 8619
rect 9137 8585 9171 8619
rect 4721 8517 4755 8551
rect 4905 8517 4939 8551
rect 5365 8517 5399 8551
rect 1869 8449 1903 8483
rect 3709 8449 3743 8483
rect 4445 8449 4479 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 6377 8449 6411 8483
rect 7021 8449 7055 8483
rect 7378 8449 7412 8483
rect 9321 8449 9355 8483
rect 1593 8381 1627 8415
rect 2237 8381 2271 8415
rect 5181 8381 5215 8415
rect 7665 8381 7699 8415
rect 4273 8313 4307 8347
rect 5089 8313 5123 8347
rect 6009 8313 6043 8347
rect 9505 8313 9539 8347
rect 1409 8245 1443 8279
rect 4629 8245 4663 8279
rect 6469 8245 6503 8279
rect 5181 8041 5215 8075
rect 5733 8041 5767 8075
rect 9413 8041 9447 8075
rect 8125 7973 8159 8007
rect 1593 7905 1627 7939
rect 1869 7905 1903 7939
rect 3341 7905 3375 7939
rect 3617 7905 3651 7939
rect 1501 7837 1535 7871
rect 4261 7837 4295 7871
rect 4353 7837 4387 7871
rect 5089 7837 5123 7871
rect 5917 7837 5951 7871
rect 6653 7837 6687 7871
rect 8033 7837 8067 7871
rect 8493 7837 8527 7871
rect 8769 7837 8803 7871
rect 6193 7769 6227 7803
rect 6561 7769 6595 7803
rect 7389 7769 7423 7803
rect 8309 7769 8343 7803
rect 1409 7701 1443 7735
rect 4997 7701 5031 7735
rect 5549 7701 5583 7735
rect 6101 7701 6135 7735
rect 6285 7701 6319 7735
rect 6377 7701 6411 7735
rect 7297 7701 7331 7735
rect 1317 7497 1351 7531
rect 9137 7497 9171 7531
rect 9413 7497 9447 7531
rect 2789 7429 2823 7463
rect 3249 7361 3283 7395
rect 3525 7361 3559 7395
rect 3893 7361 3927 7395
rect 5365 7361 5399 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6929 7361 6963 7395
rect 8401 7361 8435 7395
rect 9321 7361 9355 7395
rect 3065 7293 3099 7327
rect 5929 7225 5963 7259
rect 3341 7157 3375 7191
rect 6193 7157 6227 7191
rect 8585 7157 8619 7191
rect 8961 7157 8995 7191
rect 1764 6953 1798 6987
rect 7401 6953 7435 6987
rect 8861 6953 8895 6987
rect 9413 6953 9447 6987
rect 1501 6817 1535 6851
rect 3249 6817 3283 6851
rect 3617 6817 3651 6851
rect 4353 6817 4387 6851
rect 5917 6817 5951 6851
rect 7665 6817 7699 6851
rect 8217 6817 8251 6851
rect 4261 6749 4295 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 7849 6749 7883 6783
rect 8033 6749 8067 6783
rect 8309 6749 8343 6783
rect 8585 6749 8619 6783
rect 8769 6749 8803 6783
rect 1409 6613 1443 6647
rect 5733 6613 5767 6647
rect 9229 6613 9263 6647
rect 1409 6409 1443 6443
rect 1501 6409 1535 6443
rect 5917 6409 5951 6443
rect 7941 6341 7975 6375
rect 8217 6341 8251 6375
rect 8585 6341 8619 6375
rect 2789 6273 2823 6307
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 5181 6273 5215 6307
rect 8033 6273 8067 6307
rect 8493 6273 8527 6307
rect 8769 6273 8803 6307
rect 8953 6273 8987 6307
rect 9321 6273 9355 6307
rect 1685 6205 1719 6239
rect 2697 6205 2731 6239
rect 3709 6205 3743 6239
rect 6193 6205 6227 6239
rect 9413 6205 9447 6239
rect 2329 6137 2363 6171
rect 2973 6137 3007 6171
rect 5745 6137 5779 6171
rect 2421 6069 2455 6103
rect 3249 6069 3283 6103
rect 8309 6069 8343 6103
rect 1501 5865 1535 5899
rect 1685 5865 1719 5899
rect 3893 5865 3927 5899
rect 4261 5865 4295 5899
rect 8125 5865 8159 5899
rect 8861 5865 8895 5899
rect 3709 5797 3743 5831
rect 5917 5797 5951 5831
rect 9229 5797 9263 5831
rect 9505 5797 9539 5831
rect 1317 5729 1351 5763
rect 6193 5729 6227 5763
rect 3433 5661 3467 5695
rect 4353 5661 4387 5695
rect 4445 5661 4479 5695
rect 5641 5661 5675 5695
rect 8033 5661 8067 5695
rect 9045 5661 9079 5695
rect 9321 5661 9355 5695
rect 3157 5593 3191 5627
rect 7941 5593 7975 5627
rect 8493 5525 8527 5559
rect 6469 5321 6503 5355
rect 7481 5321 7515 5355
rect 5181 5253 5215 5287
rect 7205 5253 7239 5287
rect 8953 5253 8987 5287
rect 3341 5185 3375 5219
rect 4353 5185 4387 5219
rect 5089 5185 5123 5219
rect 7021 5185 7055 5219
rect 8125 5185 8159 5219
rect 8309 5185 8343 5219
rect 9137 5185 9171 5219
rect 9321 5185 9355 5219
rect 4169 5049 4203 5083
rect 7389 5049 7423 5083
rect 3985 4981 4019 5015
rect 4629 4981 4663 5015
rect 4813 4981 4847 5015
rect 8401 4981 8435 5015
rect 8769 4981 8803 5015
rect 9505 4981 9539 5015
rect 3341 4777 3375 4811
rect 3801 4777 3835 4811
rect 4445 4777 4479 4811
rect 6193 4777 6227 4811
rect 8873 4777 8907 4811
rect 9045 4709 9079 4743
rect 4813 4641 4847 4675
rect 6837 4641 6871 4675
rect 3525 4573 3559 4607
rect 3709 4573 3743 4607
rect 4353 4573 4387 4607
rect 5365 4573 5399 4607
rect 5549 4573 5583 4607
rect 6377 4573 6411 4607
rect 6469 4573 6503 4607
rect 8309 4573 8343 4607
rect 9229 4573 9263 4607
rect 9505 4573 9539 4607
rect 4997 4505 5031 4539
rect 5181 4505 5215 4539
rect 5733 4505 5767 4539
rect 5917 4505 5951 4539
rect 6101 4505 6135 4539
rect 4169 4437 4203 4471
rect 9321 4437 9355 4471
rect 3709 4233 3743 4267
rect 9137 4233 9171 4267
rect 6929 4165 6963 4199
rect 3617 4097 3651 4131
rect 3985 4097 4019 4131
rect 6101 4097 6135 4131
rect 7205 4097 7239 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 9229 4097 9263 4131
rect 9505 4097 9539 4131
rect 3525 4029 3559 4063
rect 4261 4029 4295 4063
rect 4629 4029 4663 4063
rect 7297 4029 7331 4063
rect 8861 4029 8895 4063
rect 7113 3961 7147 3995
rect 4169 3893 4203 3927
rect 6665 3893 6699 3927
rect 7481 3893 7515 3927
rect 9321 3893 9355 3927
rect 3341 3689 3375 3723
rect 3617 3689 3651 3723
rect 4445 3689 4479 3723
rect 6469 3689 6503 3723
rect 9149 3689 9183 3723
rect 4813 3621 4847 3655
rect 5733 3621 5767 3655
rect 5457 3553 5491 3587
rect 6745 3553 6779 3587
rect 7113 3553 7147 3587
rect 3893 3485 3927 3519
rect 3985 3485 4019 3519
rect 4261 3485 4295 3519
rect 4537 3485 4571 3519
rect 5549 3485 5583 3519
rect 6377 3485 6411 3519
rect 6653 3485 6687 3519
rect 8585 3485 8619 3519
rect 9505 3485 9539 3519
rect 4997 3417 5031 3451
rect 3801 3349 3835 3383
rect 4169 3349 4203 3383
rect 4721 3349 4755 3383
rect 5273 3349 5307 3383
rect 9321 3349 9355 3383
rect 3525 3145 3559 3179
rect 8309 3145 8343 3179
rect 6561 3077 6595 3111
rect 8861 3077 8895 3111
rect 3617 3009 3651 3043
rect 5457 3009 5491 3043
rect 8493 3009 8527 3043
rect 3985 2941 4019 2975
rect 6285 2941 6319 2975
rect 8033 2941 8067 2975
rect 8769 2941 8803 2975
rect 9413 2941 9447 2975
rect 6021 2805 6055 2839
rect 5365 2601 5399 2635
rect 8133 2601 8167 2635
rect 9137 2601 9171 2635
rect 5089 2533 5123 2567
rect 3341 2465 3375 2499
rect 5733 2465 5767 2499
rect 8309 2465 8343 2499
rect 5549 2397 5583 2431
rect 6101 2397 6135 2431
rect 7573 2397 7607 2431
rect 8861 2397 8895 2431
rect 9229 2397 9263 2431
rect 9505 2397 9539 2431
rect 3617 2329 3651 2363
rect 9321 2261 9355 2295
rect 4077 2057 4111 2091
rect 7941 2057 7975 2091
rect 4537 1989 4571 2023
rect 4261 1921 4295 1955
rect 6193 1921 6227 1955
rect 8309 1921 8343 1955
rect 6469 1853 6503 1887
rect 8861 1853 8895 1887
rect 8953 1853 8987 1887
rect 6009 1717 6043 1751
rect 9505 1717 9539 1751
rect 5733 1513 5767 1547
rect 5917 1513 5951 1547
rect 6745 1513 6779 1547
rect 7757 1513 7791 1547
rect 9321 1513 9355 1547
rect 7849 1445 7883 1479
rect 8309 1445 8343 1479
rect 8493 1445 8527 1479
rect 3341 1377 3375 1411
rect 3617 1377 3651 1411
rect 9229 1377 9263 1411
rect 5365 1309 5399 1343
rect 5457 1309 5491 1343
rect 6101 1309 6135 1343
rect 7481 1309 7515 1343
rect 7573 1309 7607 1343
rect 8861 1309 8895 1343
rect 9045 1309 9079 1343
rect 8125 1241 8159 1275
rect 5089 1173 5123 1207
rect 6837 1173 6871 1207
<< metal1 >>
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 1670 11336 1676 11348
rect 1583 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11336 1734 11348
rect 2130 11336 2136 11348
rect 1728 11308 2136 11336
rect 1728 11296 1734 11308
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 3881 11339 3939 11345
rect 3881 11336 3893 11339
rect 2464 11308 3893 11336
rect 2464 11296 2470 11308
rect 3881 11305 3893 11308
rect 3927 11336 3939 11339
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 3927 11308 4077 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11237 1823 11271
rect 1765 11231 1823 11237
rect 1780 11200 1808 11231
rect 1854 11228 1860 11280
rect 1912 11268 1918 11280
rect 3602 11268 3608 11280
rect 1912 11240 3608 11268
rect 1912 11228 1918 11240
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 2406 11200 2412 11212
rect 1780 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2516 11172 2973 11200
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1820 11104 2145 11132
rect 1820 11092 1826 11104
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2280 11104 2325 11132
rect 2280 11092 2286 11104
rect 1394 11024 1400 11076
rect 1452 11064 1458 11076
rect 2314 11064 2320 11076
rect 1452 11036 2320 11064
rect 1452 11024 1458 11036
rect 2314 11024 2320 11036
rect 2372 11064 2378 11076
rect 2516 11073 2544 11172
rect 2961 11169 2973 11172
rect 3007 11169 3019 11203
rect 2961 11163 3019 11169
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 3145 11135 3203 11141
rect 3145 11132 3157 11135
rect 2915 11104 3157 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 3145 11101 3157 11104
rect 3191 11101 3203 11135
rect 3145 11095 3203 11101
rect 2501 11067 2559 11073
rect 2501 11064 2513 11067
rect 2372 11036 2513 11064
rect 2372 11024 2378 11036
rect 2501 11033 2513 11036
rect 2547 11033 2559 11067
rect 2501 11027 2559 11033
rect 2685 11067 2743 11073
rect 2685 11033 2697 11067
rect 2731 11064 2743 11067
rect 4080 11064 4108 11299
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 6178 11336 6184 11348
rect 4672 11308 6184 11336
rect 4672 11296 4678 11308
rect 6178 11296 6184 11308
rect 6236 11336 6242 11348
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 6236 11308 6377 11336
rect 6236 11296 6242 11308
rect 6365 11305 6377 11308
rect 6411 11305 6423 11339
rect 6365 11299 6423 11305
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 7239 11308 7389 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7377 11305 7389 11308
rect 7423 11336 7435 11339
rect 9309 11339 9367 11345
rect 7423 11308 8892 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 4430 11268 4436 11280
rect 4391 11240 4436 11268
rect 4430 11228 4436 11240
rect 4488 11228 4494 11280
rect 5074 11228 5080 11280
rect 5132 11268 5138 11280
rect 5721 11271 5779 11277
rect 5721 11268 5733 11271
rect 5132 11240 5733 11268
rect 5132 11228 5138 11240
rect 5721 11237 5733 11240
rect 5767 11268 5779 11271
rect 5905 11271 5963 11277
rect 5905 11268 5917 11271
rect 5767 11240 5917 11268
rect 5767 11237 5779 11240
rect 5721 11231 5779 11237
rect 5905 11237 5917 11240
rect 5951 11237 5963 11271
rect 5905 11231 5963 11237
rect 6914 11228 6920 11280
rect 6972 11268 6978 11280
rect 7929 11271 7987 11277
rect 6972 11240 7788 11268
rect 6972 11228 6978 11240
rect 4522 11160 4528 11212
rect 4580 11200 4586 11212
rect 4580 11172 7512 11200
rect 4580 11160 4586 11172
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 7484 11141 7512 11172
rect 7760 11141 7788 11240
rect 7929 11237 7941 11271
rect 7975 11268 7987 11271
rect 8018 11268 8024 11280
rect 7975 11240 8024 11268
rect 7975 11237 7987 11240
rect 7929 11231 7987 11237
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 8297 11271 8355 11277
rect 8297 11237 8309 11271
rect 8343 11268 8355 11271
rect 8386 11268 8392 11280
rect 8343 11240 8392 11268
rect 8343 11237 8355 11240
rect 8297 11231 8355 11237
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11132 4951 11135
rect 5629 11135 5687 11141
rect 5629 11132 5641 11135
rect 4939 11104 5641 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 5629 11101 5641 11104
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 8110 11132 8116 11144
rect 8067 11104 8116 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 4338 11064 4344 11076
rect 2731 11036 3188 11064
rect 4080 11036 4344 11064
rect 2731 11033 2743 11036
rect 2685 11027 2743 11033
rect 3160 11008 3188 11036
rect 4338 11024 4344 11036
rect 4396 11064 4402 11076
rect 4525 11067 4583 11073
rect 4525 11064 4537 11067
rect 4396 11036 4537 11064
rect 4396 11024 4402 11036
rect 4525 11033 4537 11036
rect 4571 11033 4583 11067
rect 4525 11027 4583 11033
rect 4709 11067 4767 11073
rect 4709 11033 4721 11067
rect 4755 11064 4767 11067
rect 4985 11067 5043 11073
rect 4755 11036 4936 11064
rect 4755 11033 4767 11036
rect 4709 11027 4767 11033
rect 4908 11008 4936 11036
rect 4985 11033 4997 11067
rect 5031 11064 5043 11067
rect 5074 11064 5080 11076
rect 5031 11036 5080 11064
rect 5031 11033 5043 11036
rect 4985 11027 5043 11033
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 5169 11067 5227 11073
rect 5169 11033 5181 11067
rect 5215 11033 5227 11067
rect 5169 11027 5227 11033
rect 5353 11067 5411 11073
rect 5353 11033 5365 11067
rect 5399 11064 5411 11067
rect 5399 11036 5580 11064
rect 5399 11033 5411 11036
rect 5353 11027 5411 11033
rect 2038 10996 2044 11008
rect 1999 10968 2044 10996
rect 2038 10956 2044 10968
rect 2096 10956 2102 11008
rect 2409 10999 2467 11005
rect 2409 10965 2421 10999
rect 2455 10996 2467 10999
rect 2590 10996 2596 11008
rect 2455 10968 2596 10996
rect 2455 10965 2467 10968
rect 2409 10959 2467 10965
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 3142 10956 3148 11008
rect 3200 10956 3206 11008
rect 3329 10999 3387 11005
rect 3329 10965 3341 10999
rect 3375 10996 3387 10999
rect 3510 10996 3516 11008
rect 3375 10968 3516 10996
rect 3375 10965 3387 10968
rect 3329 10959 3387 10965
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 3602 10956 3608 11008
rect 3660 10996 3666 11008
rect 4890 10996 4896 11008
rect 3660 10968 3705 10996
rect 4803 10968 4896 10996
rect 3660 10956 3666 10968
rect 4890 10956 4896 10968
rect 4948 10996 4954 11008
rect 5184 10996 5212 11027
rect 5442 10996 5448 11008
rect 4948 10968 5212 10996
rect 5403 10968 5448 10996
rect 4948 10956 4954 10968
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 5552 10996 5580 11036
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 6270 11064 6276 11076
rect 5776 11036 6276 11064
rect 5776 11024 5782 11036
rect 6270 11024 6276 11036
rect 6328 11064 6334 11076
rect 6549 11067 6607 11073
rect 6549 11064 6561 11067
rect 6328 11036 6561 11064
rect 6328 11024 6334 11036
rect 6549 11033 6561 11036
rect 6595 11033 6607 11067
rect 7006 11064 7012 11076
rect 6967 11036 7012 11064
rect 6549 11027 6607 11033
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 7190 11024 7196 11076
rect 7248 11064 7254 11076
rect 7561 11067 7619 11073
rect 7561 11064 7573 11067
rect 7248 11036 7573 11064
rect 7248 11024 7254 11036
rect 7561 11033 7573 11036
rect 7607 11033 7619 11067
rect 8496 11064 8524 11095
rect 8864 11076 8892 11308
rect 9309 11305 9321 11339
rect 9355 11336 9367 11339
rect 13814 11336 13820 11348
rect 9355 11308 13820 11336
rect 9355 11305 9367 11308
rect 9309 11299 9367 11305
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9324 11132 9352 11299
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 9171 11104 9352 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 8846 11064 8852 11076
rect 7561 11027 7619 11033
rect 7668 11036 8524 11064
rect 8807 11036 8852 11064
rect 6086 10996 6092 11008
rect 5552 10968 6092 10996
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 7374 10956 7380 11008
rect 7432 10996 7438 11008
rect 7668 10996 7696 11036
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 9030 11064 9036 11076
rect 8991 11036 9036 11064
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 9401 11067 9459 11073
rect 9401 11064 9413 11067
rect 9140 11036 9413 11064
rect 8202 10996 8208 11008
rect 7432 10968 7696 10996
rect 8163 10968 8208 10996
rect 7432 10956 7438 10968
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 8864 10996 8892 11024
rect 9140 10996 9168 11036
rect 9401 11033 9413 11036
rect 9447 11033 9459 11067
rect 9401 11027 9459 11033
rect 8864 10968 9168 10996
rect 920 10906 9844 10928
rect 920 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 5194 10906
rect 5246 10854 5258 10906
rect 5310 10854 5322 10906
rect 5374 10854 9844 10906
rect 920 10832 9844 10854
rect 1394 10792 1400 10804
rect 1355 10764 1400 10792
rect 1394 10752 1400 10764
rect 1452 10752 1458 10804
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 2188 10764 5181 10792
rect 2188 10752 2194 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 6086 10752 6092 10804
rect 6144 10792 6150 10804
rect 8205 10795 8263 10801
rect 6144 10764 7788 10792
rect 6144 10752 6150 10764
rect 2590 10684 2596 10736
rect 2648 10684 2654 10736
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 5592 10696 7604 10724
rect 5592 10684 5598 10696
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 2038 10656 2044 10668
rect 1903 10628 2044 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3568 10628 3709 10656
rect 3568 10616 3574 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4396 10628 4445 10656
rect 4396 10616 4402 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5040 10628 5457 10656
rect 5040 10616 5046 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 6178 10656 6184 10668
rect 6139 10628 6184 10656
rect 5445 10619 5503 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6362 10616 6368 10668
rect 6420 10656 6426 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6420 10628 6929 10656
rect 6420 10616 6426 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 7156 10628 7205 10656
rect 7156 10616 7162 10628
rect 7193 10625 7205 10628
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 2130 10548 2136 10600
rect 2188 10588 2194 10600
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 2188 10560 2237 10588
rect 2188 10548 2194 10560
rect 2225 10557 2237 10560
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4893 10591 4951 10597
rect 4893 10588 4905 10591
rect 4304 10560 4905 10588
rect 4304 10548 4310 10560
rect 4893 10557 4905 10560
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10588 5963 10591
rect 6822 10588 6828 10600
rect 5951 10560 6828 10588
rect 5951 10557 5963 10560
rect 5905 10551 5963 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7484 10588 7512 10619
rect 7064 10560 7512 10588
rect 7576 10588 7604 10696
rect 7760 10665 7788 10764
rect 8205 10761 8217 10795
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 8573 10795 8631 10801
rect 8573 10761 8585 10795
rect 8619 10792 8631 10795
rect 13906 10792 13912 10804
rect 8619 10764 13912 10792
rect 8619 10761 8631 10764
rect 8573 10755 8631 10761
rect 8220 10724 8248 10755
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 13814 10724 13820 10736
rect 8220 10696 13820 10724
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8036 10588 8064 10619
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 8260 10628 8401 10656
rect 8260 10616 8266 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8754 10588 8760 10600
rect 7576 10560 8064 10588
rect 8715 10560 8760 10588
rect 7064 10548 7070 10560
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 9140 10560 9505 10588
rect 1762 10520 1768 10532
rect 1723 10492 1768 10520
rect 1762 10480 1768 10492
rect 1820 10480 1826 10532
rect 5626 10520 5632 10532
rect 4540 10492 5632 10520
rect 4261 10455 4319 10461
rect 4261 10421 4273 10455
rect 4307 10452 4319 10455
rect 4540 10452 4568 10492
rect 5626 10480 5632 10492
rect 5684 10520 5690 10532
rect 6730 10520 6736 10532
rect 5684 10492 6736 10520
rect 5684 10480 5690 10492
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 9140 10529 9168 10560
rect 9493 10557 9505 10560
rect 9539 10588 9551 10591
rect 13722 10588 13728 10600
rect 9539 10560 13728 10588
rect 9539 10557 9551 10560
rect 9493 10551 9551 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 7561 10523 7619 10529
rect 7561 10520 7573 10523
rect 6972 10492 7573 10520
rect 6972 10480 6978 10492
rect 7561 10489 7573 10492
rect 7607 10489 7619 10523
rect 9125 10523 9183 10529
rect 7561 10483 7619 10489
rect 7668 10492 8616 10520
rect 4307 10424 4568 10452
rect 4307 10421 4319 10424
rect 4261 10415 4319 10421
rect 4614 10412 4620 10464
rect 4672 10452 4678 10464
rect 4709 10455 4767 10461
rect 4709 10452 4721 10455
rect 4672 10424 4721 10452
rect 4672 10412 4678 10424
rect 4709 10421 4721 10424
rect 4755 10452 4767 10455
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 4755 10424 5733 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 5721 10421 5733 10424
rect 5767 10452 5779 10455
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 5767 10424 6285 10452
rect 5767 10421 5779 10424
rect 5721 10415 5779 10421
rect 6273 10421 6285 10424
rect 6319 10421 6331 10455
rect 6638 10452 6644 10464
rect 6599 10424 6644 10452
rect 6273 10415 6331 10421
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7006 10452 7012 10464
rect 6967 10424 7012 10452
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7374 10452 7380 10464
rect 7335 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 7668 10452 7696 10492
rect 7524 10424 7696 10452
rect 7929 10455 7987 10461
rect 7524 10412 7530 10424
rect 7929 10421 7941 10455
rect 7975 10452 7987 10455
rect 8478 10452 8484 10464
rect 7975 10424 8484 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 8588 10452 8616 10492
rect 9125 10489 9137 10523
rect 9171 10489 9183 10523
rect 9125 10483 9183 10489
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 8588 10424 9229 10452
rect 9217 10421 9229 10424
rect 9263 10421 9275 10455
rect 9217 10415 9275 10421
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2869 10251 2927 10257
rect 2869 10248 2881 10251
rect 2280 10220 2881 10248
rect 2280 10208 2286 10220
rect 2869 10217 2881 10220
rect 2915 10217 2927 10251
rect 2869 10211 2927 10217
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3881 10251 3939 10257
rect 3881 10248 3893 10251
rect 3283 10220 3893 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 3881 10217 3893 10220
rect 3927 10248 3939 10251
rect 4154 10248 4160 10260
rect 3927 10220 4160 10248
rect 3927 10217 3939 10220
rect 3881 10211 3939 10217
rect 4154 10208 4160 10220
rect 4212 10248 4218 10260
rect 4614 10248 4620 10260
rect 4212 10220 4620 10248
rect 4212 10208 4218 10220
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 4709 10251 4767 10257
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 6362 10248 6368 10260
rect 4755 10220 6368 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 4724 10112 4752 10211
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 8754 10248 8760 10260
rect 6788 10220 8760 10248
rect 6788 10208 6794 10220
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 1636 10084 4752 10112
rect 1636 10072 1642 10084
rect 1302 10044 1308 10056
rect 1263 10016 1308 10044
rect 1302 10004 1308 10016
rect 1360 10004 1366 10056
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2041 10047 2099 10053
rect 2041 10044 2053 10047
rect 1995 10016 2053 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 2041 10013 2053 10016
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 2314 10004 2320 10056
rect 2372 10044 2378 10056
rect 3329 10047 3387 10053
rect 3329 10044 3341 10047
rect 2372 10016 3341 10044
rect 2372 10004 2378 10016
rect 3329 10013 3341 10016
rect 3375 10013 3387 10047
rect 3602 10044 3608 10056
rect 3563 10016 3608 10044
rect 3329 10007 3387 10013
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 6086 10044 6092 10056
rect 6047 10016 6092 10044
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10044 6515 10047
rect 6546 10044 6552 10056
rect 6503 10016 6552 10044
rect 6503 10013 6515 10016
rect 6457 10007 6515 10013
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 7374 10004 7380 10056
rect 7432 10044 7438 10056
rect 7929 10047 7987 10053
rect 7929 10044 7941 10047
rect 7432 10016 7941 10044
rect 7432 10004 7438 10016
rect 7929 10013 7941 10016
rect 7975 10013 7987 10047
rect 9398 10044 9404 10056
rect 9359 10016 9404 10044
rect 7929 10007 7987 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3620 9976 3648 10004
rect 5994 9976 6000 9988
rect 3016 9948 3648 9976
rect 5955 9948 6000 9976
rect 3016 9936 3022 9948
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 7466 9936 7472 9988
rect 7524 9936 7530 9988
rect 8493 9979 8551 9985
rect 8493 9945 8505 9979
rect 8539 9976 8551 9979
rect 13538 9976 13544 9988
rect 8539 9948 13544 9976
rect 8539 9945 8551 9948
rect 8493 9939 8551 9945
rect 13538 9936 13544 9948
rect 13596 9936 13602 9988
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 2130 9908 2136 9920
rect 1912 9880 2136 9908
rect 1912 9868 1918 9880
rect 2130 9868 2136 9880
rect 2188 9908 2194 9920
rect 2685 9911 2743 9917
rect 2685 9908 2697 9911
rect 2188 9880 2697 9908
rect 2188 9868 2194 9880
rect 2685 9877 2697 9880
rect 2731 9877 2743 9911
rect 2685 9871 2743 9877
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3844 9880 4077 9908
rect 3844 9868 3850 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 7892 9880 8769 9908
rect 7892 9868 7898 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 920 9818 9844 9840
rect 920 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 5194 9818
rect 5246 9766 5258 9818
rect 5310 9766 5322 9818
rect 5374 9766 9844 9818
rect 920 9744 9844 9766
rect 1302 9704 1308 9716
rect 1263 9676 1308 9704
rect 1302 9664 1308 9676
rect 1360 9664 1366 9716
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6144 9676 6745 9704
rect 6144 9664 6150 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 7098 9704 7104 9716
rect 6733 9667 6791 9673
rect 6932 9676 7104 9704
rect 2314 9596 2320 9648
rect 2372 9596 2378 9648
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 2832 9608 2877 9636
rect 2832 9596 2838 9608
rect 4430 9596 4436 9648
rect 4488 9596 4494 9648
rect 6178 9636 6184 9648
rect 6139 9608 6184 9636
rect 6178 9596 6184 9608
rect 6236 9596 6242 9648
rect 6549 9639 6607 9645
rect 6549 9605 6561 9639
rect 6595 9636 6607 9639
rect 6932 9636 6960 9676
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 6595 9608 6960 9636
rect 6595 9605 6607 9608
rect 6549 9599 6607 9605
rect 8018 9596 8024 9648
rect 8076 9596 8082 9648
rect 3234 9568 3240 9580
rect 3195 9540 3240 9568
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 5442 9568 5448 9580
rect 5399 9540 5448 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5551 9540 6377 9568
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9469 3111 9503
rect 3510 9500 3516 9512
rect 3471 9472 3516 9500
rect 3053 9463 3111 9469
rect 3068 9432 3096 9463
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 4062 9500 4068 9512
rect 3927 9472 4068 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 3068 9404 3556 9432
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2314 9364 2320 9376
rect 1728 9336 2320 9364
rect 1728 9324 1734 9336
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3528 9364 3556 9404
rect 4890 9392 4896 9444
rect 4948 9432 4954 9444
rect 5551 9432 5579 9540
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 6730 9500 6736 9512
rect 5960 9472 6736 9500
rect 5960 9460 5966 9472
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 6840 9500 6868 9531
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 6972 9540 7017 9568
rect 6972 9528 6978 9540
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8536 9540 8769 9568
rect 8536 9528 8542 9540
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 7006 9500 7012 9512
rect 6840 9472 7012 9500
rect 7006 9460 7012 9472
rect 7064 9460 7070 9512
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9500 7343 9503
rect 7834 9500 7840 9512
rect 7331 9472 7840 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 4948 9404 5579 9432
rect 4948 9392 4954 9404
rect 4430 9364 4436 9376
rect 3528 9336 4436 9364
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 5917 9367 5975 9373
rect 5917 9333 5929 9367
rect 5963 9364 5975 9367
rect 8662 9364 8668 9376
rect 5963 9336 8668 9364
rect 5963 9333 5975 9336
rect 5917 9327 5975 9333
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 9321 9367 9379 9373
rect 9321 9333 9333 9367
rect 9367 9364 9379 9367
rect 9582 9364 9588 9376
rect 9367 9336 9588 9364
rect 9367 9333 9379 9336
rect 9321 9327 9379 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 3053 9163 3111 9169
rect 3053 9129 3065 9163
rect 3099 9160 3111 9163
rect 3234 9160 3240 9172
rect 3099 9132 3240 9160
rect 3099 9129 3111 9132
rect 3053 9123 3111 9129
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 3973 9163 4031 9169
rect 3973 9160 3985 9163
rect 3568 9132 3985 9160
rect 3568 9120 3574 9132
rect 3973 9129 3985 9132
rect 4019 9129 4031 9163
rect 4154 9160 4160 9172
rect 4115 9132 4160 9160
rect 3973 9123 4031 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 5994 9160 6000 9172
rect 5767 9132 6000 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 7098 9160 7104 9172
rect 6236 9132 7104 9160
rect 6236 9120 6242 9132
rect 7098 9120 7104 9132
rect 7156 9160 7162 9172
rect 8202 9160 8208 9172
rect 7156 9132 8208 9160
rect 7156 9120 7162 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 4430 9052 4436 9104
rect 4488 9092 4494 9104
rect 5169 9095 5227 9101
rect 5169 9092 5181 9095
rect 4488 9064 5181 9092
rect 4488 9052 4494 9064
rect 5169 9061 5181 9064
rect 5215 9092 5227 9095
rect 6196 9092 6224 9120
rect 5215 9064 6224 9092
rect 8481 9095 8539 9101
rect 5215 9061 5227 9064
rect 5169 9055 5227 9061
rect 8481 9061 8493 9095
rect 8527 9092 8539 9095
rect 13722 9092 13728 9104
rect 8527 9064 13728 9092
rect 8527 9061 8539 9064
rect 8481 9055 8539 9061
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 1762 8984 1768 9036
rect 1820 9024 1826 9036
rect 6086 9024 6092 9036
rect 1820 8996 2774 9024
rect 1820 8984 1826 8996
rect 1302 8956 1308 8968
rect 1263 8928 1308 8956
rect 1302 8916 1308 8928
rect 1360 8916 1366 8968
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1995 8928 2053 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2746 8956 2774 8996
rect 3436 8996 3924 9024
rect 3436 8965 3464 8996
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 2746 8928 3433 8956
rect 2041 8919 2099 8925
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 3786 8956 3792 8968
rect 3747 8928 3792 8956
rect 3421 8919 3479 8925
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 3896 8965 3924 8996
rect 4632 8996 6092 9024
rect 4632 8965 4660 8996
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6236 8996 6281 9024
rect 6236 8984 6242 8996
rect 3881 8959 3939 8965
rect 3881 8925 3893 8959
rect 3927 8925 3939 8959
rect 3881 8919 3939 8925
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 1762 8848 1768 8900
rect 1820 8888 1826 8900
rect 2777 8891 2835 8897
rect 2777 8888 2789 8891
rect 1820 8860 2789 8888
rect 1820 8848 1826 8860
rect 2777 8857 2789 8860
rect 2823 8888 2835 8891
rect 2866 8888 2872 8900
rect 2823 8860 2872 8888
rect 2823 8857 2835 8860
rect 2777 8851 2835 8857
rect 2866 8848 2872 8860
rect 2924 8848 2930 8900
rect 2961 8891 3019 8897
rect 2961 8857 2973 8891
rect 3007 8888 3019 8891
rect 3234 8888 3240 8900
rect 3007 8860 3240 8888
rect 3007 8857 3019 8860
rect 2961 8851 3019 8857
rect 3234 8848 3240 8860
rect 3292 8848 3298 8900
rect 4356 8888 4384 8919
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 5074 8956 5080 8968
rect 4764 8928 5080 8956
rect 4764 8916 4770 8928
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5534 8956 5540 8968
rect 5495 8928 5540 8956
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 7558 8916 7564 8968
rect 7616 8956 7622 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 7616 8928 8309 8956
rect 7616 8916 7622 8928
rect 8297 8925 8309 8928
rect 8343 8956 8355 8959
rect 8754 8956 8760 8968
rect 8343 8928 8760 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 9180 8928 9321 8956
rect 9180 8916 9186 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 5353 8891 5411 8897
rect 4356 8860 4936 8888
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2280 8792 2697 8820
rect 2280 8780 2286 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 2685 8783 2743 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 3108 8792 3341 8820
rect 3108 8780 3114 8792
rect 3329 8789 3341 8792
rect 3375 8789 3387 8823
rect 3602 8820 3608 8832
rect 3563 8792 3608 8820
rect 3329 8783 3387 8789
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 4338 8820 4344 8832
rect 3752 8792 4344 8820
rect 3752 8780 3758 8792
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4908 8829 4936 8860
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 5810 8888 5816 8900
rect 5399 8860 5816 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 5810 8848 5816 8860
rect 5868 8848 5874 8900
rect 5997 8891 6055 8897
rect 5997 8857 6009 8891
rect 6043 8888 6055 8891
rect 6457 8891 6515 8897
rect 6043 8860 6224 8888
rect 6043 8857 6055 8860
rect 5997 8851 6055 8857
rect 6196 8832 6224 8860
rect 6457 8857 6469 8891
rect 6503 8888 6515 8891
rect 6546 8888 6552 8900
rect 6503 8860 6552 8888
rect 6503 8857 6515 8860
rect 6457 8851 6515 8857
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 7834 8848 7840 8900
rect 7892 8888 7898 8900
rect 8113 8891 8171 8897
rect 8113 8888 8125 8891
rect 7892 8860 8125 8888
rect 7892 8848 7898 8860
rect 8113 8857 8125 8860
rect 8159 8857 8171 8891
rect 8113 8851 8171 8857
rect 4893 8823 4951 8829
rect 4893 8789 4905 8823
rect 4939 8820 4951 8823
rect 4982 8820 4988 8832
rect 4939 8792 4988 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 5592 8792 5917 8820
rect 5592 8780 5598 8792
rect 5905 8789 5917 8792
rect 5951 8789 5963 8823
rect 5905 8783 5963 8789
rect 6178 8780 6184 8832
rect 6236 8780 6242 8832
rect 6362 8780 6368 8832
rect 6420 8820 6426 8832
rect 6822 8820 6828 8832
rect 6420 8792 6828 8820
rect 6420 8780 6426 8792
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7929 8823 7987 8829
rect 7929 8789 7941 8823
rect 7975 8820 7987 8823
rect 8018 8820 8024 8832
rect 7975 8792 8024 8820
rect 7975 8789 7987 8792
rect 7929 8783 7987 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8757 8823 8815 8829
rect 8757 8820 8769 8823
rect 8444 8792 8769 8820
rect 8444 8780 8450 8792
rect 8757 8789 8769 8792
rect 8803 8789 8815 8823
rect 8757 8783 8815 8789
rect 920 8730 9844 8752
rect 920 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 5194 8730
rect 5246 8678 5258 8730
rect 5310 8678 5322 8730
rect 5374 8678 9844 8730
rect 920 8656 9844 8678
rect 1762 8616 1768 8628
rect 1723 8588 1768 8616
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 3050 8616 3056 8628
rect 1872 8588 3056 8616
rect 1872 8489 1900 8588
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 3694 8616 3700 8628
rect 3200 8588 3700 8616
rect 3200 8576 3206 8588
rect 3694 8576 3700 8588
rect 3752 8616 3758 8628
rect 3752 8588 4752 8616
rect 3752 8576 3758 8588
rect 3602 8548 3608 8560
rect 3358 8520 3608 8548
rect 3602 8508 3608 8520
rect 3660 8508 3666 8560
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 4724 8557 4752 8588
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 6273 8619 6331 8625
rect 5040 8588 5856 8616
rect 5040 8576 5046 8588
rect 4709 8551 4767 8557
rect 4304 8520 4660 8548
rect 4304 8508 4310 8520
rect 4632 8492 4660 8520
rect 4709 8517 4721 8551
rect 4755 8517 4767 8551
rect 4890 8548 4896 8560
rect 4851 8520 4896 8548
rect 4709 8511 4767 8517
rect 4890 8508 4896 8520
rect 4948 8548 4954 8560
rect 5258 8548 5264 8560
rect 4948 8520 5264 8548
rect 4948 8508 4954 8520
rect 5258 8508 5264 8520
rect 5316 8548 5322 8560
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 5316 8520 5365 8548
rect 5316 8508 5322 8520
rect 5353 8517 5365 8520
rect 5399 8517 5411 8551
rect 5353 8511 5411 8517
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 2056 8452 2360 8480
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8412 1639 8415
rect 2056 8412 2084 8452
rect 2222 8412 2228 8424
rect 1627 8384 2084 8412
rect 2183 8384 2228 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2332 8412 2360 8452
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3476 8452 3709 8480
rect 3476 8440 3482 8452
rect 3697 8449 3709 8452
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 2866 8412 2872 8424
rect 2332 8384 2872 8412
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 4448 8412 4476 8443
rect 4614 8440 4620 8492
rect 4672 8480 4678 8492
rect 4672 8452 5396 8480
rect 4672 8440 4678 8452
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4448 8384 5181 8412
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5368 8412 5396 8452
rect 5442 8440 5448 8492
rect 5500 8482 5506 8492
rect 5828 8489 5856 8588
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6362 8616 6368 8628
rect 6319 8588 6368 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 6825 8619 6883 8625
rect 6825 8585 6837 8619
rect 6871 8616 6883 8619
rect 6914 8616 6920 8628
rect 6871 8588 6920 8616
rect 6871 8585 6883 8588
rect 6825 8579 6883 8585
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 7193 8619 7251 8625
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 7466 8616 7472 8628
rect 7239 8588 7472 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 9122 8616 9128 8628
rect 8536 8588 8984 8616
rect 9083 8588 9128 8616
rect 8536 8576 8542 8588
rect 5537 8483 5595 8489
rect 5537 8482 5549 8483
rect 5500 8454 5549 8482
rect 5500 8440 5506 8454
rect 5537 8449 5549 8454
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 5813 8483 5871 8489
rect 5675 8452 5764 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 5368 8384 5580 8412
rect 5169 8375 5227 8381
rect 4261 8347 4319 8353
rect 4261 8313 4273 8347
rect 4307 8344 4319 8347
rect 4798 8344 4804 8356
rect 4307 8316 4804 8344
rect 4307 8313 4319 8316
rect 4261 8307 4319 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5442 8344 5448 8356
rect 5123 8316 5448 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 5552 8344 5580 8384
rect 5736 8344 5764 8452
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5994 8480 6000 8492
rect 5859 8452 6000 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6328 8452 6377 8480
rect 6328 8440 6334 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6638 8440 6644 8492
rect 6696 8480 6702 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6696 8452 7021 8480
rect 6696 8440 6702 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7366 8483 7424 8489
rect 7366 8480 7378 8483
rect 7156 8452 7378 8480
rect 7156 8440 7162 8452
rect 7366 8449 7378 8452
rect 7412 8480 7424 8483
rect 7412 8449 7432 8480
rect 7366 8443 7432 8449
rect 7404 8356 7432 8443
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 8956 8480 8984 8588
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 8956 8452 9321 8480
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 9398 8412 9404 8424
rect 7699 8384 9404 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 5552 8316 5764 8344
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8344 6055 8347
rect 6730 8344 6736 8356
rect 6043 8316 6736 8344
rect 6043 8313 6055 8316
rect 5997 8307 6055 8313
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 7374 8304 7380 8356
rect 7432 8304 7438 8356
rect 9493 8347 9551 8353
rect 9493 8313 9505 8347
rect 9539 8344 9551 8347
rect 13630 8344 13636 8356
rect 9539 8316 13636 8344
rect 9539 8313 9551 8316
rect 9493 8307 9551 8313
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 1397 8279 1455 8285
rect 1397 8245 1409 8279
rect 1443 8276 1455 8279
rect 2406 8276 2412 8288
rect 1443 8248 2412 8276
rect 1443 8245 1455 8248
rect 1397 8239 1455 8245
rect 2406 8236 2412 8248
rect 2464 8236 2470 8288
rect 4617 8279 4675 8285
rect 4617 8245 4629 8279
rect 4663 8276 4675 8279
rect 4890 8276 4896 8288
rect 4663 8248 4896 8276
rect 4663 8245 4675 8248
rect 4617 8239 4675 8245
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 5224 8248 6469 8276
rect 5224 8236 5230 8248
rect 6457 8245 6469 8248
rect 6503 8276 6515 8279
rect 7282 8276 7288 8288
rect 6503 8248 7288 8276
rect 6503 8245 6515 8248
rect 6457 8239 6515 8245
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1544 8044 4200 8072
rect 1544 8032 1550 8044
rect 1578 7936 1584 7948
rect 1539 7908 1584 7936
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 1854 7936 1860 7948
rect 1815 7908 1860 7936
rect 1854 7896 1860 7908
rect 1912 7896 1918 7948
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 3329 7939 3387 7945
rect 2372 7908 3188 7936
rect 2372 7896 2378 7908
rect 3160 7880 3188 7908
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 3605 7939 3663 7945
rect 3605 7936 3617 7939
rect 3375 7908 3617 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 3605 7905 3617 7908
rect 3651 7905 3663 7939
rect 4172 7936 4200 8044
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 5166 8072 5172 8084
rect 4304 8044 5172 8072
rect 4304 8032 4310 8044
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 5721 8075 5779 8081
rect 5721 8072 5733 8075
rect 5316 8044 5733 8072
rect 5316 8032 5322 8044
rect 5721 8041 5733 8044
rect 5767 8041 5779 8075
rect 5721 8035 5779 8041
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6454 8072 6460 8084
rect 6144 8044 6460 8072
rect 6144 8032 6150 8044
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 8018 8032 8024 8084
rect 8076 8072 8082 8084
rect 9398 8072 9404 8084
rect 8076 8044 8800 8072
rect 9359 8044 9404 8072
rect 8076 8032 8082 8044
rect 5994 7964 6000 8016
rect 6052 8004 6058 8016
rect 7834 8004 7840 8016
rect 6052 7976 7840 8004
rect 6052 7964 6058 7976
rect 7834 7964 7840 7976
rect 7892 7964 7898 8016
rect 8110 8004 8116 8016
rect 8071 7976 8116 8004
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 5350 7936 5356 7948
rect 4172 7908 5356 7936
rect 3605 7899 3663 7905
rect 1486 7868 1492 7880
rect 1447 7840 1492 7868
rect 1486 7828 1492 7840
rect 1544 7828 1550 7880
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 5092 7877 5120 7908
rect 5350 7896 5356 7908
rect 5408 7936 5414 7948
rect 5718 7936 5724 7948
rect 5408 7908 5724 7936
rect 5408 7896 5414 7908
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 6328 7908 8524 7936
rect 6328 7896 6334 7908
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4295 7840 4353 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4341 7837 4353 7840
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6052 7840 6653 7868
rect 6052 7828 6058 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 7466 7868 7472 7880
rect 6641 7831 6699 7837
rect 6840 7840 7472 7868
rect 3160 7800 3188 7828
rect 4706 7800 4712 7812
rect 3082 7772 4712 7800
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 5644 7800 5672 7828
rect 6181 7803 6239 7809
rect 6181 7800 6193 7803
rect 5644 7772 6193 7800
rect 6181 7769 6193 7772
rect 6227 7769 6239 7803
rect 6181 7763 6239 7769
rect 6549 7803 6607 7809
rect 6549 7769 6561 7803
rect 6595 7800 6607 7803
rect 6840 7800 6868 7840
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8386 7868 8392 7880
rect 8067 7840 8392 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 8496 7877 8524 7908
rect 8772 7877 8800 8044
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 6595 7772 6868 7800
rect 6595 7769 6607 7772
rect 6549 7763 6607 7769
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7377 7803 7435 7809
rect 7377 7800 7389 7803
rect 6972 7772 7389 7800
rect 6972 7760 6978 7772
rect 7377 7769 7389 7772
rect 7423 7769 7435 7803
rect 7377 7763 7435 7769
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8297 7803 8355 7809
rect 8297 7800 8309 7803
rect 8168 7772 8309 7800
rect 8168 7760 8174 7772
rect 8297 7769 8309 7772
rect 8343 7769 8355 7803
rect 8496 7800 8524 7831
rect 9398 7800 9404 7812
rect 8496 7772 9404 7800
rect 8297 7763 8355 7769
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 3142 7732 3148 7744
rect 1443 7704 3148 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 3936 7704 4997 7732
rect 3936 7692 3942 7704
rect 4985 7701 4997 7704
rect 5031 7701 5043 7735
rect 4985 7695 5043 7701
rect 5537 7735 5595 7741
rect 5537 7701 5549 7735
rect 5583 7732 5595 7735
rect 5626 7732 5632 7744
rect 5583 7704 5632 7732
rect 5583 7701 5595 7704
rect 5537 7695 5595 7701
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 6086 7732 6092 7744
rect 6047 7704 6092 7732
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6270 7732 6276 7744
rect 6231 7704 6276 7732
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 6420 7704 6465 7732
rect 6420 7692 6426 7704
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7064 7704 7297 7732
rect 7064 7692 7070 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7285 7695 7343 7701
rect 7834 7692 7840 7744
rect 7892 7732 7898 7744
rect 9306 7732 9312 7744
rect 7892 7704 9312 7732
rect 7892 7692 7898 7704
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 920 7642 9844 7664
rect 920 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 5194 7642
rect 5246 7590 5258 7642
rect 5310 7590 5322 7642
rect 5374 7590 9844 7642
rect 920 7568 9844 7590
rect 1302 7528 1308 7540
rect 1263 7500 1308 7528
rect 1302 7488 1308 7500
rect 1360 7488 1366 7540
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 4522 7528 4528 7540
rect 1544 7500 4528 7528
rect 1544 7488 1550 7500
rect 2314 7420 2320 7472
rect 2372 7420 2378 7472
rect 2774 7460 2780 7472
rect 2735 7432 2780 7460
rect 2774 7420 2780 7432
rect 2832 7420 2838 7472
rect 3068 7392 3096 7500
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 7190 7528 7196 7540
rect 6564 7500 7196 7528
rect 4988 7472 5040 7478
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 3200 7432 3556 7460
rect 3200 7420 3206 7432
rect 3528 7401 3556 7432
rect 4988 7414 5040 7420
rect 3237 7395 3295 7401
rect 3237 7392 3249 7395
rect 3068 7364 3249 7392
rect 3237 7361 3249 7364
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7361 3571 7395
rect 3878 7392 3884 7404
rect 3839 7364 3884 7392
rect 3513 7355 3571 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 4890 7352 4896 7404
rect 4948 7382 4954 7404
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 5092 7382 5365 7392
rect 4948 7364 5365 7382
rect 4948 7354 5120 7364
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 4948 7352 4954 7354
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 6564 7401 6592 7500
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 7616 7500 9137 7528
rect 7616 7488 7622 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9398 7528 9404 7540
rect 9359 7500 9404 7528
rect 9125 7491 9183 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 8294 7460 8300 7472
rect 8050 7432 8300 7460
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 5500 7364 6377 7392
rect 5500 7352 5506 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 6549 7355 6607 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 8260 7364 8401 7392
rect 8260 7352 8266 7364
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 9306 7392 9312 7404
rect 9267 7364 9312 7392
rect 8389 7355 8447 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 1544 7296 3065 7324
rect 1544 7284 1550 7296
rect 3053 7293 3065 7296
rect 3099 7324 3111 7327
rect 4430 7324 4436 7336
rect 3099 7296 4436 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 7282 7284 7288 7336
rect 7340 7324 7346 7336
rect 7558 7324 7564 7336
rect 7340 7296 7564 7324
rect 7340 7284 7346 7296
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 5917 7259 5975 7265
rect 5917 7225 5929 7259
rect 5963 7256 5975 7259
rect 6362 7256 6368 7268
rect 5963 7228 6368 7256
rect 5963 7225 5975 7228
rect 5917 7219 5975 7225
rect 6362 7216 6368 7228
rect 6420 7256 6426 7268
rect 8754 7256 8760 7268
rect 6420 7228 6696 7256
rect 6420 7216 6426 7228
rect 3326 7188 3332 7200
rect 3287 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 6144 7160 6193 7188
rect 6144 7148 6150 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 6668 7188 6696 7228
rect 7852 7228 8760 7256
rect 7852 7188 7880 7228
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 6668 7160 7880 7188
rect 8573 7191 8631 7197
rect 6181 7151 6239 7157
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 8846 7188 8852 7200
rect 8619 7160 8852 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 8938 7148 8944 7200
rect 8996 7197 9002 7200
rect 8996 7188 9007 7197
rect 8996 7160 9041 7188
rect 8996 7151 9007 7160
rect 8996 7148 9002 7151
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 1752 6987 1810 6993
rect 1752 6953 1764 6987
rect 1798 6984 1810 6987
rect 2222 6984 2228 6996
rect 1798 6956 2228 6984
rect 1798 6953 1810 6956
rect 1752 6947 1810 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 6362 6984 6368 6996
rect 5960 6956 6368 6984
rect 5960 6944 5966 6956
rect 6362 6944 6368 6956
rect 6420 6944 6426 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7389 6987 7447 6993
rect 7389 6984 7401 6987
rect 6972 6956 7401 6984
rect 6972 6944 6978 6956
rect 7389 6953 7401 6956
rect 7435 6953 7447 6987
rect 7389 6947 7447 6953
rect 8662 6944 8668 6996
rect 8720 6984 8726 6996
rect 8849 6987 8907 6993
rect 8849 6984 8861 6987
rect 8720 6956 8861 6984
rect 8720 6944 8726 6956
rect 8849 6953 8861 6956
rect 8895 6984 8907 6987
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 8895 6956 9413 6984
rect 8895 6953 8907 6956
rect 8849 6947 8907 6953
rect 9401 6953 9413 6956
rect 9447 6984 9459 6987
rect 9490 6984 9496 6996
rect 9447 6956 9496 6984
rect 9447 6953 9459 6956
rect 9401 6947 9459 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3605 6851 3663 6857
rect 3605 6848 3617 6851
rect 3283 6820 3617 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3605 6817 3617 6820
rect 3651 6817 3663 6851
rect 3605 6811 3663 6817
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4341 6851 4399 6857
rect 4341 6848 4353 6851
rect 4120 6820 4353 6848
rect 4120 6808 4126 6820
rect 4341 6817 4353 6820
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 5905 6851 5963 6857
rect 5905 6817 5917 6851
rect 5951 6817 5963 6851
rect 5905 6811 5963 6817
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 4080 6780 4108 6808
rect 3200 6752 4108 6780
rect 4249 6783 4307 6789
rect 3200 6740 3206 6752
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4295 6752 4997 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5920 6780 5948 6811
rect 7374 6808 7380 6860
rect 7432 6848 7438 6860
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7432 6820 7665 6848
rect 7432 6808 7438 6820
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 13722 6848 13728 6860
rect 8251 6820 13728 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 5123 6752 5948 6780
rect 7668 6752 7849 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 3050 6712 3056 6724
rect 2990 6684 3056 6712
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 7466 6712 7472 6724
rect 6946 6684 7472 6712
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 1397 6647 1455 6653
rect 1397 6613 1409 6647
rect 1443 6644 1455 6647
rect 1486 6644 1492 6656
rect 1443 6616 1492 6644
rect 1443 6613 1455 6616
rect 1397 6607 1455 6613
rect 1486 6604 1492 6616
rect 1544 6644 1550 6656
rect 3068 6644 3096 6672
rect 3510 6644 3516 6656
rect 1544 6616 3516 6644
rect 1544 6604 1550 6616
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 5721 6647 5779 6653
rect 5721 6613 5733 6647
rect 5767 6644 5779 6647
rect 5902 6644 5908 6656
rect 5767 6616 5908 6644
rect 5767 6613 5779 6616
rect 5721 6607 5779 6613
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 7668 6644 7696 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6749 8079 6783
rect 8294 6780 8300 6792
rect 8255 6752 8300 6780
rect 8021 6743 8079 6749
rect 8036 6712 8064 6743
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8570 6780 8576 6792
rect 8531 6752 8576 6780
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 8754 6780 8760 6792
rect 8715 6752 8760 6780
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 9030 6712 9036 6724
rect 8036 6684 9036 6712
rect 9030 6672 9036 6684
rect 9088 6672 9094 6724
rect 8386 6644 8392 6656
rect 6696 6616 8392 6644
rect 6696 6604 6702 6616
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6644 9275 6647
rect 9306 6644 9312 6656
rect 9263 6616 9312 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 920 6554 9844 6576
rect 920 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 5194 6554
rect 5246 6502 5258 6554
rect 5310 6502 5322 6554
rect 5374 6502 9844 6554
rect 920 6480 9844 6502
rect 1397 6443 1455 6449
rect 1397 6409 1409 6443
rect 1443 6440 1455 6443
rect 1486 6440 1492 6452
rect 1443 6412 1492 6440
rect 1443 6409 1455 6412
rect 1397 6403 1455 6409
rect 1486 6400 1492 6412
rect 1544 6400 1550 6452
rect 5534 6440 5540 6452
rect 3068 6412 5540 6440
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 2958 6304 2964 6316
rect 2823 6276 2964 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3068 6313 3096 6412
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5776 6412 5917 6440
rect 5776 6400 5782 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 5905 6403 5963 6409
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 6638 6440 6644 6452
rect 6420 6412 6644 6440
rect 6420 6400 6426 6412
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 4062 6332 4068 6384
rect 4120 6332 4126 6384
rect 7926 6372 7932 6384
rect 7887 6344 7932 6372
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 8205 6375 8263 6381
rect 8205 6372 8217 6375
rect 8168 6344 8217 6372
rect 8168 6332 8174 6344
rect 8205 6341 8217 6344
rect 8251 6341 8263 6375
rect 8205 6335 8263 6341
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 8573 6375 8631 6381
rect 8573 6372 8585 6375
rect 8352 6344 8585 6372
rect 8352 6332 8358 6344
rect 8573 6341 8585 6344
rect 8619 6341 8631 6375
rect 8573 6335 8631 6341
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6273 3111 6307
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 3053 6267 3111 6273
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 6086 6304 6092 6316
rect 5215 6276 6092 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7156 6276 8033 6304
rect 7156 6264 7162 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 2682 6236 2688 6248
rect 2643 6208 2688 6236
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6236 3755 6239
rect 3970 6236 3976 6248
rect 3743 6208 3976 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 6178 6236 6184 6248
rect 6139 6208 6184 6236
rect 6178 6196 6184 6208
rect 6236 6196 6242 6248
rect 8036 6236 8064 6267
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8444 6276 8493 6304
rect 8444 6264 8450 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8754 6304 8760 6316
rect 8715 6276 8760 6304
rect 8481 6267 8539 6273
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8904 6276 8953 6304
rect 8904 6264 8910 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9858 6304 9864 6316
rect 9355 6276 9864 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 8036 6208 9413 6236
rect 9401 6205 9413 6208
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 2317 6171 2375 6177
rect 2317 6137 2329 6171
rect 2363 6168 2375 6171
rect 2961 6171 3019 6177
rect 2363 6140 2774 6168
rect 2363 6137 2375 6140
rect 2317 6131 2375 6137
rect 2406 6100 2412 6112
rect 2367 6072 2412 6100
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2746 6100 2774 6140
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 5733 6171 5791 6177
rect 3007 6140 3464 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 3050 6100 3056 6112
rect 2746 6072 3056 6100
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 3234 6100 3240 6112
rect 3195 6072 3240 6100
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 3436 6100 3464 6140
rect 5733 6137 5745 6171
rect 5779 6168 5791 6171
rect 8202 6168 8208 6180
rect 5779 6140 8208 6168
rect 5779 6137 5791 6140
rect 5733 6131 5791 6137
rect 8202 6128 8208 6140
rect 8260 6128 8266 6180
rect 8662 6128 8668 6180
rect 8720 6168 8726 6180
rect 8720 6140 12434 6168
rect 8720 6128 8726 6140
rect 4062 6100 4068 6112
rect 3436 6072 4068 6100
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 9214 6100 9220 6112
rect 8343 6072 9220 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 12406 6100 12434 6140
rect 13446 6100 13452 6112
rect 12406 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 1486 5896 1492 5908
rect 1447 5868 1492 5896
rect 1486 5856 1492 5868
rect 1544 5856 1550 5908
rect 1670 5896 1676 5908
rect 1631 5868 1676 5896
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3016 5868 3893 5896
rect 3016 5856 3022 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 3881 5859 3939 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 8018 5896 8024 5908
rect 7340 5868 8024 5896
rect 7340 5856 7346 5868
rect 8018 5856 8024 5868
rect 8076 5896 8082 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 8076 5868 8125 5896
rect 8076 5856 8082 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8628 5868 8861 5896
rect 8628 5856 8634 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 3694 5828 3700 5840
rect 3655 5800 3700 5828
rect 3694 5788 3700 5800
rect 3752 5788 3758 5840
rect 5905 5831 5963 5837
rect 5905 5797 5917 5831
rect 5951 5828 5963 5831
rect 8662 5828 8668 5840
rect 5951 5800 8668 5828
rect 5951 5797 5963 5800
rect 5905 5791 5963 5797
rect 8662 5788 8668 5800
rect 8720 5788 8726 5840
rect 8754 5788 8760 5840
rect 8812 5828 8818 5840
rect 9217 5831 9275 5837
rect 9217 5828 9229 5831
rect 8812 5800 9229 5828
rect 8812 5788 8818 5800
rect 9217 5797 9229 5800
rect 9263 5797 9275 5831
rect 9217 5791 9275 5797
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 9490 5828 9496 5840
rect 9364 5800 9496 5828
rect 9364 5788 9370 5800
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 1305 5763 1363 5769
rect 1305 5729 1317 5763
rect 1351 5760 1363 5763
rect 1351 5732 5776 5760
rect 1351 5729 1363 5732
rect 1305 5723 1363 5729
rect 3418 5652 3424 5704
rect 3476 5692 3482 5704
rect 3476 5664 3521 5692
rect 3476 5652 3482 5664
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 3752 5664 4353 5692
rect 3752 5652 3758 5664
rect 4341 5661 4353 5664
rect 4387 5661 4399 5695
rect 4341 5655 4399 5661
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5661 4491 5695
rect 4433 5655 4491 5661
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5661 5687 5695
rect 5748 5692 5776 5732
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 5868 5732 6193 5760
rect 5868 5720 5874 5732
rect 6181 5729 6193 5732
rect 6227 5729 6239 5763
rect 6181 5723 6239 5729
rect 6822 5720 6828 5772
rect 6880 5760 6886 5772
rect 6880 5732 7972 5760
rect 6880 5720 6886 5732
rect 7944 5692 7972 5732
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 13814 5760 13820 5772
rect 8352 5732 13820 5760
rect 8352 5720 8358 5732
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 5748 5664 7880 5692
rect 7944 5664 8033 5692
rect 5629 5655 5687 5661
rect 1486 5584 1492 5636
rect 1544 5624 1550 5636
rect 3142 5624 3148 5636
rect 1544 5596 1978 5624
rect 3103 5596 3148 5624
rect 1544 5584 1550 5596
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 4448 5624 4476 5655
rect 3252 5596 4476 5624
rect 5644 5624 5672 5655
rect 7466 5624 7472 5636
rect 5644 5596 7472 5624
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 3252 5556 3280 5596
rect 7466 5584 7472 5596
rect 7524 5584 7530 5636
rect 7852 5624 7880 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 9030 5692 9036 5704
rect 8991 5664 9036 5692
rect 8021 5655 8079 5661
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5692 9367 5695
rect 9858 5692 9864 5704
rect 9355 5664 9864 5692
rect 9355 5661 9367 5664
rect 9309 5655 9367 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 7929 5627 7987 5633
rect 7929 5624 7941 5627
rect 7852 5596 7941 5624
rect 7929 5593 7941 5596
rect 7975 5624 7987 5627
rect 7975 5596 8064 5624
rect 7975 5593 7987 5596
rect 7929 5587 7987 5593
rect 2832 5528 3280 5556
rect 8036 5556 8064 5596
rect 8294 5556 8300 5568
rect 8036 5528 8300 5556
rect 2832 5516 2838 5528
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 920 5466 9844 5488
rect 920 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 5194 5466
rect 5246 5414 5258 5466
rect 5310 5414 5322 5466
rect 5374 5414 9844 5466
rect 920 5392 9844 5414
rect 2406 5312 2412 5364
rect 2464 5352 2470 5364
rect 4614 5352 4620 5364
rect 2464 5324 4620 5352
rect 2464 5312 2470 5324
rect 4614 5312 4620 5324
rect 4672 5352 4678 5364
rect 6454 5352 6460 5364
rect 4672 5324 5304 5352
rect 6415 5324 6460 5352
rect 4672 5312 4678 5324
rect 3234 5244 3240 5296
rect 3292 5284 3298 5296
rect 5169 5287 5227 5293
rect 5169 5284 5181 5287
rect 3292 5256 5181 5284
rect 3292 5244 3298 5256
rect 5169 5253 5181 5256
rect 5215 5253 5227 5287
rect 5169 5247 5227 5253
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3108 5188 3341 5216
rect 3108 5176 3114 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5276 5216 5304 5324
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 6604 5324 7481 5352
rect 6604 5312 6610 5324
rect 7469 5321 7481 5324
rect 7515 5321 7527 5355
rect 7469 5315 7527 5321
rect 8110 5312 8116 5364
rect 8168 5312 8174 5364
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 6270 5284 6276 5296
rect 5592 5256 6276 5284
rect 5592 5244 5598 5256
rect 6270 5244 6276 5256
rect 6328 5284 6334 5296
rect 7193 5287 7251 5293
rect 7193 5284 7205 5287
rect 6328 5256 7205 5284
rect 6328 5244 6334 5256
rect 7193 5253 7205 5256
rect 7239 5284 7251 5287
rect 8128 5284 8156 5312
rect 7239 5256 8156 5284
rect 7239 5253 7251 5256
rect 7193 5247 7251 5253
rect 8754 5244 8760 5296
rect 8812 5284 8818 5296
rect 8941 5287 8999 5293
rect 8941 5284 8953 5287
rect 8812 5256 8953 5284
rect 8812 5244 8818 5256
rect 8941 5253 8953 5256
rect 8987 5253 8999 5287
rect 8941 5247 8999 5253
rect 5123 5188 5304 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 4356 5148 4384 5179
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6086 5216 6092 5228
rect 5684 5188 6092 5216
rect 5684 5176 5690 5188
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6880 5188 7021 5216
rect 6880 5176 6886 5188
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 8110 5216 8116 5228
rect 8071 5188 8116 5216
rect 7009 5179 7067 5185
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8386 5216 8392 5228
rect 8343 5188 8392 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 9355 5188 12434 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 6178 5148 6184 5160
rect 4356 5120 6184 5148
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 9140 5148 9168 5179
rect 6420 5120 9536 5148
rect 6420 5108 6426 5120
rect 4154 5080 4160 5092
rect 4115 5052 4160 5080
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 7377 5083 7435 5089
rect 7377 5049 7389 5083
rect 7423 5080 7435 5083
rect 8202 5080 8208 5092
rect 7423 5052 8208 5080
rect 7423 5049 7435 5052
rect 7377 5043 7435 5049
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 3970 5012 3976 5024
rect 3931 4984 3976 5012
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4614 5012 4620 5024
rect 4575 4984 4620 5012
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4798 5012 4804 5024
rect 4759 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 8076 4984 8401 5012
rect 8076 4972 8082 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 8754 5012 8760 5024
rect 8715 4984 8760 5012
rect 8389 4975 8447 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 9508 5021 9536 5120
rect 9493 5015 9551 5021
rect 9493 4981 9505 5015
rect 9539 5012 9551 5015
rect 9582 5012 9588 5024
rect 9539 4984 9588 5012
rect 9539 4981 9551 4984
rect 9493 4975 9551 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 3326 4808 3332 4820
rect 3287 4780 3332 4808
rect 3326 4768 3332 4780
rect 3384 4808 3390 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3384 4780 3801 4808
rect 3384 4768 3390 4780
rect 3789 4777 3801 4780
rect 3835 4808 3847 4811
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 3835 4780 4445 4808
rect 3835 4777 3847 4780
rect 3789 4771 3847 4777
rect 4433 4777 4445 4780
rect 4479 4808 4491 4811
rect 4798 4808 4804 4820
rect 4479 4780 4804 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 5040 4780 6193 4808
rect 5040 4768 5046 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 7098 4808 7104 4820
rect 6181 4771 6239 4777
rect 6564 4780 7104 4808
rect 6564 4740 6592 4780
rect 7098 4768 7104 4780
rect 7156 4808 7162 4820
rect 8386 4808 8392 4820
rect 7156 4780 8392 4808
rect 7156 4768 7162 4780
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 8861 4811 8919 4817
rect 8861 4777 8873 4811
rect 8907 4808 8919 4811
rect 9876 4808 9904 5188
rect 8907 4780 9904 4808
rect 12406 4808 12434 5188
rect 13814 4808 13820 4820
rect 12406 4780 13820 4808
rect 8907 4777 8919 4780
rect 8861 4771 8919 4777
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 6012 4712 6592 4740
rect 8312 4712 9045 4740
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 5718 4672 5724 4684
rect 4847 4644 5724 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 3510 4604 3516 4616
rect 3471 4576 3516 4604
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 3697 4607 3755 4613
rect 3697 4604 3709 4607
rect 3660 4576 3709 4604
rect 3660 4564 3666 4576
rect 3697 4573 3709 4576
rect 3743 4573 3755 4607
rect 4338 4604 4344 4616
rect 4299 4576 4344 4604
rect 3697 4567 3755 4573
rect 3712 4536 3740 4567
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 4522 4564 4528 4616
rect 4580 4604 4586 4616
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 4580 4576 5365 4604
rect 4580 4564 4586 4576
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 6012 4604 6040 4712
rect 6086 4632 6092 4684
rect 6144 4672 6150 4684
rect 6825 4675 6883 4681
rect 6144 4644 6408 4672
rect 6144 4632 6150 4644
rect 6380 4613 6408 4644
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7006 4672 7012 4684
rect 6871 4644 7012 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 5583 4576 6040 4604
rect 6365 4607 6423 4613
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6454 4564 6460 4616
rect 6512 4604 6518 4616
rect 8312 4613 8340 4712
rect 9033 4709 9045 4712
rect 9079 4709 9091 4743
rect 9033 4703 9091 4709
rect 8754 4632 8760 4684
rect 8812 4672 8818 4684
rect 8812 4644 9536 4672
rect 8812 4632 8818 4644
rect 8297 4607 8355 4613
rect 6512 4576 6557 4604
rect 6512 4564 6518 4576
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 9214 4604 9220 4616
rect 9175 4576 9220 4604
rect 8297 4567 8355 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9508 4613 9536 4644
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 4985 4539 5043 4545
rect 4985 4536 4997 4539
rect 3712 4508 4997 4536
rect 4985 4505 4997 4508
rect 5031 4505 5043 4539
rect 4985 4499 5043 4505
rect 5169 4539 5227 4545
rect 5169 4505 5181 4539
rect 5215 4536 5227 4539
rect 5442 4536 5448 4548
rect 5215 4508 5448 4536
rect 5215 4505 5227 4508
rect 5169 4499 5227 4505
rect 5442 4496 5448 4508
rect 5500 4496 5506 4548
rect 5721 4539 5779 4545
rect 5721 4536 5733 4539
rect 5644 4508 5733 4536
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 4246 4468 4252 4480
rect 4203 4440 4252 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 5644 4468 5672 4508
rect 5721 4505 5733 4508
rect 5767 4505 5779 4539
rect 5721 4499 5779 4505
rect 5905 4539 5963 4545
rect 5905 4505 5917 4539
rect 5951 4505 5963 4539
rect 5905 4499 5963 4505
rect 4396 4440 5672 4468
rect 5920 4468 5948 4499
rect 5994 4496 6000 4548
rect 6052 4536 6058 4548
rect 6089 4539 6147 4545
rect 6089 4536 6101 4539
rect 6052 4508 6101 4536
rect 6052 4496 6058 4508
rect 6089 4505 6101 4508
rect 6135 4505 6147 4539
rect 7958 4508 9352 4536
rect 6089 4499 6147 4505
rect 6270 4468 6276 4480
rect 5920 4440 6276 4468
rect 4396 4428 4402 4440
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 9324 4477 9352 4508
rect 9309 4471 9367 4477
rect 9309 4437 9321 4471
rect 9355 4437 9367 4471
rect 9309 4431 9367 4437
rect 3036 4378 9844 4400
rect 3036 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 5194 4378
rect 5246 4326 5258 4378
rect 5310 4326 5322 4378
rect 5374 4326 9844 4378
rect 3036 4304 9844 4326
rect 3510 4224 3516 4276
rect 3568 4264 3574 4276
rect 3694 4264 3700 4276
rect 3568 4236 3700 4264
rect 3568 4224 3574 4236
rect 3694 4224 3700 4236
rect 3752 4224 3758 4276
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 9125 4267 9183 4273
rect 9125 4264 9137 4267
rect 7524 4236 9137 4264
rect 7524 4224 7530 4236
rect 9125 4233 9137 4236
rect 9171 4233 9183 4267
rect 9125 4227 9183 4233
rect 4154 4196 4160 4208
rect 3896 4168 4160 4196
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4128 3663 4131
rect 3896 4128 3924 4168
rect 4154 4156 4160 4168
rect 4212 4156 4218 4208
rect 4246 4156 4252 4208
rect 4304 4156 4310 4208
rect 5350 4156 5356 4208
rect 5408 4156 5414 4208
rect 6546 4156 6552 4208
rect 6604 4196 6610 4208
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 6604 4168 6929 4196
rect 6604 4156 6610 4168
rect 6917 4165 6929 4168
rect 6963 4165 6975 4199
rect 6917 4159 6975 4165
rect 3651 4100 3924 4128
rect 3973 4131 4031 4137
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4264 4128 4292 4156
rect 6086 4128 6092 4140
rect 4019 4100 4292 4128
rect 6047 4100 6092 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4128 7251 4131
rect 8113 4131 8171 4137
rect 7239 4100 7420 4128
rect 7239 4097 7251 4100
rect 7193 4091 7251 4097
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 3559 4032 4261 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4338 4020 4344 4072
rect 4396 4020 4402 4072
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 4798 4060 4804 4072
rect 4663 4032 4804 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 6512 4032 7297 4060
rect 6512 4020 6518 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 4120 3896 4169 3924
rect 4120 3884 4126 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4356 3924 4384 4020
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 5592 3964 7113 3992
rect 5592 3952 5598 3964
rect 7101 3961 7113 3964
rect 7147 3992 7159 3995
rect 7392 3992 7420 4100
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8159 4100 8309 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9493 4131 9551 4137
rect 9272 4100 9317 4128
rect 9272 4088 9278 4100
rect 9493 4097 9505 4131
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8444 4032 8861 4060
rect 8444 4020 8450 4032
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 7147 3964 7420 3992
rect 7147 3961 7159 3964
rect 7101 3955 7159 3961
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 9508 3992 9536 4091
rect 8260 3964 9536 3992
rect 8260 3952 8266 3964
rect 5994 3924 6000 3936
rect 4356 3896 6000 3924
rect 4157 3887 4215 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6653 3927 6711 3933
rect 6653 3893 6665 3927
rect 6699 3924 6711 3927
rect 6822 3924 6828 3936
rect 6699 3896 6828 3924
rect 6699 3893 6711 3896
rect 6653 3887 6711 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7466 3924 7472 3936
rect 7427 3896 7472 3924
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 9306 3924 9312 3936
rect 9267 3896 9312 3924
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 3329 3723 3387 3729
rect 3329 3689 3341 3723
rect 3375 3720 3387 3723
rect 3602 3720 3608 3732
rect 3375 3692 3608 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 4338 3720 4344 3732
rect 4120 3692 4344 3720
rect 4120 3680 4126 3692
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 6086 3720 6092 3732
rect 4479 3692 6092 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 6457 3723 6515 3729
rect 6457 3720 6469 3723
rect 6328 3692 6469 3720
rect 6328 3680 6334 3692
rect 6457 3689 6469 3692
rect 6503 3689 6515 3723
rect 6457 3683 6515 3689
rect 9137 3723 9195 3729
rect 9137 3689 9149 3723
rect 9183 3720 9195 3723
rect 9858 3720 9864 3732
rect 9183 3692 9864 3720
rect 9183 3689 9195 3692
rect 9137 3683 9195 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 4801 3655 4859 3661
rect 4801 3652 4813 3655
rect 3476 3624 4813 3652
rect 3476 3612 3482 3624
rect 4801 3621 4813 3624
rect 4847 3621 4859 3655
rect 5721 3655 5779 3661
rect 5721 3652 5733 3655
rect 4801 3615 4859 3621
rect 5000 3624 5733 3652
rect 4154 3584 4160 3596
rect 3896 3556 4160 3584
rect 3896 3525 3924 3556
rect 4154 3544 4160 3556
rect 4212 3584 4218 3596
rect 4890 3584 4896 3596
rect 4212 3556 4896 3584
rect 4212 3544 4218 3556
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 4246 3516 4252 3528
rect 4207 3488 4252 3516
rect 3973 3479 4031 3485
rect 3988 3448 4016 3479
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 4522 3516 4528 3528
rect 4483 3488 4528 3516
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 5000 3516 5028 3624
rect 5721 3621 5733 3624
rect 5767 3621 5779 3655
rect 5721 3615 5779 3621
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 5491 3556 6745 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 6733 3553 6745 3556
rect 6779 3553 6791 3587
rect 6733 3547 6791 3553
rect 7101 3587 7159 3593
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 7466 3584 7472 3596
rect 7147 3556 7472 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 5534 3516 5540 3528
rect 4856 3488 5028 3516
rect 5495 3488 5540 3516
rect 4856 3476 4862 3488
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 5684 3488 6377 3516
rect 5684 3476 5690 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6638 3516 6644 3528
rect 6599 3488 6644 3516
rect 6365 3479 6423 3485
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 9306 3516 9312 3528
rect 8619 3488 9312 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9456 3488 9505 3516
rect 9456 3476 9462 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 4614 3448 4620 3460
rect 3988 3420 4620 3448
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 4985 3451 5043 3457
rect 4985 3417 4997 3451
rect 5031 3448 5043 3451
rect 5810 3448 5816 3460
rect 5031 3420 5816 3448
rect 5031 3417 5043 3420
rect 4985 3411 5043 3417
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 8294 3448 8300 3460
rect 8234 3420 8300 3448
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 3660 3352 3801 3380
rect 3660 3340 3666 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 3789 3343 3847 3349
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4246 3380 4252 3392
rect 4203 3352 4252 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4706 3380 4712 3392
rect 4667 3352 4712 3380
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 5261 3383 5319 3389
rect 5261 3349 5273 3383
rect 5307 3380 5319 3383
rect 6914 3380 6920 3392
rect 5307 3352 6920 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 9306 3380 9312 3392
rect 9267 3352 9312 3380
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 3036 3290 9844 3312
rect 3036 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 5194 3290
rect 5246 3238 5258 3290
rect 5310 3238 5322 3290
rect 5374 3238 9844 3290
rect 3036 3216 9844 3238
rect 3513 3179 3571 3185
rect 3513 3145 3525 3179
rect 3559 3176 3571 3179
rect 4430 3176 4436 3188
rect 3559 3148 4436 3176
rect 3559 3145 3571 3148
rect 3513 3139 3571 3145
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 4764 3148 5212 3176
rect 4764 3136 4770 3148
rect 4338 3068 4344 3120
rect 4396 3068 4402 3120
rect 3602 3040 3608 3052
rect 3563 3012 3608 3040
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 5184 3040 5212 3148
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5718 3176 5724 3188
rect 5592 3148 5724 3176
rect 5592 3136 5598 3148
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 8294 3176 8300 3188
rect 8255 3148 8300 3176
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 9306 3136 9312 3188
rect 9364 3136 9370 3188
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 5960 3080 6561 3108
rect 5960 3068 5966 3080
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 6549 3071 6607 3077
rect 7282 3068 7288 3120
rect 7340 3068 7346 3120
rect 8849 3111 8907 3117
rect 8849 3077 8861 3111
rect 8895 3108 8907 3111
rect 9324 3108 9352 3136
rect 8895 3080 9352 3108
rect 8895 3077 8907 3080
rect 8849 3071 8907 3077
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 5184 3012 5457 3040
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 8478 3040 8484 3052
rect 8439 3012 8484 3040
rect 5445 3003 5503 3009
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3620 2944 3985 2972
rect 3620 2916 3648 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 6273 2975 6331 2981
rect 6273 2972 6285 2975
rect 6236 2944 6285 2972
rect 6236 2932 6242 2944
rect 6273 2941 6285 2944
rect 6319 2941 6331 2975
rect 6273 2935 6331 2941
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8386 2972 8392 2984
rect 8067 2944 8392 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 8754 2972 8760 2984
rect 8667 2944 8760 2972
rect 8754 2932 8760 2944
rect 8812 2972 8818 2984
rect 9214 2972 9220 2984
rect 8812 2944 9220 2972
rect 8812 2932 8818 2944
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9398 2972 9404 2984
rect 9359 2944 9404 2972
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 3602 2864 3608 2916
rect 3660 2864 3666 2916
rect 4430 2796 4436 2848
rect 4488 2836 4494 2848
rect 4706 2836 4712 2848
rect 4488 2808 4712 2836
rect 4488 2796 4494 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 6009 2839 6067 2845
rect 6009 2805 6021 2839
rect 6055 2836 6067 2839
rect 6362 2836 6368 2848
rect 6055 2808 6368 2836
rect 6055 2805 6067 2808
rect 6009 2799 6067 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 3036 2672 9844 2694
rect 5353 2635 5411 2641
rect 5353 2601 5365 2635
rect 5399 2632 5411 2635
rect 5442 2632 5448 2644
rect 5399 2604 5448 2632
rect 5399 2601 5411 2604
rect 5353 2595 5411 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 8121 2635 8179 2641
rect 8121 2601 8133 2635
rect 8167 2601 8179 2635
rect 8121 2595 8179 2601
rect 5077 2567 5135 2573
rect 5077 2533 5089 2567
rect 5123 2564 5135 2567
rect 5626 2564 5632 2576
rect 5123 2536 5632 2564
rect 5123 2533 5135 2536
rect 5077 2527 5135 2533
rect 5626 2524 5632 2536
rect 5684 2524 5690 2576
rect 8128 2564 8156 2595
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 9088 2604 9137 2632
rect 9088 2592 9094 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 8202 2564 8208 2576
rect 8128 2536 8208 2564
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 3326 2496 3332 2508
rect 3287 2468 3332 2496
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 5442 2456 5448 2508
rect 5500 2496 5506 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5500 2468 5733 2496
rect 5500 2456 5506 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 8110 2456 8116 2508
rect 8168 2496 8174 2508
rect 8297 2499 8355 2505
rect 8297 2496 8309 2499
rect 8168 2468 8309 2496
rect 8168 2456 8174 2468
rect 8297 2465 8309 2468
rect 8343 2465 8355 2499
rect 8297 2459 8355 2465
rect 5534 2428 5540 2440
rect 5495 2400 5540 2428
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 6086 2428 6092 2440
rect 6047 2400 6092 2428
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 3602 2360 3608 2372
rect 3563 2332 3608 2360
rect 3602 2320 3608 2332
rect 3660 2320 3666 2372
rect 3694 2320 3700 2372
rect 3752 2360 3758 2372
rect 4062 2360 4068 2372
rect 3752 2332 4068 2360
rect 3752 2320 3758 2332
rect 4062 2320 4068 2332
rect 4120 2320 4126 2372
rect 6380 2332 6486 2360
rect 4246 2252 4252 2304
rect 4304 2292 4310 2304
rect 6380 2292 6408 2332
rect 7466 2320 7472 2372
rect 7524 2360 7530 2372
rect 7576 2360 7604 2391
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8849 2431 8907 2437
rect 8849 2428 8861 2431
rect 7984 2400 8861 2428
rect 7984 2388 7990 2400
rect 8849 2397 8861 2400
rect 8895 2397 8907 2431
rect 9214 2428 9220 2440
rect 9175 2400 9220 2428
rect 8849 2391 8907 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9490 2428 9496 2440
rect 9451 2400 9496 2428
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 7524 2332 7604 2360
rect 7524 2320 7530 2332
rect 9306 2292 9312 2304
rect 4304 2264 6408 2292
rect 9267 2264 9312 2292
rect 4304 2252 4310 2264
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 3036 2202 9844 2224
rect 3036 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 5194 2202
rect 5246 2150 5258 2202
rect 5310 2150 5322 2202
rect 5374 2150 9844 2202
rect 3036 2128 9844 2150
rect 4062 2088 4068 2100
rect 4023 2060 4068 2088
rect 4062 2048 4068 2060
rect 4120 2048 4126 2100
rect 7926 2088 7932 2100
rect 4264 2060 5856 2088
rect 7887 2060 7932 2088
rect 3326 1912 3332 1964
rect 3384 1952 3390 1964
rect 4264 1961 4292 2060
rect 4525 2023 4583 2029
rect 4525 1989 4537 2023
rect 4571 2020 4583 2023
rect 4614 2020 4620 2032
rect 4571 1992 4620 2020
rect 4571 1989 4583 1992
rect 4525 1983 4583 1989
rect 4614 1980 4620 1992
rect 4672 1980 4678 2032
rect 4249 1955 4307 1961
rect 4249 1952 4261 1955
rect 3384 1924 4261 1952
rect 3384 1912 3390 1924
rect 4249 1921 4261 1924
rect 4295 1921 4307 1955
rect 5828 1952 5856 2060
rect 7926 2048 7932 2060
rect 7984 2048 7990 2100
rect 7190 1980 7196 2032
rect 7248 1980 7254 2032
rect 6178 1952 6184 1964
rect 4249 1915 4307 1921
rect 4062 1844 4068 1896
rect 4120 1884 4126 1896
rect 5644 1884 5672 1938
rect 5828 1924 6184 1952
rect 6178 1912 6184 1924
rect 6236 1912 6242 1964
rect 8297 1955 8355 1961
rect 8297 1921 8309 1955
rect 8343 1952 8355 1955
rect 8386 1952 8392 1964
rect 8343 1924 8392 1952
rect 8343 1921 8355 1924
rect 8297 1915 8355 1921
rect 8386 1912 8392 1924
rect 8444 1912 8450 1964
rect 5902 1884 5908 1896
rect 4120 1856 5908 1884
rect 4120 1844 4126 1856
rect 5902 1844 5908 1856
rect 5960 1844 5966 1896
rect 6086 1844 6092 1896
rect 6144 1884 6150 1896
rect 6454 1884 6460 1896
rect 6144 1856 6460 1884
rect 6144 1844 6150 1856
rect 6454 1844 6460 1856
rect 6512 1844 6518 1896
rect 8849 1887 8907 1893
rect 8849 1853 8861 1887
rect 8895 1884 8907 1887
rect 8941 1887 8999 1893
rect 8941 1884 8953 1887
rect 8895 1856 8953 1884
rect 8895 1853 8907 1856
rect 8849 1847 8907 1853
rect 8941 1853 8953 1856
rect 8987 1853 8999 1887
rect 8941 1847 8999 1853
rect 5997 1751 6055 1757
rect 5997 1717 6009 1751
rect 6043 1748 6055 1751
rect 6086 1748 6092 1760
rect 6043 1720 6092 1748
rect 6043 1717 6055 1720
rect 5997 1711 6055 1717
rect 6086 1708 6092 1720
rect 6144 1708 6150 1760
rect 9030 1708 9036 1760
rect 9088 1748 9094 1760
rect 9493 1751 9551 1757
rect 9493 1748 9505 1751
rect 9088 1720 9505 1748
rect 9088 1708 9094 1720
rect 9493 1717 9505 1720
rect 9539 1717 9551 1751
rect 9493 1711 9551 1717
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 4798 1504 4804 1556
rect 4856 1544 4862 1556
rect 5721 1547 5779 1553
rect 5721 1544 5733 1547
rect 4856 1516 5733 1544
rect 4856 1504 4862 1516
rect 5721 1513 5733 1516
rect 5767 1513 5779 1547
rect 5902 1544 5908 1556
rect 5863 1516 5908 1544
rect 5721 1507 5779 1513
rect 5902 1504 5908 1516
rect 5960 1504 5966 1556
rect 6454 1504 6460 1556
rect 6512 1544 6518 1556
rect 6733 1547 6791 1553
rect 6733 1544 6745 1547
rect 6512 1516 6745 1544
rect 6512 1504 6518 1516
rect 6733 1513 6745 1516
rect 6779 1513 6791 1547
rect 6733 1507 6791 1513
rect 7466 1504 7472 1556
rect 7524 1544 7530 1556
rect 7745 1547 7803 1553
rect 7745 1544 7757 1547
rect 7524 1516 7757 1544
rect 7524 1504 7530 1516
rect 7745 1513 7757 1516
rect 7791 1513 7803 1547
rect 7745 1507 7803 1513
rect 9214 1504 9220 1556
rect 9272 1544 9278 1556
rect 9309 1547 9367 1553
rect 9309 1544 9321 1547
rect 9272 1516 9321 1544
rect 9272 1504 9278 1516
rect 9309 1513 9321 1516
rect 9355 1513 9367 1547
rect 9309 1507 9367 1513
rect 7282 1436 7288 1488
rect 7340 1476 7346 1488
rect 7837 1479 7895 1485
rect 7837 1476 7849 1479
rect 7340 1448 7849 1476
rect 7340 1436 7346 1448
rect 7837 1445 7849 1448
rect 7883 1476 7895 1479
rect 8297 1479 8355 1485
rect 8297 1476 8309 1479
rect 7883 1448 8309 1476
rect 7883 1445 7895 1448
rect 7837 1439 7895 1445
rect 8297 1445 8309 1448
rect 8343 1476 8355 1479
rect 8481 1479 8539 1485
rect 8481 1476 8493 1479
rect 8343 1448 8493 1476
rect 8343 1445 8355 1448
rect 8297 1439 8355 1445
rect 8481 1445 8493 1448
rect 8527 1445 8539 1479
rect 8481 1439 8539 1445
rect 3326 1408 3332 1420
rect 3287 1380 3332 1408
rect 3326 1368 3332 1380
rect 3384 1368 3390 1420
rect 3605 1411 3663 1417
rect 3605 1377 3617 1411
rect 3651 1408 3663 1411
rect 3970 1408 3976 1420
rect 3651 1380 3976 1408
rect 3651 1377 3663 1380
rect 3605 1371 3663 1377
rect 3970 1368 3976 1380
rect 4028 1368 4034 1420
rect 9217 1411 9275 1417
rect 7404 1380 7604 1408
rect 4890 1300 4896 1352
rect 4948 1340 4954 1352
rect 5353 1343 5411 1349
rect 5353 1340 5365 1343
rect 4948 1312 5365 1340
rect 4948 1300 4954 1312
rect 5353 1309 5365 1312
rect 5399 1309 5411 1343
rect 5353 1303 5411 1309
rect 5442 1300 5448 1352
rect 5500 1340 5506 1352
rect 6086 1340 6092 1352
rect 5500 1312 5545 1340
rect 6047 1312 6092 1340
rect 5500 1300 5506 1312
rect 6086 1300 6092 1312
rect 6144 1300 6150 1352
rect 6730 1300 6736 1352
rect 6788 1340 6794 1352
rect 7404 1340 7432 1380
rect 7576 1349 7604 1380
rect 9217 1377 9229 1411
rect 9263 1408 9275 1411
rect 9306 1408 9312 1420
rect 9263 1380 9312 1408
rect 9263 1377 9275 1380
rect 9217 1371 9275 1377
rect 9306 1368 9312 1380
rect 9364 1408 9370 1420
rect 16574 1408 16580 1420
rect 9364 1380 16580 1408
rect 9364 1368 9370 1380
rect 16574 1368 16580 1380
rect 16632 1368 16638 1420
rect 6788 1312 7432 1340
rect 7469 1343 7527 1349
rect 6788 1300 6794 1312
rect 7469 1309 7481 1343
rect 7515 1309 7527 1343
rect 7469 1303 7527 1309
rect 7561 1343 7619 1349
rect 7561 1309 7573 1343
rect 7607 1309 7619 1343
rect 7561 1303 7619 1309
rect 4062 1232 4068 1284
rect 4120 1232 4126 1284
rect 5092 1244 7144 1272
rect 5092 1213 5120 1244
rect 5077 1207 5135 1213
rect 5077 1173 5089 1207
rect 5123 1173 5135 1207
rect 6822 1204 6828 1216
rect 6783 1176 6828 1204
rect 5077 1167 5135 1173
rect 6822 1164 6828 1176
rect 6880 1164 6886 1216
rect 7116 1204 7144 1244
rect 7484 1204 7512 1303
rect 8662 1300 8668 1352
rect 8720 1340 8726 1352
rect 8849 1343 8907 1349
rect 8849 1340 8861 1343
rect 8720 1312 8861 1340
rect 8720 1300 8726 1312
rect 8849 1309 8861 1312
rect 8895 1309 8907 1343
rect 9030 1340 9036 1352
rect 8991 1312 9036 1340
rect 8849 1303 8907 1309
rect 9030 1300 9036 1312
rect 9088 1300 9094 1352
rect 8113 1275 8171 1281
rect 8113 1241 8125 1275
rect 8159 1272 8171 1275
rect 8754 1272 8760 1284
rect 8159 1244 8760 1272
rect 8159 1241 8171 1244
rect 8113 1235 8171 1241
rect 8754 1232 8760 1244
rect 8812 1232 8818 1284
rect 7116 1176 7512 1204
rect 3036 1114 9844 1136
rect 3036 1062 5066 1114
rect 5118 1062 5130 1114
rect 5182 1062 5194 1114
rect 5246 1062 5258 1114
rect 5310 1062 5322 1114
rect 5374 1062 9844 1114
rect 3036 1040 9844 1062
rect 3602 960 3608 1012
rect 3660 1000 3666 1012
rect 6822 1000 6828 1012
rect 3660 972 6828 1000
rect 3660 960 3666 972
rect 6822 960 6828 972
rect 6880 960 6886 1012
<< via1 >>
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2136 11296 2188 11348
rect 2412 11296 2464 11348
rect 1860 11228 1912 11280
rect 3608 11228 3660 11280
rect 2412 11160 2464 11212
rect 1768 11092 1820 11144
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 1400 11024 1452 11076
rect 2320 11024 2372 11076
rect 4620 11296 4672 11348
rect 6184 11339 6236 11348
rect 6184 11305 6193 11339
rect 6193 11305 6227 11339
rect 6227 11305 6236 11339
rect 6184 11296 6236 11305
rect 4436 11271 4488 11280
rect 4436 11237 4445 11271
rect 4445 11237 4479 11271
rect 4479 11237 4488 11271
rect 4436 11228 4488 11237
rect 5080 11228 5132 11280
rect 6920 11228 6972 11280
rect 4528 11160 4580 11212
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 8024 11228 8076 11280
rect 8392 11228 8444 11280
rect 8116 11092 8168 11144
rect 4344 11024 4396 11076
rect 5080 11024 5132 11076
rect 2044 10999 2096 11008
rect 2044 10965 2053 10999
rect 2053 10965 2087 10999
rect 2087 10965 2096 10999
rect 2044 10956 2096 10965
rect 2596 10956 2648 11008
rect 3148 10956 3200 11008
rect 3516 10956 3568 11008
rect 3608 10999 3660 11008
rect 3608 10965 3617 10999
rect 3617 10965 3651 10999
rect 3651 10965 3660 10999
rect 3608 10956 3660 10965
rect 4896 10956 4948 11008
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 5724 11024 5776 11076
rect 6276 11024 6328 11076
rect 7012 11067 7064 11076
rect 7012 11033 7021 11067
rect 7021 11033 7055 11067
rect 7055 11033 7064 11067
rect 7012 11024 7064 11033
rect 7196 11024 7248 11076
rect 13820 11296 13872 11348
rect 8852 11067 8904 11076
rect 6092 10956 6144 11008
rect 7380 10956 7432 11008
rect 8852 11033 8861 11067
rect 8861 11033 8895 11067
rect 8895 11033 8904 11067
rect 8852 11024 8904 11033
rect 9036 11067 9088 11076
rect 9036 11033 9045 11067
rect 9045 11033 9079 11067
rect 9079 11033 9088 11067
rect 9036 11024 9088 11033
rect 8208 10999 8260 11008
rect 8208 10965 8217 10999
rect 8217 10965 8251 10999
rect 8251 10965 8260 10999
rect 8208 10956 8260 10965
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5194 10854 5246 10906
rect 5258 10854 5310 10906
rect 5322 10854 5374 10906
rect 1400 10795 1452 10804
rect 1400 10761 1409 10795
rect 1409 10761 1443 10795
rect 1443 10761 1452 10795
rect 1400 10752 1452 10761
rect 2136 10752 2188 10804
rect 6092 10752 6144 10804
rect 2596 10684 2648 10736
rect 5540 10684 5592 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2044 10616 2096 10668
rect 3516 10616 3568 10668
rect 4344 10616 4396 10668
rect 4988 10616 5040 10668
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 6368 10616 6420 10668
rect 7104 10616 7156 10668
rect 2136 10548 2188 10600
rect 4252 10548 4304 10600
rect 6828 10548 6880 10600
rect 7012 10548 7064 10600
rect 13912 10752 13964 10804
rect 13820 10684 13872 10736
rect 8208 10616 8260 10668
rect 8760 10591 8812 10600
rect 8760 10557 8769 10591
rect 8769 10557 8803 10591
rect 8803 10557 8812 10591
rect 8760 10548 8812 10557
rect 1768 10523 1820 10532
rect 1768 10489 1777 10523
rect 1777 10489 1811 10523
rect 1811 10489 1820 10523
rect 1768 10480 1820 10489
rect 5632 10480 5684 10532
rect 6736 10480 6788 10532
rect 6920 10480 6972 10532
rect 13728 10548 13780 10600
rect 4620 10412 4672 10464
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 7472 10412 7524 10464
rect 8484 10412 8536 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 2228 10208 2280 10260
rect 4160 10208 4212 10260
rect 4620 10208 4672 10260
rect 1584 10072 1636 10124
rect 6368 10208 6420 10260
rect 6736 10208 6788 10260
rect 8760 10208 8812 10260
rect 1308 10047 1360 10056
rect 1308 10013 1317 10047
rect 1317 10013 1351 10047
rect 1351 10013 1360 10047
rect 1308 10004 1360 10013
rect 2320 10004 2372 10056
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 6552 10004 6604 10056
rect 7380 10004 7432 10056
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 2964 9936 3016 9988
rect 6000 9979 6052 9988
rect 6000 9945 6009 9979
rect 6009 9945 6043 9979
rect 6043 9945 6052 9979
rect 6000 9936 6052 9945
rect 7472 9936 7524 9988
rect 13544 9936 13596 9988
rect 1860 9868 1912 9920
rect 2136 9868 2188 9920
rect 3792 9868 3844 9920
rect 7840 9868 7892 9920
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5194 9766 5246 9818
rect 5258 9766 5310 9818
rect 5322 9766 5374 9818
rect 1308 9707 1360 9716
rect 1308 9673 1317 9707
rect 1317 9673 1351 9707
rect 1351 9673 1360 9707
rect 1308 9664 1360 9673
rect 6092 9664 6144 9716
rect 2320 9596 2372 9648
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 4436 9596 4488 9648
rect 6184 9639 6236 9648
rect 6184 9605 6193 9639
rect 6193 9605 6227 9639
rect 6227 9605 6236 9639
rect 6184 9596 6236 9605
rect 7104 9664 7156 9716
rect 8024 9596 8076 9648
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 5448 9528 5500 9580
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 4068 9460 4120 9512
rect 1676 9324 1728 9376
rect 2320 9324 2372 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 4896 9392 4948 9444
rect 5908 9460 5960 9512
rect 6736 9460 6788 9512
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 8484 9528 8536 9580
rect 7012 9460 7064 9512
rect 7840 9460 7892 9512
rect 4436 9324 4488 9376
rect 8668 9324 8720 9376
rect 9588 9324 9640 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 3240 9120 3292 9172
rect 3516 9120 3568 9172
rect 4160 9163 4212 9172
rect 4160 9129 4169 9163
rect 4169 9129 4203 9163
rect 4203 9129 4212 9163
rect 4160 9120 4212 9129
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 6000 9120 6052 9172
rect 6184 9120 6236 9172
rect 7104 9120 7156 9172
rect 8208 9120 8260 9172
rect 4436 9052 4488 9104
rect 13728 9052 13780 9104
rect 1768 8984 1820 9036
rect 1308 8959 1360 8968
rect 1308 8925 1317 8959
rect 1317 8925 1351 8959
rect 1351 8925 1360 8959
rect 1308 8916 1360 8925
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 6092 8984 6144 9036
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 1768 8848 1820 8900
rect 2872 8848 2924 8900
rect 3240 8848 3292 8900
rect 4712 8916 4764 8968
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 7564 8916 7616 8968
rect 8760 8916 8812 8968
rect 9128 8916 9180 8968
rect 2228 8780 2280 8832
rect 3056 8780 3108 8832
rect 3608 8823 3660 8832
rect 3608 8789 3617 8823
rect 3617 8789 3651 8823
rect 3651 8789 3660 8823
rect 3608 8780 3660 8789
rect 3700 8780 3752 8832
rect 4344 8780 4396 8832
rect 5816 8848 5868 8900
rect 6552 8848 6604 8900
rect 7840 8848 7892 8900
rect 4988 8780 5040 8832
rect 5540 8780 5592 8832
rect 6184 8780 6236 8832
rect 6368 8780 6420 8832
rect 6828 8780 6880 8832
rect 8024 8780 8076 8832
rect 8392 8780 8444 8832
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5194 8678 5246 8730
rect 5258 8678 5310 8730
rect 5322 8678 5374 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 3056 8576 3108 8628
rect 3148 8576 3200 8628
rect 3700 8576 3752 8628
rect 3608 8508 3660 8560
rect 4252 8508 4304 8560
rect 4988 8576 5040 8628
rect 4896 8551 4948 8560
rect 4896 8517 4905 8551
rect 4905 8517 4939 8551
rect 4939 8517 4948 8551
rect 4896 8508 4948 8517
rect 5264 8508 5316 8560
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 3424 8440 3476 8492
rect 2872 8372 2924 8424
rect 4620 8440 4672 8492
rect 5448 8440 5500 8492
rect 6368 8576 6420 8628
rect 6920 8576 6972 8628
rect 7472 8576 7524 8628
rect 8484 8576 8536 8628
rect 9128 8619 9180 8628
rect 4804 8304 4856 8356
rect 5448 8304 5500 8356
rect 6000 8440 6052 8492
rect 6276 8440 6328 8492
rect 6644 8440 6696 8492
rect 7104 8440 7156 8492
rect 8760 8440 8812 8492
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 9404 8372 9456 8424
rect 6736 8304 6788 8356
rect 7380 8304 7432 8356
rect 13636 8304 13688 8356
rect 2412 8236 2464 8288
rect 4896 8236 4948 8288
rect 5172 8236 5224 8288
rect 7288 8236 7340 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 1492 8032 1544 8084
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 1860 7939 1912 7948
rect 1860 7905 1869 7939
rect 1869 7905 1903 7939
rect 1903 7905 1912 7939
rect 1860 7896 1912 7905
rect 2320 7896 2372 7948
rect 4252 8032 4304 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 5264 8032 5316 8084
rect 6092 8032 6144 8084
rect 6460 8032 6512 8084
rect 8024 8032 8076 8084
rect 9404 8075 9456 8084
rect 6000 7964 6052 8016
rect 7840 7964 7892 8016
rect 8116 8007 8168 8016
rect 8116 7973 8125 8007
rect 8125 7973 8159 8007
rect 8159 7973 8168 8007
rect 8116 7964 8168 7973
rect 1492 7871 1544 7880
rect 1492 7837 1501 7871
rect 1501 7837 1535 7871
rect 1535 7837 1544 7871
rect 1492 7828 1544 7837
rect 3148 7828 3200 7880
rect 5356 7896 5408 7948
rect 5724 7896 5776 7948
rect 6276 7896 6328 7948
rect 5632 7828 5684 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6000 7828 6052 7880
rect 4712 7760 4764 7812
rect 7472 7828 7524 7880
rect 8392 7828 8444 7880
rect 9404 8041 9413 8075
rect 9413 8041 9447 8075
rect 9447 8041 9456 8075
rect 9404 8032 9456 8041
rect 6920 7760 6972 7812
rect 8116 7760 8168 7812
rect 9404 7760 9456 7812
rect 3148 7692 3200 7744
rect 3884 7692 3936 7744
rect 5632 7692 5684 7744
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 6368 7735 6420 7744
rect 6368 7701 6377 7735
rect 6377 7701 6411 7735
rect 6411 7701 6420 7735
rect 6368 7692 6420 7701
rect 7012 7692 7064 7744
rect 7840 7692 7892 7744
rect 9312 7692 9364 7744
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 5194 7590 5246 7642
rect 5258 7590 5310 7642
rect 5322 7590 5374 7642
rect 1308 7531 1360 7540
rect 1308 7497 1317 7531
rect 1317 7497 1351 7531
rect 1351 7497 1360 7531
rect 1308 7488 1360 7497
rect 1492 7488 1544 7540
rect 2320 7420 2372 7472
rect 2780 7463 2832 7472
rect 2780 7429 2789 7463
rect 2789 7429 2823 7463
rect 2823 7429 2832 7463
rect 2780 7420 2832 7429
rect 4528 7488 4580 7540
rect 3148 7420 3200 7472
rect 4988 7420 5040 7472
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4896 7352 4948 7404
rect 5448 7352 5500 7404
rect 7196 7488 7248 7540
rect 7564 7488 7616 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 8300 7420 8352 7472
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 8208 7352 8260 7404
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 1492 7284 1544 7336
rect 4436 7284 4488 7336
rect 7288 7284 7340 7336
rect 7564 7284 7616 7336
rect 6368 7216 6420 7268
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 6092 7148 6144 7200
rect 8760 7216 8812 7268
rect 8852 7148 8904 7200
rect 8944 7191 8996 7200
rect 8944 7157 8961 7191
rect 8961 7157 8995 7191
rect 8995 7157 8996 7191
rect 8944 7148 8996 7157
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 2228 6944 2280 6996
rect 5908 6944 5960 6996
rect 6368 6944 6420 6996
rect 6920 6944 6972 6996
rect 8668 6944 8720 6996
rect 9496 6944 9548 6996
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 4068 6808 4120 6860
rect 3148 6740 3200 6792
rect 7380 6808 7432 6860
rect 13728 6808 13780 6860
rect 3056 6672 3108 6724
rect 7472 6672 7524 6724
rect 1492 6604 1544 6656
rect 3516 6604 3568 6656
rect 5908 6604 5960 6656
rect 6644 6604 6696 6656
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 9036 6672 9088 6724
rect 8392 6604 8444 6656
rect 9312 6604 9364 6656
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5194 6502 5246 6554
rect 5258 6502 5310 6554
rect 5322 6502 5374 6554
rect 1492 6443 1544 6452
rect 1492 6409 1501 6443
rect 1501 6409 1535 6443
rect 1535 6409 1544 6443
rect 1492 6400 1544 6409
rect 2964 6264 3016 6316
rect 5540 6400 5592 6452
rect 5724 6400 5776 6452
rect 6368 6400 6420 6452
rect 6644 6400 6696 6452
rect 4068 6332 4120 6384
rect 7932 6375 7984 6384
rect 7932 6341 7941 6375
rect 7941 6341 7975 6375
rect 7975 6341 7984 6375
rect 7932 6332 7984 6341
rect 8116 6332 8168 6384
rect 8300 6332 8352 6384
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 6092 6264 6144 6316
rect 7104 6264 7156 6316
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 3976 6196 4028 6248
rect 6184 6239 6236 6248
rect 6184 6205 6193 6239
rect 6193 6205 6227 6239
rect 6227 6205 6236 6239
rect 6184 6196 6236 6205
rect 8392 6264 8444 6316
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 8852 6264 8904 6316
rect 9864 6264 9916 6316
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 3056 6060 3108 6112
rect 3240 6103 3292 6112
rect 3240 6069 3249 6103
rect 3249 6069 3283 6103
rect 3283 6069 3292 6103
rect 3240 6060 3292 6069
rect 8208 6128 8260 6180
rect 8668 6128 8720 6180
rect 4068 6060 4120 6112
rect 9220 6060 9272 6112
rect 13452 6060 13504 6112
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 1676 5899 1728 5908
rect 1676 5865 1685 5899
rect 1685 5865 1719 5899
rect 1719 5865 1728 5899
rect 1676 5856 1728 5865
rect 2964 5856 3016 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 7288 5856 7340 5908
rect 8024 5856 8076 5908
rect 8576 5856 8628 5908
rect 3700 5831 3752 5840
rect 3700 5797 3709 5831
rect 3709 5797 3743 5831
rect 3743 5797 3752 5831
rect 3700 5788 3752 5797
rect 8668 5788 8720 5840
rect 8760 5788 8812 5840
rect 9312 5788 9364 5840
rect 9496 5831 9548 5840
rect 9496 5797 9505 5831
rect 9505 5797 9539 5831
rect 9539 5797 9548 5831
rect 9496 5788 9548 5797
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 3700 5652 3752 5704
rect 5816 5720 5868 5772
rect 6828 5720 6880 5772
rect 8300 5720 8352 5772
rect 13820 5720 13872 5772
rect 1492 5584 1544 5636
rect 3148 5627 3200 5636
rect 3148 5593 3157 5627
rect 3157 5593 3191 5627
rect 3191 5593 3200 5627
rect 3148 5584 3200 5593
rect 2780 5516 2832 5568
rect 7472 5584 7524 5636
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 9864 5652 9916 5704
rect 8300 5516 8352 5568
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5194 5414 5246 5466
rect 5258 5414 5310 5466
rect 5322 5414 5374 5466
rect 2412 5312 2464 5364
rect 4620 5312 4672 5364
rect 6460 5355 6512 5364
rect 3240 5244 3292 5296
rect 3056 5176 3108 5228
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 6552 5312 6604 5364
rect 8116 5312 8168 5364
rect 5540 5244 5592 5296
rect 6276 5244 6328 5296
rect 8760 5244 8812 5296
rect 5632 5176 5684 5228
rect 6092 5176 6144 5228
rect 6828 5176 6880 5228
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 8392 5176 8444 5228
rect 6184 5108 6236 5160
rect 6368 5108 6420 5160
rect 4160 5083 4212 5092
rect 4160 5049 4169 5083
rect 4169 5049 4203 5083
rect 4203 5049 4212 5083
rect 4160 5040 4212 5049
rect 8208 5040 8260 5092
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 4620 5015 4672 5024
rect 4620 4981 4629 5015
rect 4629 4981 4663 5015
rect 4663 4981 4672 5015
rect 4620 4972 4672 4981
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 8024 4972 8076 5024
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 9588 4972 9640 5024
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 4804 4768 4856 4820
rect 4988 4768 5040 4820
rect 7104 4768 7156 4820
rect 8392 4768 8444 4820
rect 13820 4768 13872 4820
rect 5724 4632 5776 4684
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 3608 4564 3660 4616
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4528 4564 4580 4616
rect 6092 4632 6144 4684
rect 7012 4632 7064 4684
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 8760 4632 8812 4684
rect 6460 4564 6512 4573
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 5448 4496 5500 4548
rect 4252 4428 4304 4480
rect 4344 4428 4396 4480
rect 6000 4496 6052 4548
rect 6276 4428 6328 4480
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 5194 4326 5246 4378
rect 5258 4326 5310 4378
rect 5322 4326 5374 4378
rect 3516 4224 3568 4276
rect 3700 4267 3752 4276
rect 3700 4233 3709 4267
rect 3709 4233 3743 4267
rect 3743 4233 3752 4267
rect 3700 4224 3752 4233
rect 7472 4224 7524 4276
rect 4160 4156 4212 4208
rect 4252 4156 4304 4208
rect 5356 4156 5408 4208
rect 6552 4156 6604 4208
rect 6092 4131 6144 4140
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 4344 4020 4396 4072
rect 4804 4020 4856 4072
rect 6460 4020 6512 4072
rect 4068 3884 4120 3936
rect 5540 3952 5592 4004
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 8392 4020 8444 4072
rect 8208 3952 8260 4004
rect 6000 3884 6052 3936
rect 6828 3884 6880 3936
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 4068 3680 4120 3732
rect 4344 3680 4396 3732
rect 6092 3680 6144 3732
rect 6276 3680 6328 3732
rect 9864 3680 9916 3732
rect 3424 3612 3476 3664
rect 4160 3544 4212 3596
rect 4896 3544 4948 3596
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 4804 3476 4856 3528
rect 7472 3544 7524 3596
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 5632 3476 5684 3528
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 6644 3476 6696 3485
rect 9312 3476 9364 3528
rect 9404 3476 9456 3528
rect 4620 3408 4672 3460
rect 5816 3408 5868 3460
rect 8300 3408 8352 3460
rect 3608 3340 3660 3392
rect 4252 3340 4304 3392
rect 4712 3383 4764 3392
rect 4712 3349 4721 3383
rect 4721 3349 4755 3383
rect 4755 3349 4764 3383
rect 4712 3340 4764 3349
rect 6920 3340 6972 3392
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5194 3238 5246 3290
rect 5258 3238 5310 3290
rect 5322 3238 5374 3290
rect 4436 3136 4488 3188
rect 4712 3136 4764 3188
rect 4344 3068 4396 3120
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 5540 3136 5592 3188
rect 5724 3136 5776 3188
rect 8300 3179 8352 3188
rect 8300 3145 8309 3179
rect 8309 3145 8343 3179
rect 8343 3145 8352 3179
rect 8300 3136 8352 3145
rect 9312 3136 9364 3188
rect 5908 3068 5960 3120
rect 7288 3068 7340 3120
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 6184 2932 6236 2984
rect 8392 2932 8444 2984
rect 8760 2975 8812 2984
rect 8760 2941 8769 2975
rect 8769 2941 8803 2975
rect 8803 2941 8812 2975
rect 8760 2932 8812 2941
rect 9220 2932 9272 2984
rect 9404 2975 9456 2984
rect 9404 2941 9413 2975
rect 9413 2941 9447 2975
rect 9447 2941 9456 2975
rect 9404 2932 9456 2941
rect 3608 2864 3660 2916
rect 4436 2796 4488 2848
rect 4712 2796 4764 2848
rect 6368 2796 6420 2848
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 5448 2592 5500 2644
rect 5632 2524 5684 2576
rect 9036 2592 9088 2644
rect 8208 2524 8260 2576
rect 3332 2499 3384 2508
rect 3332 2465 3341 2499
rect 3341 2465 3375 2499
rect 3375 2465 3384 2499
rect 3332 2456 3384 2465
rect 5448 2456 5500 2508
rect 8116 2456 8168 2508
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 6092 2431 6144 2440
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 3608 2363 3660 2372
rect 3608 2329 3617 2363
rect 3617 2329 3651 2363
rect 3651 2329 3660 2363
rect 3608 2320 3660 2329
rect 3700 2320 3752 2372
rect 4068 2320 4120 2372
rect 4252 2252 4304 2304
rect 7472 2320 7524 2372
rect 7932 2388 7984 2440
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 5194 2150 5246 2202
rect 5258 2150 5310 2202
rect 5322 2150 5374 2202
rect 4068 2091 4120 2100
rect 4068 2057 4077 2091
rect 4077 2057 4111 2091
rect 4111 2057 4120 2091
rect 4068 2048 4120 2057
rect 7932 2091 7984 2100
rect 3332 1912 3384 1964
rect 4620 1980 4672 2032
rect 7932 2057 7941 2091
rect 7941 2057 7975 2091
rect 7975 2057 7984 2091
rect 7932 2048 7984 2057
rect 7196 1980 7248 2032
rect 6184 1955 6236 1964
rect 4068 1844 4120 1896
rect 6184 1921 6193 1955
rect 6193 1921 6227 1955
rect 6227 1921 6236 1955
rect 6184 1912 6236 1921
rect 8392 1912 8444 1964
rect 5908 1844 5960 1896
rect 6092 1844 6144 1896
rect 6460 1887 6512 1896
rect 6460 1853 6469 1887
rect 6469 1853 6503 1887
rect 6503 1853 6512 1887
rect 6460 1844 6512 1853
rect 6092 1708 6144 1760
rect 9036 1708 9088 1760
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 4804 1504 4856 1556
rect 5908 1547 5960 1556
rect 5908 1513 5917 1547
rect 5917 1513 5951 1547
rect 5951 1513 5960 1547
rect 5908 1504 5960 1513
rect 6460 1504 6512 1556
rect 7472 1504 7524 1556
rect 9220 1504 9272 1556
rect 7288 1436 7340 1488
rect 3332 1411 3384 1420
rect 3332 1377 3341 1411
rect 3341 1377 3375 1411
rect 3375 1377 3384 1411
rect 3332 1368 3384 1377
rect 3976 1368 4028 1420
rect 4896 1300 4948 1352
rect 5448 1343 5500 1352
rect 5448 1309 5457 1343
rect 5457 1309 5491 1343
rect 5491 1309 5500 1343
rect 6092 1343 6144 1352
rect 5448 1300 5500 1309
rect 6092 1309 6101 1343
rect 6101 1309 6135 1343
rect 6135 1309 6144 1343
rect 6092 1300 6144 1309
rect 6736 1300 6788 1352
rect 9312 1368 9364 1420
rect 16580 1368 16632 1420
rect 4068 1232 4120 1284
rect 6828 1207 6880 1216
rect 6828 1173 6837 1207
rect 6837 1173 6871 1207
rect 6871 1173 6880 1207
rect 6828 1164 6880 1173
rect 8668 1300 8720 1352
rect 9036 1343 9088 1352
rect 9036 1309 9045 1343
rect 9045 1309 9079 1343
rect 9079 1309 9088 1343
rect 9036 1300 9088 1309
rect 8760 1232 8812 1284
rect 5066 1062 5118 1114
rect 5130 1062 5182 1114
rect 5194 1062 5246 1114
rect 5258 1062 5310 1114
rect 5322 1062 5374 1114
rect 3608 960 3660 1012
rect 6828 960 6880 1012
<< metal2 >>
rect 938 12322 994 13000
rect 1398 12322 1454 13000
rect 938 12294 1348 12322
rect 938 12200 994 12294
rect 1320 10962 1348 12294
rect 1398 12294 1532 12322
rect 1398 12200 1454 12294
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1412 10962 1440 11018
rect 1320 10934 1440 10962
rect 1412 10810 1440 10934
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1320 9722 1348 9998
rect 1308 9716 1360 9722
rect 1308 9658 1360 9664
rect 1308 8968 1360 8974
rect 1308 8910 1360 8916
rect 1320 7546 1348 8910
rect 1504 8090 1532 12294
rect 1858 12200 1914 13000
rect 2318 12322 2374 13000
rect 2778 12322 2834 13000
rect 2318 12294 2452 12322
rect 2318 12200 2374 12294
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10130 1624 10610
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1688 9382 1716 11290
rect 1872 11286 1900 12200
rect 2424 11354 2452 12294
rect 2778 12294 3096 12322
rect 2778 12200 2834 12294
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10538 1808 11086
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2056 10674 2084 10950
rect 2148 10810 2176 11290
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 1768 10532 1820 10538
rect 1768 10474 1820 10480
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1780 9042 1808 10474
rect 2148 9926 2176 10542
rect 2240 10266 2268 11086
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2332 10062 2360 11018
rect 2424 10146 2452 11154
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2608 10742 2636 10950
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2424 10118 2820 10146
rect 2320 10056 2372 10062
rect 2792 10033 2820 10118
rect 2320 9998 2372 10004
rect 2778 10024 2834 10033
rect 2778 9959 2834 9968
rect 2964 9988 3016 9994
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1780 8634 1808 8842
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1872 7954 1900 9862
rect 2792 9654 2820 9959
rect 2964 9930 3016 9936
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2332 9382 2360 9590
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8430 2268 8774
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1504 7546 1532 7822
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1492 7336 1544 7342
rect 1596 7324 1624 7890
rect 1544 7296 1624 7324
rect 1492 7278 1544 7284
rect 1504 6866 1532 7278
rect 2240 7002 2268 8366
rect 2332 7954 2360 9318
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2976 9058 3004 9930
rect 2884 9030 3004 9058
rect 2884 8906 2912 9030
rect 3068 8922 3096 12294
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 13818 12336 13874 12345
rect 13818 12271 13874 12280
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 9058 3188 10950
rect 3252 9738 3280 12200
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3620 11014 3648 11222
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3528 10674 3556 10950
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3620 10062 3648 10950
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3252 9710 3372 9738
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3252 9178 3280 9522
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3160 9030 3280 9058
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2976 8894 3188 8922
rect 3252 8906 3280 9030
rect 2976 8514 3004 8894
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8634 3096 8774
rect 3160 8634 3188 8894
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2884 8486 3004 8514
rect 2884 8430 2912 8486
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2332 7478 2360 7890
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6458 1532 6598
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1504 5914 1532 6394
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1688 5914 1716 6190
rect 2424 6118 2452 8230
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 3148 7880 3200 7886
rect 3068 7840 3148 7868
rect 2780 7472 2832 7478
rect 2778 7440 2780 7449
rect 2832 7440 2834 7449
rect 2778 7375 2834 7384
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 3068 6730 3096 7840
rect 3148 7822 3200 7828
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 7478 3188 7686
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2688 6248 2740 6254
rect 2686 6216 2688 6225
rect 2740 6216 2742 6225
rect 2686 6151 2742 6160
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1504 5642 1532 5850
rect 1492 5636 1544 5642
rect 1492 5578 1544 5584
rect 2424 5370 2452 6054
rect 2566 6012 2874 6032
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5936 2874 5956
rect 2976 5914 3004 6258
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2792 3505 2820 5510
rect 3068 5234 3096 6054
rect 3160 5642 3188 6734
rect 3252 6202 3280 8842
rect 3344 7290 3372 9710
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 8498 3464 9318
rect 3528 9178 3556 9454
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3712 8838 3740 12200
rect 4172 10418 4200 12200
rect 4632 11354 4660 12200
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 5092 11286 5120 12200
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10606 4292 11086
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4356 10674 4384 11018
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4172 10390 4292 10418
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 8974 3832 9862
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3620 8566 3648 8774
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3344 7262 3648 7290
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 6322 3372 7142
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3252 6174 3372 6202
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3252 5302 3280 6054
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3344 4826 3372 6174
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3436 3670 3464 5646
rect 3528 4622 3556 6598
rect 3620 4622 3648 7262
rect 3712 5846 3740 8570
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7449 3924 7686
rect 3882 7440 3938 7449
rect 3882 7375 3884 7384
rect 3936 7375 3938 7384
rect 3884 7346 3936 7352
rect 3896 7315 3924 7346
rect 4080 6866 4108 9454
rect 4172 9178 4200 10202
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4264 8566 4292 10390
rect 4448 9654 4476 11222
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4448 9110 4476 9318
rect 4540 9178 4568 11154
rect 5092 11082 5120 11222
rect 5080 11076 5132 11082
rect 5000 11036 5080 11064
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10266 4660 10406
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4908 9450 4936 10950
rect 5000 10674 5028 11036
rect 5552 11064 5580 12200
rect 5724 11076 5776 11082
rect 5552 11036 5724 11064
rect 5080 11018 5132 11024
rect 5724 11018 5776 11024
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5066 10908 5374 10928
rect 5066 10906 5072 10908
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5368 10906 5374 10908
rect 5128 10854 5130 10906
rect 5310 10854 5312 10906
rect 5066 10852 5072 10854
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5368 10852 5374 10854
rect 5066 10832 5374 10852
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5066 9820 5374 9840
rect 5066 9818 5072 9820
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5368 9818 5374 9820
rect 5128 9766 5130 9818
rect 5310 9766 5312 9818
rect 5066 9764 5072 9766
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5368 9764 5374 9766
rect 5066 9744 5374 9764
rect 5460 9586 5488 10950
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4436 9104 4488 9110
rect 4436 9046 4488 9052
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3712 5710 3740 5782
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3988 5030 4016 6190
rect 4080 6118 4108 6326
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4264 5914 4292 8026
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3528 4282 3556 4558
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3620 3738 3648 4558
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 2778 3496 2834 3505
rect 2778 3431 2834 3440
rect 3436 2774 3464 3606
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 3058 3648 3334
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3344 2746 3464 2774
rect 3344 2514 3372 2746
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3344 1970 3372 2450
rect 3620 2378 3648 2858
rect 3712 2378 3740 4218
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 3344 1426 3372 1906
rect 3332 1420 3384 1426
rect 3332 1362 3384 1368
rect 3620 1018 3648 2314
rect 3988 1426 4016 4966
rect 4172 4214 4200 5034
rect 4356 4622 4384 8774
rect 4448 7342 4476 9046
rect 4540 7546 4568 9114
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4632 5370 4660 8434
rect 4724 7818 4752 8910
rect 4908 8566 4936 9386
rect 5552 8974 5580 10678
rect 5632 10532 5684 10538
rect 5632 10474 5684 10480
rect 5080 8968 5132 8974
rect 5078 8936 5080 8945
rect 5540 8968 5592 8974
rect 5132 8936 5134 8945
rect 5540 8910 5592 8916
rect 5078 8871 5134 8880
rect 5552 8838 5580 8910
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5000 8634 5028 8774
rect 5066 8732 5374 8752
rect 5066 8730 5072 8732
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5368 8730 5374 8732
rect 5128 8678 5130 8730
rect 5310 8678 5312 8730
rect 5066 8676 5072 8678
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5368 8676 5374 8678
rect 5066 8656 5374 8676
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5446 8528 5502 8537
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4816 5137 4844 8298
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 4908 7410 4936 8230
rect 5184 8090 5212 8230
rect 5276 8090 5304 8502
rect 5368 8472 5446 8480
rect 5368 8452 5448 8472
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5368 7954 5396 8452
rect 5500 8463 5502 8472
rect 5448 8434 5500 8440
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5066 7644 5374 7664
rect 5066 7642 5072 7644
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5368 7642 5374 7644
rect 5128 7590 5130 7642
rect 5310 7590 5312 7642
rect 5066 7588 5072 7590
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5368 7588 5374 7590
rect 5066 7568 5374 7588
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4802 5128 4858 5137
rect 4802 5063 4858 5072
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4356 4486 4384 4558
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4264 4214 4292 4422
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4356 4162 4384 4422
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3738 4108 3878
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4172 3602 4200 4150
rect 4356 4134 4476 4162
rect 4344 4072 4396 4078
rect 4264 4020 4344 4026
rect 4264 4014 4396 4020
rect 4264 3998 4384 4014
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4264 3534 4292 3998
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4080 2106 4108 2314
rect 4264 2310 4292 3334
rect 4356 3126 4384 3674
rect 4448 3194 4476 4134
rect 4540 3534 4568 4558
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4632 3466 4660 4966
rect 4816 4826 4844 4966
rect 5000 4826 5028 7414
rect 5460 7410 5488 8298
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5066 6556 5374 6576
rect 5066 6554 5072 6556
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5368 6554 5374 6556
rect 5128 6502 5130 6554
rect 5310 6502 5312 6554
rect 5066 6500 5072 6502
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5368 6500 5374 6502
rect 5066 6480 5374 6500
rect 5552 6458 5580 8774
rect 5644 7886 5672 10474
rect 6012 10146 6040 12200
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6104 10810 6132 10950
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6196 10674 6224 11290
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 5920 10118 6040 10146
rect 5920 9518 5948 10118
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 6012 9178 6040 9930
rect 6104 9722 6132 9998
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6196 9654 6224 10610
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6196 9042 6224 9114
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5632 7880 5684 7886
rect 5630 7848 5632 7857
rect 5684 7848 5686 7857
rect 5630 7783 5686 7792
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5066 5468 5374 5488
rect 5066 5466 5072 5468
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5368 5466 5374 5468
rect 5128 5414 5130 5466
rect 5310 5414 5312 5466
rect 5066 5412 5072 5414
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5368 5412 5374 5414
rect 5066 5392 5374 5412
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5552 4570 5580 5238
rect 5644 5234 5672 7686
rect 5736 6458 5764 7890
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5828 5778 5856 8842
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 8022 6040 8434
rect 6104 8090 6132 8978
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6000 8016 6052 8022
rect 5920 7964 6000 7970
rect 5920 7958 6052 7964
rect 5920 7942 6040 7958
rect 5920 7886 5948 7942
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5920 7002 5948 7822
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5908 6656 5960 6662
rect 6012 6644 6040 7822
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 7313 6132 7686
rect 6090 7304 6146 7313
rect 6090 7239 6146 7248
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 5960 6616 6040 6644
rect 5908 6598 5960 6604
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5460 4554 5580 4570
rect 5448 4548 5580 4554
rect 5500 4542 5580 4548
rect 5448 4490 5500 4496
rect 5066 4380 5374 4400
rect 5066 4378 5072 4380
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5368 4378 5374 4380
rect 5128 4326 5130 4378
rect 5310 4326 5312 4378
rect 5066 4324 5072 4326
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5368 4324 5374 4326
rect 5066 4304 5374 4324
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4816 3534 4844 4014
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3194 4752 3334
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4448 2854 4476 3130
rect 4816 3074 4844 3470
rect 4632 3046 4844 3074
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4080 1902 4108 2042
rect 4632 2038 4660 3046
rect 4712 2848 4764 2854
rect 4764 2796 4844 2802
rect 4712 2790 4844 2796
rect 4724 2774 4844 2790
rect 4620 2032 4672 2038
rect 4620 1974 4672 1980
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 4080 1290 4108 1838
rect 4816 1562 4844 2774
rect 4804 1556 4856 1562
rect 4804 1498 4856 1504
rect 4908 1358 4936 3538
rect 5368 3482 5396 4150
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5552 3534 5580 3946
rect 5540 3528 5592 3534
rect 5368 3454 5488 3482
rect 5540 3470 5592 3476
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5066 3292 5374 3312
rect 5066 3290 5072 3292
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5368 3290 5374 3292
rect 5128 3238 5130 3290
rect 5310 3238 5312 3290
rect 5066 3236 5072 3238
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5368 3236 5374 3238
rect 5066 3216 5374 3236
rect 5460 2650 5488 3454
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5066 2204 5374 2224
rect 5066 2202 5072 2204
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5368 2202 5374 2204
rect 5128 2150 5130 2202
rect 5310 2150 5312 2202
rect 5066 2148 5072 2150
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5368 2148 5374 2150
rect 5066 2128 5374 2148
rect 5460 1358 5488 2450
rect 5552 2446 5580 3130
rect 5644 2582 5672 3470
rect 5736 3194 5764 4626
rect 5828 3466 5856 5714
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5920 3126 5948 6598
rect 6104 6322 6132 7142
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6196 6254 6224 8774
rect 6288 8498 6316 11018
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6380 10266 6408 10610
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6472 9674 6500 12200
rect 13726 11928 13782 11937
rect 13726 11863 13782 11872
rect 13450 11520 13506 11529
rect 7566 11452 7874 11472
rect 13450 11455 13506 11464
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11376 7874 11396
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 6932 10690 6960 11222
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7024 10713 7052 11018
rect 6840 10662 6960 10690
rect 7010 10704 7066 10713
rect 6840 10606 6868 10662
rect 7010 10639 7066 10648
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6380 9646 6500 9674
rect 6380 8838 6408 9646
rect 6564 8906 6592 9998
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6288 7954 6316 8434
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6380 7834 6408 8570
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6288 7806 6408 7834
rect 6288 7750 6316 7806
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6104 4690 6132 5170
rect 6196 5166 6224 6190
rect 6288 5794 6316 7686
rect 6380 7274 6408 7686
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6380 6458 6408 6938
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6288 5766 6408 5794
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6012 3942 6040 4490
rect 6288 4486 6316 5238
rect 6380 5166 6408 5766
rect 6472 5370 6500 8026
rect 6564 5370 6592 8842
rect 6656 8498 6684 10406
rect 6748 10266 6776 10474
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6932 9586 6960 10474
rect 7024 10470 7052 10542
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7024 9518 7052 10406
rect 7116 9722 7144 10610
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6748 8922 6776 9454
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6748 8894 7052 8922
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6642 7848 6698 7857
rect 6642 7783 6698 7792
rect 6656 6662 6684 7783
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6472 4706 6500 5306
rect 6472 4678 6592 4706
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6104 3738 6132 4082
rect 6288 3738 6316 4422
rect 6472 4078 6500 4558
rect 6564 4214 6592 4678
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6656 3534 6684 6394
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6104 1902 6132 2382
rect 6196 1970 6224 2926
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6380 2417 6408 2790
rect 6366 2408 6422 2417
rect 6366 2343 6422 2352
rect 6184 1964 6236 1970
rect 6184 1906 6236 1912
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 6092 1896 6144 1902
rect 6092 1838 6144 1844
rect 6460 1896 6512 1902
rect 6460 1838 6512 1844
rect 5920 1562 5948 1838
rect 6092 1760 6144 1766
rect 6092 1702 6144 1708
rect 5908 1556 5960 1562
rect 5908 1498 5960 1504
rect 6104 1358 6132 1702
rect 6472 1562 6500 1838
rect 6460 1556 6512 1562
rect 6460 1498 6512 1504
rect 6748 1358 6776 8298
rect 6840 6225 6868 8774
rect 6918 8664 6974 8673
rect 6918 8599 6920 8608
rect 6972 8599 6974 8608
rect 6920 8570 6972 8576
rect 7024 7834 7052 8894
rect 7116 8498 7144 9114
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6920 7812 6972 7818
rect 7024 7806 7144 7834
rect 6920 7754 6972 7760
rect 6932 7410 6960 7754
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6932 7002 6960 7346
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6826 6216 6882 6225
rect 6826 6151 6882 6160
rect 6840 5778 6868 6151
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6840 5234 6868 5714
rect 6828 5228 6880 5234
rect 6880 5188 6960 5216
rect 6828 5170 6880 5176
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3369 6868 3878
rect 6932 3398 6960 5188
rect 7024 4690 7052 7686
rect 7116 6322 7144 7806
rect 7208 7546 7236 11018
rect 7380 11008 7432 11014
rect 7300 10968 7380 10996
rect 7300 8673 7328 10968
rect 7380 10950 7432 10956
rect 7930 10704 7986 10713
rect 7930 10639 7986 10648
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7392 10062 7420 10406
rect 7484 10146 7512 10406
rect 7566 10364 7874 10384
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10288 7874 10308
rect 7484 10118 7696 10146
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7378 9480 7434 9489
rect 7378 9415 7434 9424
rect 7286 8664 7342 8673
rect 7286 8599 7342 8608
rect 7392 8514 7420 9415
rect 7484 8634 7512 9930
rect 7668 9489 7696 10118
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9518 7880 9862
rect 7840 9512 7892 9518
rect 7654 9480 7710 9489
rect 7840 9454 7892 9460
rect 7654 9415 7710 9424
rect 7566 9276 7874 9296
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9200 7874 9220
rect 7564 8968 7616 8974
rect 7562 8936 7564 8945
rect 7616 8936 7618 8945
rect 7562 8871 7618 8880
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7852 8537 7880 8842
rect 7838 8528 7894 8537
rect 7392 8486 7512 8514
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7300 7342 7328 8230
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7116 4826 7144 6258
rect 7300 5914 7328 7278
rect 7392 6866 7420 8298
rect 7484 7886 7512 8486
rect 7838 8463 7894 8472
rect 7566 8188 7874 8208
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8112 7874 8132
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7852 7750 7880 7958
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7470 7440 7526 7449
rect 7470 7375 7526 7384
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7484 6730 7512 7375
rect 7576 7342 7604 7482
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7566 7100 7874 7120
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7024 7874 7044
rect 7472 6724 7524 6730
rect 7392 6684 7472 6712
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6920 3392 6972 3398
rect 6826 3360 6882 3369
rect 6920 3334 6972 3340
rect 6826 3295 6882 3304
rect 7288 3120 7340 3126
rect 7392 3108 7420 6684
rect 7472 6666 7524 6672
rect 7944 6390 7972 10639
rect 8036 9654 8064 11222
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8090 8064 8774
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8128 8022 8156 11086
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10826 8248 10950
rect 8220 10798 8340 10826
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8220 9178 8248 10610
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8312 9058 8340 10798
rect 8220 9030 8340 9058
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8128 6390 8156 7754
rect 8220 7410 8248 9030
rect 8404 8922 8432 11222
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8496 9586 8524 10406
rect 8772 10266 8800 10542
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8864 9874 8892 11018
rect 8772 9846 8892 9874
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8312 8894 8432 8922
rect 8312 7478 8340 8894
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 7886 8432 8774
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8312 6390 8340 6734
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 7566 6012 7874 6032
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5936 7874 5956
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7484 4282 7512 5578
rect 8036 5030 8064 5850
rect 8128 5370 8156 6326
rect 8404 6322 8432 6598
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8220 5409 8248 6122
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8312 5574 8340 5714
rect 8496 5658 8524 8570
rect 8680 7002 8708 9318
rect 8772 8974 8800 9846
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 8498 8800 8910
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8772 8265 8800 8434
rect 8758 8256 8814 8265
rect 8758 8191 8814 8200
rect 8772 7449 8800 8191
rect 8758 7440 8814 7449
rect 8758 7375 8814 7384
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8772 6798 8800 7210
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8588 5914 8616 6734
rect 8864 6322 8892 7142
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8680 5846 8708 6122
rect 8772 5846 8800 6258
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8496 5630 8708 5658
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8206 5400 8262 5409
rect 8116 5364 8168 5370
rect 8206 5335 8262 5344
rect 8116 5306 8168 5312
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7566 4924 7874 4944
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4848 7874 4868
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3602 7512 3878
rect 7566 3836 7874 3856
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3760 7874 3780
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7340 3080 7420 3108
rect 7288 3062 7340 3068
rect 7196 2032 7248 2038
rect 7300 2020 7328 3062
rect 7566 2748 7874 2768
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2672 7874 2692
rect 8128 2514 8156 5170
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8220 4010 8248 5034
rect 8404 4826 8432 5170
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8312 3194 8340 3402
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8404 2990 8432 4014
rect 8496 3058 8524 5510
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8392 2984 8444 2990
rect 8206 2952 8262 2961
rect 8392 2926 8444 2932
rect 8206 2887 8262 2896
rect 8220 2582 8248 2887
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7248 1992 7328 2020
rect 7196 1974 7248 1980
rect 7300 1494 7328 1992
rect 7484 1562 7512 2314
rect 7944 2106 7972 2382
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8404 1970 8432 2926
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 7566 1660 7874 1680
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1584 7874 1604
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 7288 1488 7340 1494
rect 7288 1430 7340 1436
rect 8680 1358 8708 5630
rect 8772 5302 8800 5782
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8772 4690 8800 4966
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8956 3777 8984 7142
rect 9048 6730 9076 11018
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9140 8634 9168 8910
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9416 8430 9444 9998
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9416 8090 9444 8366
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9600 7857 9628 9318
rect 9586 7848 9642 7857
rect 9404 7812 9456 7818
rect 9586 7783 9642 7792
rect 9404 7754 9456 7760
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7410 9352 7686
rect 9416 7546 9444 7754
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9312 6656 9364 6662
rect 9364 6616 9444 6644
rect 9312 6598 9364 6604
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8942 3768 8998 3777
rect 8942 3703 8998 3712
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 4896 1352 4948 1358
rect 4896 1294 4948 1300
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 6092 1352 6144 1358
rect 6092 1294 6144 1300
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 8772 1290 8800 2926
rect 9048 2650 9076 5646
rect 9232 4622 9260 6054
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9324 4298 9352 5782
rect 9232 4270 9352 4298
rect 9232 4146 9260 4270
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9232 2990 9260 4082
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3534 9352 3878
rect 9416 3534 9444 6616
rect 9508 6225 9536 6938
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9494 6216 9550 6225
rect 9494 6151 9550 6160
rect 9496 5840 9548 5846
rect 9494 5808 9496 5817
rect 9548 5808 9550 5817
rect 9494 5743 9550 5752
rect 9876 5710 9904 6258
rect 13464 6118 13492 11455
rect 13740 10606 13768 11863
rect 13832 11354 13860 12271
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13818 11112 13874 11121
rect 13818 11047 13874 11056
rect 13832 10742 13860 11047
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13634 10296 13690 10305
rect 13634 10231 13690 10240
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13556 7449 13584 9930
rect 13648 8362 13676 10231
rect 13818 9480 13874 9489
rect 13924 9466 13952 10746
rect 13874 9438 13952 9466
rect 13818 9415 13874 9424
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13818 9072 13874 9081
rect 13740 8673 13768 9046
rect 13818 9007 13874 9016
rect 13726 8664 13782 8673
rect 13726 8599 13782 8608
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13542 7440 13598 7449
rect 13542 7375 13598 7384
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13740 6633 13768 6802
rect 13726 6624 13782 6633
rect 13726 6559 13782 6568
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13832 5778 13860 9007
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3194 9352 3334
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9232 2145 9260 2382
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9218 2136 9274 2145
rect 9218 2071 9274 2080
rect 9036 1760 9088 1766
rect 9036 1702 9088 1708
rect 9048 1358 9076 1702
rect 9232 1562 9260 2071
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 9324 1426 9352 2246
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 4068 1284 4120 1290
rect 4068 1226 4120 1232
rect 8760 1284 8812 1290
rect 8760 1226 8812 1232
rect 6828 1216 6880 1222
rect 6828 1158 6880 1164
rect 5066 1116 5374 1136
rect 5066 1114 5072 1116
rect 5128 1114 5152 1116
rect 5208 1114 5232 1116
rect 5288 1114 5312 1116
rect 5368 1114 5374 1116
rect 5128 1062 5130 1114
rect 5310 1062 5312 1114
rect 5066 1060 5072 1062
rect 5128 1060 5152 1062
rect 5208 1060 5232 1062
rect 5288 1060 5312 1062
rect 5368 1060 5374 1062
rect 5066 1040 5374 1060
rect 6840 1018 6868 1158
rect 3608 1012 3660 1018
rect 3608 954 3660 960
rect 6828 1012 6880 1018
rect 6828 954 6880 960
rect 9416 921 9444 2926
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9402 912 9458 921
rect 9402 847 9458 856
rect 9508 513 9536 2382
rect 9600 1737 9628 4966
rect 9876 4593 9904 5646
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 9862 4584 9918 4593
rect 9862 4519 9918 4528
rect 9876 3738 9904 4519
rect 13832 4185 13860 4762
rect 13818 4176 13874 4185
rect 13818 4111 13874 4120
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 16580 1420 16632 1426
rect 16580 1362 16632 1368
rect 16592 1329 16620 1362
rect 16578 1320 16634 1329
rect 16578 1255 16634 1264
rect 9494 504 9550 513
rect 9494 439 9550 448
<< via2 >>
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2778 9968 2834 10024
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 13818 12280 13874 12336
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2778 7420 2780 7440
rect 2780 7420 2832 7440
rect 2832 7420 2834 7440
rect 2778 7384 2834 7420
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2686 6196 2688 6216
rect 2688 6196 2740 6216
rect 2740 6196 2742 6216
rect 2686 6160 2742 6196
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 3882 7404 3938 7440
rect 3882 7384 3884 7404
rect 3884 7384 3936 7404
rect 3936 7384 3938 7404
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5118 10906
rect 5118 10854 5128 10906
rect 5152 10854 5182 10906
rect 5182 10854 5194 10906
rect 5194 10854 5208 10906
rect 5232 10854 5246 10906
rect 5246 10854 5258 10906
rect 5258 10854 5288 10906
rect 5312 10854 5322 10906
rect 5322 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5118 9818
rect 5118 9766 5128 9818
rect 5152 9766 5182 9818
rect 5182 9766 5194 9818
rect 5194 9766 5208 9818
rect 5232 9766 5246 9818
rect 5246 9766 5258 9818
rect 5258 9766 5288 9818
rect 5312 9766 5322 9818
rect 5322 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 2778 3440 2834 3496
rect 5078 8916 5080 8936
rect 5080 8916 5132 8936
rect 5132 8916 5134 8936
rect 5078 8880 5134 8916
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5118 8730
rect 5118 8678 5128 8730
rect 5152 8678 5182 8730
rect 5182 8678 5194 8730
rect 5194 8678 5208 8730
rect 5232 8678 5246 8730
rect 5246 8678 5258 8730
rect 5258 8678 5288 8730
rect 5312 8678 5322 8730
rect 5322 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 5446 8492 5502 8528
rect 5446 8472 5448 8492
rect 5448 8472 5500 8492
rect 5500 8472 5502 8492
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5118 7642
rect 5118 7590 5128 7642
rect 5152 7590 5182 7642
rect 5182 7590 5194 7642
rect 5194 7590 5208 7642
rect 5232 7590 5246 7642
rect 5246 7590 5258 7642
rect 5258 7590 5288 7642
rect 5312 7590 5322 7642
rect 5322 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 4802 5072 4858 5128
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5118 6554
rect 5118 6502 5128 6554
rect 5152 6502 5182 6554
rect 5182 6502 5194 6554
rect 5194 6502 5208 6554
rect 5232 6502 5246 6554
rect 5246 6502 5258 6554
rect 5258 6502 5288 6554
rect 5312 6502 5322 6554
rect 5322 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5630 7828 5632 7848
rect 5632 7828 5684 7848
rect 5684 7828 5686 7848
rect 5630 7792 5686 7828
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5118 5466
rect 5118 5414 5128 5466
rect 5152 5414 5182 5466
rect 5182 5414 5194 5466
rect 5194 5414 5208 5466
rect 5232 5414 5246 5466
rect 5246 5414 5258 5466
rect 5258 5414 5288 5466
rect 5312 5414 5322 5466
rect 5322 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 6090 7248 6146 7304
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5118 4378
rect 5118 4326 5128 4378
rect 5152 4326 5182 4378
rect 5182 4326 5194 4378
rect 5194 4326 5208 4378
rect 5232 4326 5246 4378
rect 5246 4326 5258 4378
rect 5258 4326 5288 4378
rect 5312 4326 5322 4378
rect 5322 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5118 3290
rect 5118 3238 5128 3290
rect 5152 3238 5182 3290
rect 5182 3238 5194 3290
rect 5194 3238 5208 3290
rect 5232 3238 5246 3290
rect 5246 3238 5258 3290
rect 5258 3238 5288 3290
rect 5312 3238 5322 3290
rect 5322 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5118 2202
rect 5118 2150 5128 2202
rect 5152 2150 5182 2202
rect 5182 2150 5194 2202
rect 5194 2150 5208 2202
rect 5232 2150 5246 2202
rect 5246 2150 5258 2202
rect 5258 2150 5288 2202
rect 5312 2150 5322 2202
rect 5322 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 13726 11872 13782 11928
rect 13450 11464 13506 11520
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 7010 10648 7066 10704
rect 6642 7792 6698 7848
rect 6366 2352 6422 2408
rect 6918 8628 6974 8664
rect 6918 8608 6920 8628
rect 6920 8608 6972 8628
rect 6972 8608 6974 8628
rect 6826 6160 6882 6216
rect 7930 10648 7986 10704
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 7378 9424 7434 9480
rect 7286 8608 7342 8664
rect 7654 9424 7710 9480
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 7562 8916 7564 8936
rect 7564 8916 7616 8936
rect 7616 8916 7618 8936
rect 7562 8880 7618 8916
rect 7838 8472 7894 8528
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 7470 7384 7526 7440
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 6826 3304 6882 3360
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 8758 8200 8814 8256
rect 8758 7384 8814 7440
rect 8206 5344 8262 5400
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 8206 2896 8262 2952
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 9586 7792 9642 7848
rect 8942 3712 8998 3768
rect 9494 6160 9550 6216
rect 9494 5788 9496 5808
rect 9496 5788 9548 5808
rect 9548 5788 9550 5808
rect 9494 5752 9550 5788
rect 13818 11056 13874 11112
rect 13634 10240 13690 10296
rect 13818 9424 13874 9480
rect 13818 9016 13874 9072
rect 13726 8608 13782 8664
rect 13542 7384 13598 7440
rect 13726 6568 13782 6624
rect 9218 2080 9274 2136
rect 5072 1114 5128 1116
rect 5152 1114 5208 1116
rect 5232 1114 5288 1116
rect 5312 1114 5368 1116
rect 5072 1062 5118 1114
rect 5118 1062 5128 1114
rect 5152 1062 5182 1114
rect 5182 1062 5194 1114
rect 5194 1062 5208 1114
rect 5232 1062 5246 1114
rect 5246 1062 5258 1114
rect 5258 1062 5288 1114
rect 5312 1062 5322 1114
rect 5322 1062 5368 1114
rect 5072 1060 5128 1062
rect 5152 1060 5208 1062
rect 5232 1060 5288 1062
rect 5312 1060 5368 1062
rect 9402 856 9458 912
rect 9862 4528 9918 4584
rect 13818 4120 13874 4176
rect 9586 1672 9642 1728
rect 16578 1264 16634 1320
rect 9494 448 9550 504
<< metal3 >>
rect 13813 12338 13879 12341
rect 14000 12338 34000 12368
rect 13813 12336 34000 12338
rect 13813 12280 13818 12336
rect 13874 12280 34000 12336
rect 13813 12278 34000 12280
rect 13813 12275 13879 12278
rect 14000 12248 34000 12278
rect 13721 11930 13787 11933
rect 14000 11930 34000 11960
rect 13721 11928 34000 11930
rect 13721 11872 13726 11928
rect 13782 11872 34000 11928
rect 13721 11870 34000 11872
rect 13721 11867 13787 11870
rect 14000 11840 34000 11870
rect 13445 11522 13511 11525
rect 14000 11522 34000 11552
rect 13445 11520 34000 11522
rect 13445 11464 13450 11520
rect 13506 11464 34000 11520
rect 13445 11462 34000 11464
rect 13445 11459 13511 11462
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 7560 11456 7880 11457
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 14000 11432 34000 11462
rect 7560 11391 7880 11392
rect 13813 11114 13879 11117
rect 14000 11114 34000 11144
rect 13813 11112 34000 11114
rect 13813 11056 13818 11112
rect 13874 11056 34000 11112
rect 13813 11054 34000 11056
rect 13813 11051 13879 11054
rect 14000 11024 34000 11054
rect 5060 10912 5380 10913
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 10847 5380 10848
rect 7005 10706 7071 10709
rect 7925 10706 7991 10709
rect 14000 10706 34000 10736
rect 7005 10704 34000 10706
rect 7005 10648 7010 10704
rect 7066 10648 7930 10704
rect 7986 10648 34000 10704
rect 7005 10646 34000 10648
rect 7005 10643 7071 10646
rect 7925 10643 7991 10646
rect 14000 10616 34000 10646
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 7560 10368 7880 10369
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 10303 7880 10304
rect 13629 10298 13695 10301
rect 14000 10298 34000 10328
rect 13629 10296 34000 10298
rect 13629 10240 13634 10296
rect 13690 10240 34000 10296
rect 13629 10238 34000 10240
rect 13629 10235 13695 10238
rect 14000 10208 34000 10238
rect 2773 10026 2839 10029
rect 2773 10024 12450 10026
rect 2773 9968 2778 10024
rect 2834 9968 12450 10024
rect 2773 9966 12450 9968
rect 2773 9963 2839 9966
rect 12390 9890 12450 9966
rect 14000 9890 34000 9920
rect 12390 9830 34000 9890
rect 5060 9824 5380 9825
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 14000 9800 34000 9830
rect 5060 9759 5380 9760
rect 7373 9482 7439 9485
rect 7649 9482 7715 9485
rect 7373 9480 7715 9482
rect 7373 9424 7378 9480
rect 7434 9424 7654 9480
rect 7710 9424 7715 9480
rect 7373 9422 7715 9424
rect 7373 9419 7439 9422
rect 7649 9419 7715 9422
rect 13813 9482 13879 9485
rect 14000 9482 34000 9512
rect 13813 9480 34000 9482
rect 13813 9424 13818 9480
rect 13874 9424 34000 9480
rect 13813 9422 34000 9424
rect 13813 9419 13879 9422
rect 14000 9392 34000 9422
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 7560 9280 7880 9281
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 9215 7880 9216
rect 13813 9074 13879 9077
rect 14000 9074 34000 9104
rect 13813 9072 34000 9074
rect 13813 9016 13818 9072
rect 13874 9016 34000 9072
rect 13813 9014 34000 9016
rect 13813 9011 13879 9014
rect 14000 8984 34000 9014
rect 5073 8938 5139 8941
rect 7557 8938 7623 8941
rect 5073 8936 7623 8938
rect 5073 8880 5078 8936
rect 5134 8880 7562 8936
rect 7618 8880 7623 8936
rect 5073 8878 7623 8880
rect 5073 8875 5139 8878
rect 7557 8875 7623 8878
rect 5060 8736 5380 8737
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 8671 5380 8672
rect 6913 8666 6979 8669
rect 7281 8666 7347 8669
rect 6913 8664 7347 8666
rect 6913 8608 6918 8664
rect 6974 8608 7286 8664
rect 7342 8608 7347 8664
rect 6913 8606 7347 8608
rect 6913 8603 6979 8606
rect 7281 8603 7347 8606
rect 13721 8666 13787 8669
rect 14000 8666 34000 8696
rect 13721 8664 34000 8666
rect 13721 8608 13726 8664
rect 13782 8608 34000 8664
rect 13721 8606 34000 8608
rect 13721 8603 13787 8606
rect 14000 8576 34000 8606
rect 5441 8530 5507 8533
rect 7833 8530 7899 8533
rect 5441 8528 7899 8530
rect 5441 8472 5446 8528
rect 5502 8472 7838 8528
rect 7894 8472 7899 8528
rect 5441 8470 7899 8472
rect 5441 8467 5507 8470
rect 7833 8467 7899 8470
rect 8753 8258 8819 8261
rect 14000 8258 34000 8288
rect 8753 8256 34000 8258
rect 8753 8200 8758 8256
rect 8814 8200 34000 8256
rect 8753 8198 34000 8200
rect 8753 8195 8819 8198
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 7560 8192 7880 8193
rect 7560 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7880 8192
rect 14000 8168 34000 8198
rect 7560 8127 7880 8128
rect 5625 7850 5691 7853
rect 6637 7850 6703 7853
rect 5625 7848 6703 7850
rect 5625 7792 5630 7848
rect 5686 7792 6642 7848
rect 6698 7792 6703 7848
rect 5625 7790 6703 7792
rect 5625 7787 5691 7790
rect 6637 7787 6703 7790
rect 9581 7850 9647 7853
rect 14000 7850 34000 7880
rect 9581 7848 34000 7850
rect 9581 7792 9586 7848
rect 9642 7792 34000 7848
rect 9581 7790 34000 7792
rect 9581 7787 9647 7790
rect 14000 7760 34000 7790
rect 5060 7648 5380 7649
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 7583 5380 7584
rect 2773 7442 2839 7445
rect 3877 7442 3943 7445
rect 2773 7440 3943 7442
rect 2773 7384 2778 7440
rect 2834 7384 3882 7440
rect 3938 7384 3943 7440
rect 2773 7382 3943 7384
rect 2773 7379 2839 7382
rect 3877 7379 3943 7382
rect 7465 7442 7531 7445
rect 8753 7442 8819 7445
rect 7465 7440 8819 7442
rect 7465 7384 7470 7440
rect 7526 7384 8758 7440
rect 8814 7384 8819 7440
rect 7465 7382 8819 7384
rect 7465 7379 7531 7382
rect 8753 7379 8819 7382
rect 13537 7442 13603 7445
rect 14000 7442 34000 7472
rect 13537 7440 34000 7442
rect 13537 7384 13542 7440
rect 13598 7384 34000 7440
rect 13537 7382 34000 7384
rect 13537 7379 13603 7382
rect 14000 7352 34000 7382
rect 6085 7306 6151 7309
rect 6085 7304 12450 7306
rect 6085 7248 6090 7304
rect 6146 7248 12450 7304
rect 6085 7246 12450 7248
rect 6085 7243 6151 7246
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 7560 7104 7880 7105
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 7039 7880 7040
rect 12390 7034 12450 7246
rect 14000 7034 34000 7064
rect 12390 6974 34000 7034
rect 14000 6944 34000 6974
rect 13721 6626 13787 6629
rect 14000 6626 34000 6656
rect 13721 6624 34000 6626
rect 13721 6568 13726 6624
rect 13782 6568 34000 6624
rect 13721 6566 34000 6568
rect 13721 6563 13787 6566
rect 5060 6560 5380 6561
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 14000 6536 34000 6566
rect 5060 6495 5380 6496
rect 2681 6218 2747 6221
rect 6821 6218 6887 6221
rect 2681 6216 6887 6218
rect 2681 6160 2686 6216
rect 2742 6160 6826 6216
rect 6882 6160 6887 6216
rect 2681 6158 6887 6160
rect 2681 6155 2747 6158
rect 6821 6155 6887 6158
rect 9489 6218 9555 6221
rect 14000 6218 34000 6248
rect 9489 6216 34000 6218
rect 9489 6160 9494 6216
rect 9550 6160 34000 6216
rect 9489 6158 34000 6160
rect 9489 6155 9555 6158
rect 14000 6128 34000 6158
rect 2560 6016 2880 6017
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5951 2880 5952
rect 7560 6016 7880 6017
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 5951 7880 5952
rect 9489 5810 9555 5813
rect 14000 5810 34000 5840
rect 9489 5808 34000 5810
rect 9489 5752 9494 5808
rect 9550 5752 34000 5808
rect 9489 5750 34000 5752
rect 9489 5747 9555 5750
rect 14000 5720 34000 5750
rect 5060 5472 5380 5473
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 5407 5380 5408
rect 8201 5402 8267 5405
rect 14000 5402 34000 5432
rect 8201 5400 34000 5402
rect 8201 5344 8206 5400
rect 8262 5344 34000 5400
rect 8201 5342 34000 5344
rect 8201 5339 8267 5342
rect 14000 5312 34000 5342
rect 4797 5130 4863 5133
rect 4797 5128 12450 5130
rect 4797 5072 4802 5128
rect 4858 5072 12450 5128
rect 4797 5070 12450 5072
rect 4797 5067 4863 5070
rect 12390 4994 12450 5070
rect 14000 4994 34000 5024
rect 12390 4934 34000 4994
rect 7560 4928 7880 4929
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 14000 4904 34000 4934
rect 7560 4863 7880 4864
rect 9857 4586 9923 4589
rect 14000 4586 34000 4616
rect 9857 4584 34000 4586
rect 9857 4528 9862 4584
rect 9918 4528 34000 4584
rect 9857 4526 34000 4528
rect 9857 4523 9923 4526
rect 14000 4496 34000 4526
rect 5060 4384 5380 4385
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 4319 5380 4320
rect 13813 4178 13879 4181
rect 14000 4178 34000 4208
rect 13813 4176 34000 4178
rect 13813 4120 13818 4176
rect 13874 4120 34000 4176
rect 13813 4118 34000 4120
rect 13813 4115 13879 4118
rect 14000 4088 34000 4118
rect 7560 3840 7880 3841
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 3775 7880 3776
rect 8937 3770 9003 3773
rect 14000 3770 34000 3800
rect 8937 3768 34000 3770
rect 8937 3712 8942 3768
rect 8998 3712 34000 3768
rect 8937 3710 34000 3712
rect 8937 3707 9003 3710
rect 14000 3680 34000 3710
rect 2773 3498 2839 3501
rect 2730 3496 2839 3498
rect 2730 3440 2778 3496
rect 2834 3440 2839 3496
rect 2730 3438 2839 3440
rect 2484 3435 2839 3438
rect 2484 3378 2790 3435
rect 6821 3362 6887 3365
rect 14000 3362 34000 3392
rect 6821 3360 34000 3362
rect 6821 3304 6826 3360
rect 6882 3304 34000 3360
rect 6821 3302 34000 3304
rect 6821 3299 6887 3302
rect 5060 3296 5380 3297
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 14000 3272 34000 3302
rect 5060 3231 5380 3232
rect 8201 2954 8267 2957
rect 14000 2954 34000 2984
rect 8201 2952 34000 2954
rect 8201 2896 8206 2952
rect 8262 2896 34000 2952
rect 8201 2894 34000 2896
rect 8201 2891 8267 2894
rect 14000 2864 34000 2894
rect 7560 2752 7880 2753
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 2687 7880 2688
rect 14000 2546 34000 2576
rect 6870 2486 34000 2546
rect 6361 2410 6427 2413
rect 6870 2410 6930 2486
rect 14000 2456 34000 2486
rect 6361 2408 6930 2410
rect 6361 2352 6366 2408
rect 6422 2352 6930 2408
rect 6361 2350 6930 2352
rect 6361 2347 6427 2350
rect 5060 2208 5380 2209
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 2143 5380 2144
rect 9213 2138 9279 2141
rect 14000 2138 34000 2168
rect 9213 2136 34000 2138
rect 9213 2080 9218 2136
rect 9274 2080 34000 2136
rect 9213 2078 34000 2080
rect 9213 2075 9279 2078
rect 14000 2048 34000 2078
rect 9581 1730 9647 1733
rect 14000 1730 34000 1760
rect 9581 1728 34000 1730
rect 9581 1672 9586 1728
rect 9642 1672 34000 1728
rect 9581 1670 34000 1672
rect 9581 1667 9647 1670
rect 7560 1664 7880 1665
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 14000 1640 34000 1670
rect 7560 1599 7880 1600
rect 14000 1320 34000 1352
rect 14000 1264 16578 1320
rect 16634 1264 34000 1320
rect 14000 1232 34000 1264
rect 5060 1120 5380 1121
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 5060 1055 5380 1056
rect 9397 914 9463 917
rect 14000 914 34000 944
rect 9397 912 34000 914
rect 9397 856 9402 912
rect 9458 856 34000 912
rect 9397 854 34000 856
rect 9397 851 9463 854
rect 14000 824 34000 854
rect 9489 506 9555 509
rect 14000 506 34000 536
rect 9489 504 34000 506
rect 9489 448 9494 504
rect 9550 448 34000 504
rect 9489 446 34000 448
rect 9489 443 9555 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 5068 1116 5132 1120
rect 5068 1060 5072 1116
rect 5072 1060 5128 1116
rect 5128 1060 5132 1116
rect 5068 1056 5132 1060
rect 5148 1116 5212 1120
rect 5148 1060 5152 1116
rect 5152 1060 5208 1116
rect 5208 1060 5212 1116
rect 5148 1056 5212 1060
rect 5228 1116 5292 1120
rect 5228 1060 5232 1116
rect 5232 1060 5288 1116
rect 5288 1060 5292 1116
rect 5228 1056 5292 1060
rect 5308 1116 5372 1120
rect 5308 1060 5312 1116
rect 5312 1060 5368 1116
rect 5368 1060 5372 1116
rect 5308 1056 5372 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1088 2880 1222
rect 3560 9266 3880 11424
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1088 3880 2270
rect 5060 10912 5380 11472
rect 7560 11456 7880 11472
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 9908 5380 10848
rect 5060 9824 5102 9908
rect 5338 9824 5380 9908
rect 5060 9760 5068 9824
rect 5372 9760 5380 9824
rect 5060 9672 5102 9760
rect 5338 9672 5380 9760
rect 5060 8736 5380 9672
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 6560 5380 7584
rect 5060 6496 5068 6560
rect 5132 6528 5148 6560
rect 5212 6528 5228 6560
rect 5292 6528 5308 6560
rect 5372 6496 5380 6560
rect 5060 6292 5102 6496
rect 5338 6292 5380 6496
rect 5060 5472 5380 6292
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3296 5380 4320
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 3148 5380 3232
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2208 5380 2912
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1120 5380 2144
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 6060 10956 6380 11424
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 1088 6380 3960
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 8218 7880 9216
rect 7560 8192 7602 8218
rect 7838 8192 7880 8218
rect 7560 8128 7568 8192
rect 7872 8128 7880 8192
rect 7560 7982 7602 8128
rect 7838 7982 7880 8128
rect 7560 7104 7880 7982
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 4928 7880 5952
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 4838 7880 4864
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 3840 7880 4602
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1458 7880 1600
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 5060 1040 5380 1056
rect 7560 1040 7880 1222
rect 8560 9266 8880 11424
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 8560 1088 8880 2270
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 5102 9824 5338 9908
rect 5102 9760 5132 9824
rect 5132 9760 5148 9824
rect 5148 9760 5212 9824
rect 5212 9760 5228 9824
rect 5228 9760 5292 9824
rect 5292 9760 5308 9824
rect 5308 9760 5338 9824
rect 5102 9672 5338 9760
rect 5102 6496 5132 6528
rect 5132 6496 5148 6528
rect 5148 6496 5212 6528
rect 5212 6496 5228 6528
rect 5228 6496 5292 6528
rect 5292 6496 5308 6528
rect 5308 6496 5338 6528
rect 5102 6292 5338 6496
rect 5102 2912 5338 3148
rect 6102 10720 6338 10956
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 7602 8192 7838 8218
rect 7602 8128 7632 8192
rect 7632 8128 7648 8192
rect 7648 8128 7712 8192
rect 7712 8128 7728 8192
rect 7728 8128 7792 8192
rect 7792 8128 7808 8192
rect 7808 8128 7838 8192
rect 7602 7982 7838 8128
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 920 10956 9844 10998
rect 920 10720 6102 10956
rect 6338 10720 9844 10956
rect 920 10678 9844 10720
rect 920 9908 9844 9950
rect 920 9672 5102 9908
rect 5338 9672 9844 9908
rect 920 9630 9844 9672
rect 920 9266 9844 9308
rect 920 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 9844 9266
rect 920 8988 9844 9030
rect 920 8218 9844 8260
rect 920 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 9844 8218
rect 920 7940 9844 7982
rect 920 7576 9844 7618
rect 920 7340 6102 7576
rect 6338 7340 9844 7576
rect 920 7298 9844 7340
rect 920 6528 9844 6570
rect 920 6292 5102 6528
rect 5338 6292 9844 6528
rect 920 6250 9844 6292
rect 920 5886 9844 5928
rect 920 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 9844 5886
rect 920 5608 9844 5650
rect 920 4838 9844 4880
rect 920 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 9844 4838
rect 920 4560 9844 4602
rect 920 4196 9844 4238
rect 920 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 9844 4196
rect 920 3918 9844 3960
rect 920 3148 9844 3190
rect 920 2912 5102 3148
rect 5338 2912 9844 3148
rect 920 2870 9844 2912
rect 920 2506 9844 2548
rect 920 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 9844 2506
rect 920 2228 9844 2270
rect 920 1458 9844 1500
rect 920 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 9844 1458
rect 920 1180 9844 1222
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__B
timestamp 1648946573
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A2
timestamp 1648946573
transform -1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1648946573
transform 1 0 9200 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1648946573
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1648946573
transform -1 0 9476 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1648946573
transform 1 0 9384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1648946573
transform 1 0 3680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__B
timestamp 1648946573
transform -1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1648946573
transform 1 0 5152 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__B_N
timestamp 1648946573
transform 1 0 1288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__B
timestamp 1648946573
transform -1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__B_N
timestamp 1648946573
transform -1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__B
timestamp 1648946573
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__B_N
timestamp 1648946573
transform -1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__B
timestamp 1648946573
transform 1 0 5704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__B_N
timestamp 1648946573
transform -1 0 6072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__B
timestamp 1648946573
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__B_N
timestamp 1648946573
transform 1 0 3864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__B
timestamp 1648946573
transform -1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__B_N
timestamp 1648946573
transform 1 0 3588 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__B
timestamp 1648946573
transform -1 0 8280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__B_N
timestamp 1648946573
transform -1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__B
timestamp 1648946573
transform -1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__B_N
timestamp 1648946573
transform 1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__B
timestamp 1648946573
transform -1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__B_N
timestamp 1648946573
transform -1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__B
timestamp 1648946573
transform -1 0 5336 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__B_N
timestamp 1648946573
transform -1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__B
timestamp 1648946573
transform -1 0 3680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__B_N
timestamp 1648946573
transform -1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__B
timestamp 1648946573
transform -1 0 5888 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__B_N
timestamp 1648946573
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__B
timestamp 1648946573
transform -1 0 1472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__B_N
timestamp 1648946573
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__D
timestamp 1648946573
transform -1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__RESET_B
timestamp 1648946573
transform -1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__RESET_B
timestamp 1648946573
transform -1 0 1472 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__RESET_B
timestamp 1648946573
transform 1 0 1472 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__RESET_B
timestamp 1648946573
transform -1 0 1472 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__RESET_B
timestamp 1648946573
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__RESET_B
timestamp 1648946573
transform 1 0 5888 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__RESET_B
timestamp 1648946573
transform 1 0 4048 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__RESET_B
timestamp 1648946573
transform 1 0 7820 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__RESET_B
timestamp 1648946573
transform 1 0 8280 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__RESET_B
timestamp 1648946573
transform -1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__RESET_B
timestamp 1648946573
transform -1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__RESET_B
timestamp 1648946573
transform -1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__RESET_B
timestamp 1648946573
transform 1 0 8464 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1648946573
transform -1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1648946573
transform -1 0 8188 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1648946573
transform -1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1648946573
transform -1 0 7084 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 5244 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84
timestamp 1648946573
transform 1 0 8648 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1648946573
transform 1 0 9476 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 3312 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_78
timestamp 1648946573
transform 1 0 8096 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1648946573
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_26
timestamp 1648946573
transform 1 0 3312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1648946573
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_83
timestamp 1648946573
transform 1 0 8556 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1648946573
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_26
timestamp 1648946573
transform 1 0 3312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_32
timestamp 1648946573
transform 1 0 3864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1648946573
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_34
timestamp 1648946573
transform 1 0 4048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1648946573
transform 1 0 1196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1648946573
transform 1 0 1196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1648946573
transform 1 0 3404 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_24
timestamp 1648946573
transform 1 0 3128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1648946573
transform 1 0 6440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1648946573
transform 1 0 1196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1648946573
transform 1 0 8556 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1648946573
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1648946573
transform 1 0 1196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_69
timestamp 1648946573
transform 1 0 7268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1648946573
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_42
timestamp 1648946573
transform 1 0 4784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1648946573
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 1648946573
transform 1 0 3128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_93
timestamp 1648946573
transform 1 0 9476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1648946573
transform 1 0 1196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1648946573
transform 1 0 3404 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1648946573
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1648946573
transform 1 0 1196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_45
timestamp 1648946573
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_48
timestamp 1648946573
transform 1 0 5336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 1196 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1648946573
transform 1 0 3404 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_31
timestamp 1648946573
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 6716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1648946573
transform 1 0 8556 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1648946573
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1648946573
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1648946573
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1648946573
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1648946573
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1648946573
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1648946573
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1648946573
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1648946573
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1648946573
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1648946573
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1648946573
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1648946573
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1648946573
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1648946573
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1648946573
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1648946573
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1648946573
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1648946573
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1648946573
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1648946573
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1648946573
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1648946573
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1648946573
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1648946573
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1648946573
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1648946573
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1648946573
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1648946573
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1648946573
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1648946573
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1648946573
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1648946573
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1648946573
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1648946573
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1648946573
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1648946573
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1648946573
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1648946573
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1648946573
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1648946573
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1648946573
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1648946573
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1648946573
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1648946573
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1648946573
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1648946573
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1648946573
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1648946573
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1648946573
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1648946573
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1648946573
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1648946573
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1648946573
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1648946573
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1648946573
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1648946573
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1648946573
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1648946573
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1648946573
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1648946573
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1648946573
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1648946573
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1648946573
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_2  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8740 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8740 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 5980 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9384 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1648946573
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8740 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9384 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o22ai_2  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 8648 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1648946573
transform -1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 9292 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _108_
timestamp 1648946573
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _109_
timestamp 1648946573
transform -1 0 3588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 2484 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _111_
timestamp 1648946573
transform 1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1648946573
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113__4
timestamp 1648946573
transform -1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _114_
timestamp 1648946573
transform -1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _115_
timestamp 1648946573
transform -1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _116_
timestamp 1648946573
transform -1 0 3404 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _117_
timestamp 1648946573
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _118_
timestamp 1648946573
transform 1 0 2760 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp 1648946573
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120__5
timestamp 1648946573
transform -1 0 3496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _121_
timestamp 1648946573
transform 1 0 3588 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _122_
timestamp 1648946573
transform -1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _123_
timestamp 1648946573
transform -1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _124_
timestamp 1648946573
transform 1 0 6164 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _125_
timestamp 1648946573
transform 1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126__6
timestamp 1648946573
transform -1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _127_
timestamp 1648946573
transform 1 0 6164 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp 1648946573
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _129_
timestamp 1648946573
transform 1 0 4968 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _130_
timestamp 1648946573
transform 1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131__7
timestamp 1648946573
transform 1 0 7452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _132_
timestamp 1648946573
transform 1 0 5428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _133_
timestamp 1648946573
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _134_
timestamp 1648946573
transform 1 0 4508 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 1648946573
transform -1 0 5704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136__8
timestamp 1648946573
transform 1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _137_
timestamp 1648946573
transform 1 0 4416 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _138_
timestamp 1648946573
transform 1 0 4232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _139_
timestamp 1648946573
transform 1 0 4692 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _140_
timestamp 1648946573
transform -1 0 6440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1648946573
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142__9
timestamp 1648946573
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1648946573
transform -1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _144_
timestamp 1648946573
transform -1 0 4416 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp 1648946573
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _146_
timestamp 1648946573
transform -1 0 5612 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1648946573
transform 1 0 4416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148__10
timestamp 1648946573
transform -1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _149_
timestamp 1648946573
transform 1 0 5060 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1648946573
transform -1 0 6440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _151_
timestamp 1648946573
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _152_
timestamp 1648946573
transform -1 0 8556 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp 1648946573
transform 1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154__11
timestamp 1648946573
transform 1 0 7452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _155_
timestamp 1648946573
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1648946573
transform -1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _157_
timestamp 1648946573
transform 1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp 1648946573
transform -1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159__12
timestamp 1648946573
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _160_
timestamp 1648946573
transform 1 0 8280 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1648946573
transform -1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _162_
timestamp 1648946573
transform 1 0 6992 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp 1648946573
transform -1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164__13
timestamp 1648946573
transform -1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _165_
timestamp 1648946573
transform 1 0 8004 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _166_
timestamp 1648946573
transform -1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _167_
timestamp 1648946573
transform 1 0 4968 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp 1648946573
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169__1
timestamp 1648946573
transform -1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _170_
timestamp 1648946573
transform 1 0 3680 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp 1648946573
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _172_
timestamp 1648946573
transform 1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1648946573
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174__2
timestamp 1648946573
transform -1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _175_
timestamp 1648946573
transform 1 0 4324 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _176_
timestamp 1648946573
transform -1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _177_
timestamp 1648946573
transform 1 0 5612 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _178_
timestamp 1648946573
transform 1 0 7544 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179__3
timestamp 1648946573
transform 1 0 5336 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _180_
timestamp 1648946573
transform -1 0 5152 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp 1648946573
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 1840 0 -1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _183_
timestamp 1648946573
transform 1 0 1840 0 -1 8704
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _184_
timestamp 1648946573
transform 1 0 6072 0 1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _185_
timestamp 1648946573
transform 1 0 6900 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _186_
timestamp 1648946573
transform 1 0 3496 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _187_
timestamp 1648946573
transform 1 0 3312 0 -1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _188_
timestamp 1648946573
transform 1 0 3496 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _189_
timestamp 1648946573
transform 1 0 6532 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _190_
timestamp 1648946573
transform 1 0 6440 0 1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _191_
timestamp 1648946573
transform 1 0 6716 0 1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _192_
timestamp 1648946573
transform 1 0 3588 0 -1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _193_
timestamp 1648946573
transform 1 0 4232 0 -1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _194_
timestamp 1648946573
transform 1 0 5704 0 1 2176
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_2  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 3128 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _196_
timestamp 1648946573
transform 1 0 1564 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _197_
timestamp 1648946573
transform -1 0 3128 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _198_
timestamp 1648946573
transform 1 0 1472 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _199_
timestamp 1648946573
transform -1 0 3496 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _200_
timestamp 1648946573
transform 1 0 3312 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _201_
timestamp 1648946573
transform 1 0 3312 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _202_
timestamp 1648946573
transform 1 0 4232 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _203_
timestamp 1648946573
transform 1 0 6164 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _204_
timestamp 1648946573
transform 1 0 6164 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _205_
timestamp 1648946573
transform 1 0 7360 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _206_
timestamp 1648946573
transform -1 0 7728 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _207_
timestamp 1648946573
transform 1 0 6256 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8280 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _209_
timestamp 1648946573
transform 1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _210_
timestamp 1648946573
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8648 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 5152 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__077_
timestamp 1648946573
transform -1 0 6072 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock
timestamp 1648946573
transform -1 0 8004 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1648946573
transform -1 0 8004 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__077_
timestamp 1648946573
transform 1 0 1472 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock
timestamp 1648946573
transform -1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_load
timestamp 1648946573
transform -1 0 4508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__049_
timestamp 1648946573
transform -1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__077_
timestamp 1648946573
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1648946573
transform -1 0 5520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_load
timestamp 1648946573
transform -1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd2_1  data_delay_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 8280 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd2_1  data_delay_2
timestamp 1648946573
transform 1 0 8924 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 4416 0 1 5440
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 1638030917
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 1656 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform 1 0 3312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1648946573
transform -1 0 9016 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1648946573
transform -1 0 8188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1648946573
transform -1 0 9476 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold6
timestamp 1648946573
transform -1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1648946573
transform 1 0 3588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1648946573
transform 1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1648946573
transform 1 0 1288 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold10
timestamp 1648946573
transform 1 0 2024 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1648946573
transform 1 0 1288 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold12
timestamp 1648946573
transform 1 0 2024 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1648946573
transform 1 0 3588 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold14
timestamp 1648946573
transform -1 0 5060 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1648946573
transform -1 0 9016 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold16
timestamp 1648946573
transform -1 0 8188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold17
timestamp 1648946573
transform 1 0 8740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold18
timestamp 1648946573
transform 1 0 5060 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1648946573
transform 1 0 6072 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold20
timestamp 1648946573
transform -1 0 6440 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold21
timestamp 1648946573
transform -1 0 7544 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1648946573
transform -1 0 9476 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1648946573
transform 1 0 6624 0 1 7616
box -38 -48 774 592
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 42 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 42 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 7560 1040 7880 11472 6 vccd
port 42 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 43 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 43 nsew power input
rlabel metal4 s 8560 1088 8880 11424 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 44 nsew ground input
rlabel metal4 s 5060 1040 5380 11472 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 45 nsew ground input
rlabel metal4 s 6060 1088 6380 11424 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
