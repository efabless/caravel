magic
tech sky130A
magscale 1 2
timestamp 1637516397
<< error_s >>
rect 55754 272986 55762 273304
rect 55754 272984 56074 272986
<< metal1 >>
rect 145190 1007428 145196 1007480
rect 145248 1007468 145254 1007480
rect 154574 1007468 154580 1007480
rect 145248 1007440 154580 1007468
rect 145248 1007428 145254 1007440
rect 154574 1007428 154580 1007440
rect 154632 1007428 154638 1007480
rect 501322 1007360 501328 1007412
rect 501380 1007400 501386 1007412
rect 517330 1007400 517336 1007412
rect 501380 1007372 517336 1007400
rect 501380 1007360 501386 1007372
rect 517330 1007360 517336 1007372
rect 517388 1007360 517394 1007412
rect 424686 1006000 424692 1006052
rect 424744 1006040 424750 1006052
rect 466454 1006040 466460 1006052
rect 424744 1006012 466460 1006040
rect 424744 1006000 424750 1006012
rect 466454 1006000 466460 1006012
rect 466512 1006000 466518 1006052
rect 423858 1005864 423864 1005916
rect 423916 1005904 423922 1005916
rect 440142 1005904 440148 1005916
rect 423916 1005876 440148 1005904
rect 423916 1005864 423922 1005876
rect 440142 1005864 440148 1005876
rect 440200 1005864 440206 1005916
rect 424318 1005796 424324 1005848
rect 424376 1005836 424382 1005848
rect 440418 1005836 440424 1005848
rect 424376 1005808 440424 1005836
rect 424376 1005796 424382 1005808
rect 440418 1005796 440424 1005808
rect 440476 1005796 440482 1005848
rect 503346 1005796 503352 1005848
rect 503404 1005836 503410 1005848
rect 520182 1005836 520188 1005848
rect 503404 1005808 520188 1005836
rect 503404 1005796 503410 1005808
rect 520182 1005796 520188 1005808
rect 520240 1005796 520246 1005848
rect 502978 1005728 502984 1005780
rect 503036 1005768 503042 1005780
rect 519998 1005768 520004 1005780
rect 503036 1005740 520004 1005768
rect 503036 1005728 503042 1005740
rect 519998 1005728 520004 1005740
rect 520056 1005728 520062 1005780
rect 356054 1005660 356060 1005712
rect 356112 1005700 356118 1005712
rect 374270 1005700 374276 1005712
rect 356112 1005672 374276 1005700
rect 356112 1005660 356118 1005672
rect 374270 1005660 374276 1005672
rect 374328 1005660 374334 1005712
rect 502518 1005660 502524 1005712
rect 502576 1005700 502582 1005712
rect 519170 1005700 519176 1005712
rect 502576 1005672 519176 1005700
rect 502576 1005660 502582 1005672
rect 519170 1005660 519176 1005672
rect 519228 1005660 519234 1005712
rect 356514 1005592 356520 1005644
rect 356572 1005632 356578 1005644
rect 377306 1005632 377312 1005644
rect 356572 1005604 377312 1005632
rect 356572 1005592 356578 1005604
rect 377306 1005592 377312 1005604
rect 377364 1005592 377370 1005644
rect 504542 1005592 504548 1005644
rect 504600 1005632 504606 1005644
rect 517238 1005632 517244 1005644
rect 504600 1005604 517244 1005632
rect 504600 1005592 504606 1005604
rect 517238 1005592 517244 1005604
rect 517296 1005592 517302 1005644
rect 200022 1005524 200028 1005576
rect 200080 1005564 200086 1005576
rect 207198 1005564 207204 1005576
rect 200080 1005536 207204 1005564
rect 200080 1005524 200086 1005536
rect 207198 1005524 207204 1005536
rect 207256 1005524 207262 1005576
rect 505830 1005524 505836 1005576
rect 505888 1005564 505894 1005576
rect 517606 1005564 517612 1005576
rect 505888 1005536 517612 1005564
rect 505888 1005524 505894 1005536
rect 517606 1005524 517612 1005536
rect 517664 1005524 517670 1005576
rect 144822 1005456 144828 1005508
rect 144880 1005496 144886 1005508
rect 160278 1005496 160284 1005508
rect 144880 1005468 160284 1005496
rect 144880 1005456 144886 1005468
rect 160278 1005456 160284 1005468
rect 160336 1005456 160342 1005508
rect 195330 1005456 195336 1005508
rect 195388 1005496 195394 1005508
rect 209590 1005496 209596 1005508
rect 195388 1005468 209596 1005496
rect 195388 1005456 195394 1005468
rect 209590 1005456 209596 1005468
rect 209648 1005456 209654 1005508
rect 361022 1005456 361028 1005508
rect 361080 1005496 361086 1005508
rect 377950 1005496 377956 1005508
rect 361080 1005468 377956 1005496
rect 361080 1005456 361086 1005468
rect 377950 1005456 377956 1005468
rect 378008 1005456 378014 1005508
rect 505370 1005456 505376 1005508
rect 505428 1005496 505434 1005508
rect 517422 1005496 517428 1005508
rect 505428 1005468 517428 1005496
rect 505428 1005456 505434 1005468
rect 517422 1005456 517428 1005468
rect 517480 1005456 517486 1005508
rect 145098 1005388 145104 1005440
rect 145156 1005428 145162 1005440
rect 154942 1005428 154948 1005440
rect 145156 1005400 154948 1005428
rect 145156 1005388 145162 1005400
rect 154942 1005388 154948 1005400
rect 155000 1005388 155006 1005440
rect 92494 1005320 92500 1005372
rect 92552 1005360 92558 1005372
rect 109310 1005360 109316 1005372
rect 92552 1005332 109316 1005360
rect 92552 1005320 92558 1005332
rect 109310 1005320 109316 1005332
rect 109368 1005320 109374 1005372
rect 145006 1005320 145012 1005372
rect 145064 1005360 145070 1005372
rect 153746 1005360 153752 1005372
rect 145064 1005332 153752 1005360
rect 145064 1005320 145070 1005332
rect 153746 1005320 153752 1005332
rect 153804 1005320 153810 1005372
rect 360194 1005320 360200 1005372
rect 360252 1005360 360258 1005372
rect 380802 1005360 380808 1005372
rect 360252 1005332 380808 1005360
rect 360252 1005320 360258 1005332
rect 380802 1005320 380808 1005332
rect 380860 1005320 380866 1005372
rect 423490 1005320 423496 1005372
rect 423548 1005360 423554 1005372
rect 467834 1005360 467840 1005372
rect 423548 1005332 467840 1005360
rect 423548 1005320 423554 1005332
rect 467834 1005320 467840 1005332
rect 467892 1005320 467898 1005372
rect 144914 1005252 144920 1005304
rect 144972 1005292 144978 1005304
rect 153286 1005292 153292 1005304
rect 144972 1005264 153292 1005292
rect 144972 1005252 144978 1005264
rect 153286 1005252 153292 1005264
rect 153344 1005252 153350 1005304
rect 259822 1005252 259828 1005304
rect 259880 1005292 259886 1005304
rect 280338 1005292 280344 1005304
rect 259880 1005264 280344 1005292
rect 259880 1005252 259886 1005264
rect 280338 1005252 280344 1005264
rect 280396 1005252 280402 1005304
rect 428366 1005252 428372 1005304
rect 428424 1005292 428430 1005304
rect 453942 1005292 453948 1005304
rect 428424 1005264 453948 1005292
rect 428424 1005252 428430 1005264
rect 453942 1005252 453948 1005264
rect 454000 1005252 454006 1005304
rect 148870 1005184 148876 1005236
rect 148928 1005224 148934 1005236
rect 151262 1005224 151268 1005236
rect 148928 1005196 151268 1005224
rect 148928 1005184 148934 1005196
rect 151262 1005184 151268 1005196
rect 151320 1005184 151326 1005236
rect 260190 1005184 260196 1005236
rect 260248 1005224 260254 1005236
rect 265250 1005224 265256 1005236
rect 260248 1005196 265256 1005224
rect 260248 1005184 260254 1005196
rect 265250 1005184 265256 1005196
rect 265308 1005184 265314 1005236
rect 359734 1005184 359740 1005236
rect 359792 1005224 359798 1005236
rect 370406 1005224 370412 1005236
rect 359792 1005196 370412 1005224
rect 359792 1005184 359798 1005196
rect 370406 1005184 370412 1005196
rect 370464 1005184 370470 1005236
rect 106458 1005116 106464 1005168
rect 106516 1005156 106522 1005168
rect 125594 1005156 125600 1005168
rect 106516 1005128 125600 1005156
rect 106516 1005116 106522 1005128
rect 125594 1005116 125600 1005128
rect 125652 1005116 125658 1005168
rect 201862 1005116 201868 1005168
rect 201920 1005156 201926 1005168
rect 227622 1005156 227628 1005168
rect 201920 1005128 227628 1005156
rect 201920 1005116 201926 1005128
rect 227622 1005116 227628 1005128
rect 227680 1005116 227686 1005168
rect 261846 1005116 261852 1005168
rect 261904 1005156 261910 1005168
rect 261904 1005128 265774 1005156
rect 261904 1005116 261910 1005128
rect 149698 1005048 149704 1005100
rect 149756 1005088 149762 1005100
rect 150434 1005088 150440 1005100
rect 149756 1005060 150440 1005088
rect 149756 1005048 149762 1005060
rect 150434 1005048 150440 1005060
rect 150492 1005088 150498 1005100
rect 175182 1005088 175188 1005100
rect 150492 1005060 175188 1005088
rect 150492 1005048 150498 1005060
rect 175182 1005048 175188 1005060
rect 175240 1005048 175246 1005100
rect 208394 1005048 208400 1005100
rect 208452 1005088 208458 1005100
rect 227806 1005088 227812 1005100
rect 208452 1005060 227812 1005088
rect 208452 1005048 208458 1005060
rect 227806 1005048 227812 1005060
rect 227864 1005048 227870 1005100
rect 263042 1005048 263048 1005100
rect 263100 1005088 263106 1005100
rect 265530 1005088 265536 1005100
rect 263100 1005060 265536 1005088
rect 263100 1005048 263106 1005060
rect 265530 1005048 265536 1005060
rect 265588 1005048 265594 1005100
rect 265746 1005088 265774 1005128
rect 504174 1005116 504180 1005168
rect 504232 1005156 504238 1005168
rect 520366 1005156 520372 1005168
rect 504232 1005128 520372 1005156
rect 504232 1005116 504238 1005128
rect 520366 1005116 520372 1005128
rect 520424 1005116 520430 1005168
rect 270462 1005088 270468 1005100
rect 265746 1005060 270468 1005088
rect 270462 1005048 270468 1005060
rect 270520 1005048 270526 1005100
rect 358170 1005048 358176 1005100
rect 358228 1005088 358234 1005100
rect 366726 1005088 366732 1005100
rect 358228 1005060 366732 1005088
rect 358228 1005048 358234 1005060
rect 366726 1005048 366732 1005060
rect 366784 1005048 366790 1005100
rect 428826 1005048 428832 1005100
rect 428884 1005088 428890 1005100
rect 464246 1005088 464252 1005100
rect 428884 1005060 464252 1005088
rect 428884 1005048 428890 1005060
rect 464246 1005048 464252 1005060
rect 464304 1005048 464310 1005100
rect 551922 1005048 551928 1005100
rect 551980 1005088 551986 1005100
rect 568574 1005088 568580 1005100
rect 551980 1005060 568580 1005088
rect 551980 1005048 551986 1005060
rect 568574 1005048 568580 1005060
rect 568632 1005048 568638 1005100
rect 148870 1004980 148876 1005032
rect 148928 1005020 148934 1005032
rect 150894 1005020 150900 1005032
rect 148928 1004992 150900 1005020
rect 148928 1004980 148934 1004992
rect 150894 1004980 150900 1004992
rect 150952 1004980 150958 1005032
rect 211614 1005020 211620 1005032
rect 206986 1004992 211620 1005020
rect 148134 1004912 148140 1004964
rect 148192 1004952 148198 1004964
rect 154114 1004952 154120 1004964
rect 148192 1004924 154120 1004952
rect 148192 1004912 148198 1004924
rect 154114 1004912 154120 1004924
rect 154172 1004912 154178 1004964
rect 159450 1004912 159456 1004964
rect 159508 1004952 159514 1004964
rect 173894 1004952 173900 1004964
rect 159508 1004924 173900 1004952
rect 159508 1004912 159514 1004924
rect 173894 1004912 173900 1004924
rect 173952 1004912 173958 1004964
rect 204162 1004912 204168 1004964
rect 204220 1004952 204226 1004964
rect 206986 1004952 207014 1004992
rect 211614 1004980 211620 1004992
rect 211672 1004980 211678 1005032
rect 260650 1004980 260656 1005032
rect 260708 1005020 260714 1005032
rect 260708 1004992 265774 1005020
rect 260708 1004980 260714 1004992
rect 204220 1004924 207014 1004952
rect 204220 1004912 204226 1004924
rect 209222 1004912 209228 1004964
rect 209280 1004952 209286 1004964
rect 227714 1004952 227720 1004964
rect 209280 1004924 227720 1004952
rect 209280 1004912 209286 1004924
rect 227714 1004912 227720 1004924
rect 227772 1004912 227778 1004964
rect 262674 1004912 262680 1004964
rect 262732 1004952 262738 1004964
rect 265530 1004952 265536 1004964
rect 262732 1004924 265536 1004952
rect 262732 1004912 262738 1004924
rect 265530 1004912 265536 1004924
rect 265588 1004912 265594 1004964
rect 265746 1004952 265774 1004992
rect 356882 1004980 356888 1005032
rect 356940 1005020 356946 1005032
rect 378042 1005020 378048 1005032
rect 356940 1004992 378048 1005020
rect 356940 1004980 356946 1004992
rect 378042 1004980 378048 1004992
rect 378100 1004980 378106 1005032
rect 425514 1004980 425520 1005032
rect 425572 1005020 425578 1005032
rect 455598 1005020 455604 1005032
rect 425572 1004992 455604 1005020
rect 425572 1004980 425578 1004992
rect 455598 1004980 455604 1004992
rect 455656 1004980 455662 1005032
rect 280154 1004952 280160 1004964
rect 265746 1004924 280160 1004952
rect 280154 1004912 280160 1004924
rect 280212 1004912 280218 1004964
rect 358538 1004912 358544 1004964
rect 358596 1004952 358602 1004964
rect 383092 1004952 383098 1004964
rect 358596 1004924 383098 1004952
rect 358596 1004912 358602 1004924
rect 383092 1004912 383098 1004924
rect 383150 1004912 383156 1004964
rect 426802 1004912 426808 1004964
rect 426860 1004952 426866 1004964
rect 455506 1004952 455512 1004964
rect 426860 1004924 455512 1004952
rect 426860 1004912 426866 1004924
rect 455506 1004912 455512 1004924
rect 455564 1004912 455570 1004964
rect 505002 1004912 505008 1004964
rect 505060 1004952 505066 1004964
rect 522942 1004952 522948 1004964
rect 505060 1004924 522948 1004952
rect 505060 1004912 505066 1004924
rect 522942 1004912 522948 1004924
rect 523000 1004912 523006 1004964
rect 551646 1004912 551652 1004964
rect 551704 1004952 551710 1004964
rect 554774 1004952 554780 1004964
rect 551704 1004924 554780 1004952
rect 551704 1004912 551710 1004924
rect 554774 1004912 554780 1004924
rect 554832 1004912 554838 1004964
rect 108022 1004844 108028 1004896
rect 108080 1004884 108086 1004896
rect 108080 1004856 109732 1004884
rect 108080 1004844 108086 1004856
rect 108850 1004816 108856 1004828
rect 102106 1004788 108856 1004816
rect 92954 1004708 92960 1004760
rect 93012 1004748 93018 1004760
rect 102106 1004748 102134 1004788
rect 108850 1004776 108856 1004788
rect 108908 1004776 108914 1004828
rect 109704 1004816 109732 1004856
rect 148870 1004844 148876 1004896
rect 148928 1004884 148934 1004896
rect 152090 1004884 152096 1004896
rect 148928 1004856 152096 1004884
rect 148928 1004844 148934 1004856
rect 152090 1004844 152096 1004856
rect 152148 1004844 152154 1004896
rect 210878 1004844 210884 1004896
rect 210936 1004884 210942 1004896
rect 210936 1004856 215692 1004884
rect 210936 1004844 210942 1004856
rect 125686 1004816 125692 1004828
rect 109704 1004788 125692 1004816
rect 125686 1004776 125692 1004788
rect 125744 1004776 125750 1004828
rect 148778 1004776 148784 1004828
rect 148836 1004816 148842 1004828
rect 152918 1004816 152924 1004828
rect 148836 1004788 152924 1004816
rect 148836 1004776 148842 1004788
rect 152918 1004776 152924 1004788
rect 152976 1004776 152982 1004828
rect 156966 1004776 156972 1004828
rect 157024 1004816 157030 1004828
rect 174078 1004816 174084 1004828
rect 157024 1004788 174084 1004816
rect 157024 1004776 157030 1004788
rect 174078 1004776 174084 1004788
rect 174136 1004776 174142 1004828
rect 195698 1004776 195704 1004828
rect 195756 1004816 195762 1004828
rect 206370 1004816 206376 1004828
rect 195756 1004788 206376 1004816
rect 195756 1004776 195762 1004788
rect 206370 1004776 206376 1004788
rect 206428 1004776 206434 1004828
rect 215664 1004816 215692 1004856
rect 261018 1004844 261024 1004896
rect 261076 1004884 261082 1004896
rect 265066 1004884 265072 1004896
rect 261076 1004856 265072 1004884
rect 261076 1004844 261082 1004856
rect 265066 1004844 265072 1004856
rect 265124 1004844 265130 1004896
rect 357342 1004844 357348 1004896
rect 357400 1004884 357406 1004896
rect 362494 1004884 362500 1004896
rect 357400 1004856 362500 1004884
rect 357400 1004844 357406 1004856
rect 362494 1004844 362500 1004856
rect 362552 1004844 362558 1004896
rect 427170 1004844 427176 1004896
rect 427228 1004884 427234 1004896
rect 455414 1004884 455420 1004896
rect 427228 1004856 455420 1004884
rect 427228 1004844 427234 1004856
rect 455414 1004844 455420 1004856
rect 455472 1004844 455478 1004896
rect 553118 1004844 553124 1004896
rect 553176 1004884 553182 1004896
rect 555510 1004884 555516 1004896
rect 553176 1004856 555516 1004884
rect 553176 1004844 553182 1004856
rect 555510 1004844 555516 1004856
rect 555568 1004844 555574 1004896
rect 571242 1004884 571248 1004896
rect 557368 1004856 571248 1004884
rect 227898 1004816 227904 1004828
rect 215664 1004788 227904 1004816
rect 227898 1004776 227904 1004788
rect 227956 1004776 227962 1004828
rect 262214 1004776 262220 1004828
rect 262272 1004816 262278 1004828
rect 280246 1004816 280252 1004828
rect 262272 1004788 280252 1004816
rect 262272 1004776 262278 1004788
rect 280246 1004776 280252 1004788
rect 280304 1004776 280310 1004828
rect 357710 1004776 357716 1004828
rect 357768 1004816 357774 1004828
rect 364242 1004816 364248 1004828
rect 357768 1004788 364248 1004816
rect 357768 1004776 357774 1004788
rect 364242 1004776 364248 1004788
rect 364300 1004776 364306 1004828
rect 427538 1004776 427544 1004828
rect 427596 1004816 427602 1004828
rect 466546 1004816 466552 1004828
rect 427596 1004788 466552 1004816
rect 427596 1004776 427602 1004788
rect 466546 1004776 466552 1004788
rect 466604 1004776 466610 1004828
rect 500494 1004776 500500 1004828
rect 500552 1004816 500558 1004828
rect 509326 1004816 509332 1004828
rect 500552 1004788 509332 1004816
rect 500552 1004776 500558 1004788
rect 509326 1004776 509332 1004788
rect 509384 1004776 509390 1004828
rect 553946 1004776 553952 1004828
rect 554004 1004816 554010 1004828
rect 555694 1004816 555700 1004828
rect 554004 1004788 555700 1004816
rect 554004 1004776 554010 1004788
rect 555694 1004776 555700 1004788
rect 555752 1004776 555758 1004828
rect 93012 1004720 102134 1004748
rect 93012 1004708 93018 1004720
rect 105630 1004708 105636 1004760
rect 105688 1004748 105694 1004760
rect 125778 1004748 125784 1004760
rect 105688 1004720 125784 1004748
rect 105688 1004708 105694 1004720
rect 125778 1004708 125784 1004720
rect 125836 1004708 125842 1004760
rect 148870 1004708 148876 1004760
rect 148928 1004748 148934 1004760
rect 151722 1004748 151728 1004760
rect 148928 1004720 151728 1004748
rect 148928 1004708 148934 1004720
rect 151722 1004708 151728 1004720
rect 151780 1004708 151786 1004760
rect 157794 1004708 157800 1004760
rect 157852 1004748 157858 1004760
rect 173986 1004748 173992 1004760
rect 157852 1004720 173992 1004748
rect 157852 1004708 157858 1004720
rect 173986 1004708 173992 1004720
rect 174044 1004708 174050 1004760
rect 201034 1004708 201040 1004760
rect 201092 1004748 201098 1004760
rect 201862 1004748 201868 1004760
rect 201092 1004720 201868 1004748
rect 201092 1004708 201098 1004720
rect 201862 1004708 201868 1004720
rect 201920 1004708 201926 1004760
rect 261478 1004708 261484 1004760
rect 261536 1004748 261542 1004760
rect 265158 1004748 265164 1004760
rect 261536 1004720 265164 1004748
rect 261536 1004708 261542 1004720
rect 265158 1004708 265164 1004720
rect 265216 1004708 265222 1004760
rect 360562 1004708 360568 1004760
rect 360620 1004748 360626 1004760
rect 366358 1004748 366364 1004760
rect 360620 1004720 366364 1004748
rect 360620 1004708 360626 1004720
rect 366358 1004708 366364 1004720
rect 366416 1004708 366422 1004760
rect 419074 1004708 419080 1004760
rect 419132 1004748 419138 1004760
rect 421834 1004748 421840 1004760
rect 419132 1004720 421840 1004748
rect 419132 1004708 419138 1004720
rect 421834 1004708 421840 1004720
rect 421892 1004748 421898 1004760
rect 422662 1004748 422668 1004760
rect 421892 1004720 422668 1004748
rect 421892 1004708 421898 1004720
rect 422662 1004708 422668 1004720
rect 422720 1004708 422726 1004760
rect 425146 1004708 425152 1004760
rect 425204 1004748 425210 1004760
rect 467742 1004748 467748 1004760
rect 425204 1004720 467748 1004748
rect 425204 1004708 425210 1004720
rect 467742 1004708 467748 1004720
rect 467800 1004708 467806 1004760
rect 496630 1004708 496636 1004760
rect 496688 1004748 496694 1004760
rect 498838 1004748 498844 1004760
rect 496688 1004720 498844 1004748
rect 496688 1004708 496694 1004720
rect 498838 1004708 498844 1004720
rect 498896 1004748 498902 1004760
rect 499666 1004748 499672 1004760
rect 498896 1004720 499672 1004748
rect 498896 1004708 498902 1004720
rect 499666 1004708 499672 1004720
rect 499724 1004708 499730 1004760
rect 501690 1004708 501696 1004760
rect 501748 1004748 501754 1004760
rect 509234 1004748 509240 1004760
rect 501748 1004720 509240 1004748
rect 501748 1004708 501754 1004720
rect 509234 1004708 509240 1004720
rect 509292 1004708 509298 1004760
rect 549438 1004708 549444 1004760
rect 549496 1004748 549502 1004760
rect 550266 1004748 550272 1004760
rect 549496 1004720 550272 1004748
rect 549496 1004708 549502 1004720
rect 550266 1004708 550272 1004720
rect 550324 1004748 550330 1004760
rect 551094 1004748 551100 1004760
rect 550324 1004720 551100 1004748
rect 550324 1004708 550330 1004720
rect 551094 1004708 551100 1004720
rect 551152 1004708 551158 1004760
rect 552750 1004708 552756 1004760
rect 552808 1004748 552814 1004760
rect 557368 1004748 557396 1004856
rect 571242 1004844 571248 1004856
rect 571300 1004844 571306 1004896
rect 552808 1004720 557396 1004748
rect 552808 1004708 552814 1004720
rect 98270 1004640 98276 1004692
rect 98328 1004680 98334 1004692
rect 99098 1004680 99104 1004692
rect 98328 1004652 99104 1004680
rect 98328 1004640 98334 1004652
rect 99098 1004640 99104 1004652
rect 99156 1004680 99162 1004692
rect 125502 1004680 125508 1004692
rect 99156 1004652 125508 1004680
rect 99156 1004640 99162 1004652
rect 125502 1004640 125508 1004652
rect 125560 1004640 125566 1004692
rect 148962 1004640 148968 1004692
rect 149020 1004680 149026 1004692
rect 152550 1004680 152556 1004692
rect 149020 1004652 152556 1004680
rect 149020 1004640 149026 1004652
rect 152550 1004640 152556 1004652
rect 152608 1004640 152614 1004692
rect 154482 1004640 154488 1004692
rect 154540 1004680 154546 1004692
rect 160646 1004680 160652 1004692
rect 154540 1004652 160652 1004680
rect 154540 1004640 154546 1004652
rect 160646 1004640 160652 1004652
rect 160704 1004640 160710 1004692
rect 195146 1004640 195152 1004692
rect 195204 1004680 195210 1004692
rect 205910 1004680 205916 1004692
rect 195204 1004652 205916 1004680
rect 195204 1004640 195210 1004652
rect 205910 1004640 205916 1004652
rect 205968 1004640 205974 1004692
rect 252462 1004640 252468 1004692
rect 252520 1004680 252526 1004692
rect 253290 1004680 253296 1004692
rect 252520 1004652 253296 1004680
rect 252520 1004640 252526 1004652
rect 253290 1004640 253296 1004652
rect 253348 1004680 253354 1004692
rect 280062 1004680 280068 1004692
rect 253348 1004652 280068 1004680
rect 253348 1004640 253354 1004652
rect 280062 1004640 280068 1004652
rect 280120 1004640 280126 1004692
rect 315114 1004640 315120 1004692
rect 315172 1004680 315178 1004692
rect 331214 1004680 331220 1004692
rect 315172 1004652 331220 1004680
rect 315172 1004640 315178 1004652
rect 331214 1004640 331220 1004652
rect 331272 1004640 331278 1004692
rect 361390 1004640 361396 1004692
rect 361448 1004680 361454 1004692
rect 365438 1004680 365444 1004692
rect 361448 1004652 365444 1004680
rect 361448 1004640 361454 1004652
rect 365438 1004640 365444 1004652
rect 365496 1004640 365502 1004692
rect 366726 1004640 366732 1004692
rect 366784 1004680 366790 1004692
rect 383276 1004680 383282 1004692
rect 366784 1004652 383282 1004680
rect 366784 1004640 366790 1004652
rect 383276 1004640 383282 1004652
rect 383334 1004640 383340 1004692
rect 466454 1004640 466460 1004692
rect 466512 1004680 466518 1004692
rect 472250 1004680 472256 1004692
rect 466512 1004652 472256 1004680
rect 466512 1004640 466518 1004652
rect 472250 1004640 472256 1004652
rect 472308 1004640 472314 1004692
rect 502150 1004640 502156 1004692
rect 502208 1004680 502214 1004692
rect 509142 1004680 509148 1004692
rect 502208 1004652 509148 1004680
rect 502208 1004640 502214 1004652
rect 509142 1004640 509148 1004652
rect 509200 1004640 509206 1004692
rect 517330 1004640 517336 1004692
rect 517388 1004680 517394 1004692
rect 523586 1004680 523592 1004692
rect 517388 1004652 523592 1004680
rect 517388 1004640 517394 1004652
rect 523586 1004640 523592 1004652
rect 523644 1004640 523650 1004692
rect 555694 1004164 555700 1004216
rect 555752 1004204 555758 1004216
rect 569862 1004204 569868 1004216
rect 555752 1004176 569868 1004204
rect 555752 1004164 555758 1004176
rect 569862 1004164 569868 1004176
rect 569920 1004164 569926 1004216
rect 555510 1003892 555516 1003944
rect 555568 1003932 555574 1003944
rect 569954 1003932 569960 1003944
rect 555568 1003904 569960 1003932
rect 555568 1003892 555574 1003904
rect 569954 1003892 569960 1003904
rect 570012 1003892 570018 1003944
rect 553486 1003484 553492 1003536
rect 553544 1003524 553550 1003536
rect 556154 1003524 556160 1003536
rect 553544 1003496 556160 1003524
rect 553544 1003484 553550 1003496
rect 556154 1003484 556160 1003496
rect 556212 1003484 556218 1003536
rect 455414 1003280 455420 1003332
rect 455472 1003320 455478 1003332
rect 469030 1003320 469036 1003332
rect 455472 1003292 469036 1003320
rect 455472 1003280 455478 1003292
rect 469030 1003280 469036 1003292
rect 469088 1003280 469094 1003332
rect 554682 1003280 554688 1003332
rect 554740 1003320 554746 1003332
rect 571610 1003320 571616 1003332
rect 554740 1003292 571616 1003320
rect 554740 1003280 554746 1003292
rect 571610 1003280 571616 1003292
rect 571668 1003280 571674 1003332
rect 455506 1003212 455512 1003264
rect 455564 1003252 455570 1003264
rect 469122 1003252 469128 1003264
rect 455564 1003224 469128 1003252
rect 455564 1003212 455570 1003224
rect 469122 1003212 469128 1003224
rect 469180 1003212 469186 1003264
rect 554314 1003212 554320 1003264
rect 554372 1003252 554378 1003264
rect 571426 1003252 571432 1003264
rect 554372 1003224 571432 1003252
rect 554372 1003212 554378 1003224
rect 571426 1003212 571432 1003224
rect 571484 1003212 571490 1003264
rect 568574 1002056 568580 1002108
rect 568632 1002096 568638 1002108
rect 571518 1002096 571524 1002108
rect 568632 1002068 571524 1002096
rect 568632 1002056 568638 1002068
rect 571518 1002056 571524 1002068
rect 571576 1002056 571582 1002108
rect 440142 1001988 440148 1002040
rect 440200 1002028 440206 1002040
rect 440200 1002000 444512 1002028
rect 440200 1001988 440206 1002000
rect 440418 1001920 440424 1001972
rect 440476 1001960 440482 1001972
rect 444484 1001960 444512 1002000
rect 440476 1001932 444420 1001960
rect 444484 1001932 447272 1001960
rect 440476 1001920 440482 1001932
rect 143902 1001852 143908 1001904
rect 143960 1001892 143966 1001904
rect 148778 1001892 148784 1001904
rect 143960 1001864 148784 1001892
rect 143960 1001852 143966 1001864
rect 148778 1001852 148784 1001864
rect 148836 1001852 148842 1001904
rect 362494 1001852 362500 1001904
rect 362552 1001892 362558 1001904
rect 364426 1001892 364432 1001904
rect 362552 1001864 364432 1001892
rect 362552 1001852 362558 1001864
rect 364426 1001852 364432 1001864
rect 364484 1001852 364490 1001904
rect 444392 1001892 444420 1001932
rect 447134 1001892 447140 1001904
rect 444392 1001864 447140 1001892
rect 447134 1001852 447140 1001864
rect 447192 1001852 447198 1001904
rect 447244 1001892 447272 1001932
rect 466546 1001920 466552 1001972
rect 466604 1001960 466610 1001972
rect 472618 1001960 472624 1001972
rect 466604 1001932 472624 1001960
rect 466604 1001920 466610 1001932
rect 472618 1001920 472624 1001932
rect 472676 1001920 472682 1001972
rect 519170 1001920 519176 1001972
rect 519228 1001960 519234 1001972
rect 523770 1001960 523776 1001972
rect 519228 1001932 523776 1001960
rect 519228 1001920 519234 1001932
rect 523770 1001920 523776 1001932
rect 523828 1001920 523834 1001972
rect 590654 1001920 590660 1001972
rect 590712 1001960 590718 1001972
rect 625798 1001960 625804 1001972
rect 590712 1001932 625804 1001960
rect 590712 1001920 590718 1001932
rect 625798 1001920 625804 1001932
rect 625856 1001920 625862 1001972
rect 447318 1001892 447324 1001904
rect 447244 1001864 447324 1001892
rect 447318 1001852 447324 1001864
rect 447376 1001852 447382 1001904
rect 377306 1001716 377312 1001768
rect 377364 1001756 377370 1001768
rect 378318 1001756 378324 1001768
rect 377364 1001728 378324 1001756
rect 377364 1001716 377370 1001728
rect 378318 1001716 378324 1001728
rect 378376 1001716 378382 1001768
rect 556154 1001240 556160 1001292
rect 556212 1001280 556218 1001292
rect 571242 1001280 571248 1001292
rect 556212 1001252 571248 1001280
rect 556212 1001240 556218 1001252
rect 571242 1001240 571248 1001252
rect 571300 1001240 571306 1001292
rect 366358 1000764 366364 1000816
rect 366416 1000804 366422 1000816
rect 383552 1000804 383558 1000816
rect 366416 1000776 383558 1000804
rect 366416 1000764 366422 1000776
rect 383552 1000764 383558 1000776
rect 383610 1000764 383616 1000816
rect 455598 1000696 455604 1000748
rect 455656 1000736 455662 1000748
rect 472158 1000736 472164 1000748
rect 455656 1000708 472164 1000736
rect 455656 1000696 455662 1000708
rect 472158 1000696 472164 1000708
rect 472216 1000696 472222 1000748
rect 365438 1000628 365444 1000680
rect 365496 1000668 365502 1000680
rect 383368 1000668 383374 1000680
rect 365496 1000640 383374 1000668
rect 365496 1000628 365502 1000640
rect 383368 1000628 383374 1000640
rect 383426 1000628 383432 1000680
rect 427998 1000628 428004 1000680
rect 428056 1000668 428062 1000680
rect 472618 1000668 472624 1000680
rect 428056 1000640 472624 1000668
rect 428056 1000628 428062 1000640
rect 472618 1000628 472624 1000640
rect 472676 1000628 472682 1000680
rect 370406 1000560 370412 1000612
rect 370464 1000600 370470 1000612
rect 383460 1000600 383466 1000612
rect 370464 1000572 383466 1000600
rect 370464 1000560 370470 1000572
rect 383460 1000560 383466 1000572
rect 383518 1000560 383524 1000612
rect 426342 1000560 426348 1000612
rect 426400 1000600 426406 1000612
rect 472526 1000600 472532 1000612
rect 426400 1000572 472532 1000600
rect 426400 1000560 426406 1000572
rect 472526 1000560 472532 1000572
rect 472584 1000560 472590 1000612
rect 358906 1000492 358912 1000544
rect 358964 1000532 358970 1000544
rect 383552 1000532 383558 1000544
rect 358964 1000504 383558 1000532
rect 358964 1000492 358970 1000504
rect 383552 1000492 383558 1000504
rect 383610 1000492 383616 1000544
rect 425974 1000492 425980 1000544
rect 426032 1000532 426038 1000544
rect 472342 1000532 472348 1000544
rect 426032 1000504 472348 1000532
rect 426032 1000492 426038 1000504
rect 472342 1000492 472348 1000504
rect 472400 1000492 472406 1000544
rect 374270 1000424 374276 1000476
rect 374328 1000464 374334 1000476
rect 380986 1000464 380992 1000476
rect 374328 1000436 380992 1000464
rect 374328 1000424 374334 1000436
rect 380986 1000424 380992 1000436
rect 381044 1000424 381050 1000476
rect 380894 1000356 380900 1000408
rect 380952 1000396 380958 1000408
rect 383552 1000396 383558 1000408
rect 380952 1000368 383558 1000396
rect 380952 1000356 380958 1000368
rect 383552 1000356 383558 1000368
rect 383610 1000356 383616 1000408
rect 555970 1000016 555976 1000068
rect 556028 1000056 556034 1000068
rect 567010 1000056 567016 1000068
rect 556028 1000028 567016 1000056
rect 556028 1000016 556034 1000028
rect 567010 1000016 567016 1000028
rect 567068 1000016 567074 1000068
rect 564250 999988 564256 1000000
rect 554746 999960 564256 999988
rect 92402 999880 92408 999932
rect 92460 999920 92466 999932
rect 118694 999920 118700 999932
rect 92460 999892 118700 999920
rect 92460 999880 92466 999892
rect 118694 999880 118700 999892
rect 118752 999880 118758 999932
rect 246758 999880 246764 999932
rect 246816 999920 246822 999932
rect 258626 999920 258632 999932
rect 246816 999892 258632 999920
rect 246816 999880 246822 999892
rect 258626 999880 258632 999892
rect 258684 999880 258690 999932
rect 92586 999812 92592 999864
rect 92644 999852 92650 999864
rect 104342 999852 104348 999864
rect 92644 999824 104348 999852
rect 92644 999812 92650 999824
rect 104342 999812 104348 999824
rect 104400 999812 104406 999864
rect 246666 999812 246672 999864
rect 246724 999852 246730 999864
rect 257338 999852 257344 999864
rect 246724 999824 257344 999852
rect 246724 999812 246730 999824
rect 257338 999812 257344 999824
rect 257396 999812 257402 999864
rect 312170 999812 312176 999864
rect 312228 999852 312234 999864
rect 318886 999852 318892 999864
rect 312228 999824 318892 999852
rect 312228 999812 312234 999824
rect 318886 999812 318892 999824
rect 318944 999812 318950 999864
rect 430850 999812 430856 999864
rect 430908 999852 430914 999864
rect 439818 999852 439824 999864
rect 430908 999824 439824 999852
rect 430908 999812 430914 999824
rect 439818 999812 439824 999824
rect 439876 999812 439882 999864
rect 93046 999744 93052 999796
rect 93104 999784 93110 999796
rect 102778 999784 102784 999796
rect 93104 999756 102784 999784
rect 93104 999744 93110 999756
rect 102778 999744 102784 999756
rect 102836 999744 102842 999796
rect 246574 999744 246580 999796
rect 246632 999784 246638 999796
rect 256970 999784 256976 999796
rect 246632 999756 256976 999784
rect 246632 999744 246638 999756
rect 256970 999744 256976 999756
rect 257028 999744 257034 999796
rect 310146 999744 310152 999796
rect 310204 999784 310210 999796
rect 314930 999784 314936 999796
rect 310204 999756 314936 999784
rect 310204 999744 310210 999756
rect 314930 999744 314936 999756
rect 314988 999744 314994 999796
rect 431678 999744 431684 999796
rect 431736 999784 431742 999796
rect 437934 999784 437940 999796
rect 431736 999756 437940 999784
rect 431736 999744 431742 999756
rect 437934 999744 437940 999756
rect 437992 999744 437998 999796
rect 508682 999744 508688 999796
rect 508740 999784 508746 999796
rect 515214 999784 515220 999796
rect 508740 999756 515220 999784
rect 508740 999744 508746 999756
rect 515214 999744 515220 999756
rect 515272 999744 515278 999796
rect 92310 999676 92316 999728
rect 92368 999716 92374 999728
rect 100662 999716 100668 999728
rect 92368 999688 100668 999716
rect 92368 999676 92374 999688
rect 100662 999676 100668 999688
rect 100720 999676 100726 999728
rect 195422 999676 195428 999728
rect 195480 999716 195486 999728
rect 205542 999716 205548 999728
rect 195480 999688 205548 999716
rect 195480 999676 195486 999688
rect 205542 999676 205548 999688
rect 205600 999676 205606 999728
rect 246850 999676 246856 999728
rect 246908 999716 246914 999728
rect 257798 999716 257804 999728
rect 246908 999688 257804 999716
rect 246908 999676 246914 999688
rect 257798 999676 257804 999688
rect 257856 999676 257862 999728
rect 311434 999676 311440 999728
rect 311492 999716 311498 999728
rect 315942 999716 315948 999728
rect 311492 999688 315948 999716
rect 311492 999676 311498 999688
rect 315942 999676 315948 999688
rect 316000 999676 316006 999728
rect 361850 999676 361856 999728
rect 361908 999716 361914 999728
rect 368750 999716 368756 999728
rect 361908 999688 368756 999716
rect 361908 999676 361914 999688
rect 368750 999676 368756 999688
rect 368808 999676 368814 999728
rect 429194 999676 429200 999728
rect 429252 999716 429258 999728
rect 434622 999716 434628 999728
rect 429252 999688 434628 999716
rect 429252 999676 429258 999688
rect 434622 999676 434628 999688
rect 434680 999676 434686 999728
rect 506198 999676 506204 999728
rect 506256 999716 506262 999728
rect 512086 999716 512092 999728
rect 506256 999688 512092 999716
rect 506256 999676 506262 999688
rect 512086 999676 512092 999688
rect 512144 999676 512150 999728
rect 92862 999608 92868 999660
rect 92920 999648 92926 999660
rect 102318 999648 102324 999660
rect 92920 999620 102324 999648
rect 92920 999608 92926 999620
rect 102318 999608 102324 999620
rect 102376 999608 102382 999660
rect 195514 999608 195520 999660
rect 195572 999648 195578 999660
rect 203886 999648 203892 999660
rect 195572 999620 203892 999648
rect 195572 999608 195578 999620
rect 203886 999608 203892 999620
rect 203944 999608 203950 999660
rect 249702 999608 249708 999660
rect 249760 999648 249766 999660
rect 254854 999648 254860 999660
rect 249760 999620 254860 999648
rect 249760 999608 249766 999620
rect 254854 999608 254860 999620
rect 254912 999608 254918 999660
rect 313826 999608 313832 999660
rect 313884 999648 313890 999660
rect 318702 999648 318708 999660
rect 313884 999620 318708 999648
rect 313884 999608 313890 999620
rect 318702 999608 318708 999620
rect 318760 999608 318766 999660
rect 362586 999608 362592 999660
rect 362644 999648 362650 999660
rect 368566 999648 368572 999660
rect 362644 999620 368572 999648
rect 362644 999608 362650 999620
rect 368566 999608 368572 999620
rect 368624 999608 368630 999660
rect 430022 999608 430028 999660
rect 430080 999648 430086 999660
rect 434806 999648 434812 999660
rect 430080 999620 434812 999648
rect 430080 999608 430086 999620
rect 434806 999608 434812 999620
rect 434864 999608 434870 999660
rect 508222 999608 508228 999660
rect 508280 999648 508286 999660
rect 513466 999648 513472 999660
rect 508280 999620 513472 999648
rect 508280 999608 508286 999620
rect 513466 999608 513472 999620
rect 513524 999608 513530 999660
rect 92770 999540 92776 999592
rect 92828 999580 92834 999592
rect 101950 999580 101956 999592
rect 92828 999552 101956 999580
rect 92828 999540 92834 999552
rect 101950 999540 101956 999552
rect 102008 999540 102014 999592
rect 155770 999540 155776 999592
rect 155828 999580 155834 999592
rect 160278 999580 160284 999592
rect 155828 999552 160284 999580
rect 155828 999540 155834 999552
rect 160278 999540 160284 999552
rect 160336 999540 160342 999592
rect 195606 999540 195612 999592
rect 195664 999580 195670 999592
rect 203518 999580 203524 999592
rect 195664 999552 203524 999580
rect 195664 999540 195670 999552
rect 203518 999540 203524 999552
rect 203576 999540 203582 999592
rect 250438 999540 250444 999592
rect 250496 999580 250502 999592
rect 256142 999580 256148 999592
rect 250496 999552 256148 999580
rect 250496 999540 250502 999552
rect 256142 999540 256148 999552
rect 256200 999540 256206 999592
rect 312630 999540 312636 999592
rect 312688 999580 312694 999592
rect 315114 999580 315120 999592
rect 312688 999552 315120 999580
rect 312688 999540 312694 999552
rect 315114 999540 315120 999552
rect 315172 999540 315178 999592
rect 363414 999540 363420 999592
rect 363472 999580 363478 999592
rect 368934 999580 368940 999592
rect 363472 999552 368940 999580
rect 363472 999540 363478 999552
rect 368934 999540 368940 999552
rect 368992 999540 368998 999592
rect 431218 999540 431224 999592
rect 431276 999580 431282 999592
rect 436186 999580 436192 999592
rect 431276 999552 436192 999580
rect 431276 999540 431282 999552
rect 436186 999540 436192 999552
rect 436244 999540 436250 999592
rect 507026 999540 507032 999592
rect 507084 999580 507090 999592
rect 511902 999580 511908 999592
rect 507084 999552 511908 999580
rect 507084 999540 507090 999552
rect 511902 999540 511908 999552
rect 511960 999540 511966 999592
rect 95142 999472 95148 999524
rect 95200 999512 95206 999524
rect 101490 999512 101496 999524
rect 95200 999484 101496 999512
rect 95200 999472 95206 999484
rect 101490 999472 101496 999484
rect 101548 999472 101554 999524
rect 159082 999472 159088 999524
rect 159140 999512 159146 999524
rect 162854 999512 162860 999524
rect 159140 999484 162860 999512
rect 159140 999472 159146 999484
rect 162854 999472 162860 999484
rect 162912 999472 162918 999524
rect 198458 999472 198464 999524
rect 198516 999512 198522 999524
rect 204346 999512 204352 999524
rect 198516 999484 204352 999512
rect 198516 999472 198522 999484
rect 204346 999472 204352 999484
rect 204404 999472 204410 999524
rect 250254 999472 250260 999524
rect 250312 999512 250318 999524
rect 255682 999512 255688 999524
rect 250312 999484 255688 999512
rect 250312 999472 250318 999484
rect 255682 999472 255688 999484
rect 255740 999472 255746 999524
rect 314838 999472 314844 999524
rect 314896 999512 314902 999524
rect 319070 999512 319076 999524
rect 314896 999484 319076 999512
rect 314896 999472 314902 999484
rect 319070 999472 319076 999484
rect 319128 999472 319134 999524
rect 365070 999472 365076 999524
rect 365128 999512 365134 999524
rect 371510 999512 371516 999524
rect 365128 999484 371516 999512
rect 365128 999472 365134 999484
rect 371510 999472 371516 999484
rect 371568 999472 371574 999524
rect 432414 999472 432420 999524
rect 432472 999512 432478 999524
rect 437566 999512 437572 999524
rect 432472 999484 437572 999512
rect 432472 999472 432478 999484
rect 437566 999472 437572 999484
rect 437624 999472 437630 999524
rect 507854 999472 507860 999524
rect 507912 999512 507918 999524
rect 512270 999512 512276 999524
rect 507912 999484 512276 999512
rect 507912 999472 507918 999484
rect 512270 999472 512276 999484
rect 512328 999472 512334 999524
rect 97902 999404 97908 999456
rect 97960 999444 97966 999456
rect 103146 999444 103152 999456
rect 97960 999416 103152 999444
rect 97960 999404 97966 999416
rect 103146 999404 103152 999416
rect 103204 999404 103210 999456
rect 198366 999404 198372 999456
rect 198424 999444 198430 999456
rect 204714 999444 204720 999456
rect 198424 999416 204720 999444
rect 198424 999404 198430 999416
rect 204714 999404 204720 999416
rect 204772 999404 204778 999456
rect 208854 999404 208860 999456
rect 208912 999444 208918 999456
rect 212718 999444 212724 999456
rect 208912 999416 212724 999444
rect 208912 999404 208918 999416
rect 212718 999404 212724 999416
rect 212776 999404 212782 999456
rect 250070 999404 250076 999456
rect 250128 999444 250134 999456
rect 255314 999444 255320 999456
rect 250128 999416 255320 999444
rect 250128 999404 250134 999416
rect 255314 999404 255320 999416
rect 255372 999404 255378 999456
rect 362218 999404 362224 999456
rect 362276 999444 362282 999456
rect 367186 999444 367192 999456
rect 362276 999416 367192 999444
rect 362276 999404 362282 999416
rect 367186 999404 367192 999416
rect 367244 999404 367250 999456
rect 432874 999404 432880 999456
rect 432932 999444 432938 999456
rect 437750 999444 437756 999456
rect 432932 999416 437756 999444
rect 432932 999404 432938 999416
rect 437750 999404 437756 999416
rect 437808 999404 437814 999456
rect 506658 999404 506664 999456
rect 506716 999444 506722 999456
rect 510706 999444 510712 999456
rect 506716 999416 510712 999444
rect 506716 999404 506722 999416
rect 510706 999404 510712 999416
rect 510764 999404 510770 999456
rect 92678 999336 92684 999388
rect 92736 999376 92742 999388
rect 99466 999376 99472 999388
rect 92736 999348 99472 999376
rect 92736 999336 92742 999348
rect 99466 999336 99472 999348
rect 99524 999336 99530 999388
rect 195238 999336 195244 999388
rect 195296 999376 195302 999388
rect 202230 999376 202236 999388
rect 195296 999348 202236 999376
rect 195296 999336 195302 999348
rect 202230 999336 202236 999348
rect 202288 999336 202294 999388
rect 210418 999336 210424 999388
rect 210476 999376 210482 999388
rect 218966 999376 218972 999388
rect 210476 999348 218972 999376
rect 210476 999336 210482 999348
rect 218966 999336 218972 999348
rect 219024 999336 219030 999388
rect 246942 999336 246948 999388
rect 247000 999376 247006 999388
rect 253658 999376 253664 999388
rect 247000 999348 253664 999376
rect 247000 999336 247006 999348
rect 253658 999336 253664 999348
rect 253716 999336 253722 999388
rect 364702 999336 364708 999388
rect 364760 999376 364766 999388
rect 369854 999376 369860 999388
rect 364760 999348 369860 999376
rect 364760 999336 364766 999348
rect 369854 999336 369860 999348
rect 369912 999336 369918 999388
rect 429654 999336 429660 999388
rect 429712 999376 429718 999388
rect 433334 999376 433340 999388
rect 429712 999348 433340 999376
rect 429712 999336 429718 999348
rect 433334 999336 433340 999348
rect 433392 999336 433398 999388
rect 509050 999336 509056 999388
rect 509108 999376 509114 999388
rect 513374 999376 513380 999388
rect 509108 999348 513380 999376
rect 509108 999336 509114 999348
rect 513374 999336 513380 999348
rect 513432 999336 513438 999388
rect 95694 999268 95700 999320
rect 95752 999308 95758 999320
rect 101122 999308 101128 999320
rect 95752 999280 101128 999308
rect 95752 999268 95758 999280
rect 101122 999268 101128 999280
rect 101180 999268 101186 999320
rect 200114 999268 200120 999320
rect 200172 999308 200178 999320
rect 205174 999308 205180 999320
rect 200172 999280 205180 999308
rect 200172 999268 200178 999280
rect 205174 999268 205180 999280
rect 205232 999268 205238 999320
rect 209590 999268 209596 999320
rect 209648 999308 209654 999320
rect 212626 999308 212632 999320
rect 209648 999280 212632 999308
rect 209648 999268 209654 999280
rect 212626 999268 212632 999280
rect 212684 999268 212690 999320
rect 249886 999268 249892 999320
rect 249944 999308 249950 999320
rect 254486 999308 254492 999320
rect 249944 999280 254492 999308
rect 249944 999268 249950 999280
rect 254486 999268 254492 999280
rect 254544 999268 254550 999320
rect 365438 999268 365444 999320
rect 365496 999308 365502 999320
rect 371142 999308 371148 999320
rect 365496 999280 371148 999308
rect 365496 999268 365502 999280
rect 371142 999268 371148 999280
rect 371200 999268 371206 999320
rect 430390 999268 430396 999320
rect 430448 999308 430454 999320
rect 433426 999308 433432 999320
rect 430448 999280 433432 999308
rect 430448 999268 430454 999280
rect 433426 999268 433432 999280
rect 433484 999268 433490 999320
rect 507394 999268 507400 999320
rect 507452 999308 507458 999320
rect 510614 999308 510620 999320
rect 507452 999280 510620 999308
rect 507452 999268 507458 999280
rect 510614 999268 510620 999280
rect 510672 999268 510678 999320
rect 540330 999268 540336 999320
rect 540388 999308 540394 999320
rect 554746 999308 554774 999960
rect 564250 999948 564256 999960
rect 564308 999948 564314 1000000
rect 558454 999880 558460 999932
rect 558512 999920 558518 999932
rect 564526 999920 564532 999932
rect 558512 999892 564532 999920
rect 558512 999880 558518 999892
rect 564526 999880 564532 999892
rect 564584 999880 564590 999932
rect 560846 999812 560852 999864
rect 560904 999852 560910 999864
rect 567286 999852 567292 999864
rect 560904 999824 567292 999852
rect 560904 999812 560910 999824
rect 567286 999812 567292 999824
rect 567344 999812 567350 999864
rect 556338 999744 556344 999796
rect 556396 999784 556402 999796
rect 562134 999784 562140 999796
rect 556396 999756 562140 999784
rect 556396 999744 556402 999756
rect 562134 999744 562140 999756
rect 562192 999744 562198 999796
rect 560478 999676 560484 999728
rect 560536 999716 560542 999728
rect 565814 999716 565820 999728
rect 560536 999688 565820 999716
rect 560536 999676 560542 999688
rect 565814 999676 565820 999688
rect 565872 999676 565878 999728
rect 559190 999608 559196 999660
rect 559248 999648 559254 999660
rect 564342 999648 564348 999660
rect 559248 999620 564348 999648
rect 559248 999608 559254 999620
rect 564342 999608 564348 999620
rect 564400 999608 564406 999660
rect 560018 999540 560024 999592
rect 560076 999580 560082 999592
rect 564710 999580 564716 999592
rect 560076 999552 564716 999580
rect 560076 999540 560082 999552
rect 564710 999540 564716 999552
rect 564768 999540 564774 999592
rect 557994 999472 558000 999524
rect 558052 999512 558058 999524
rect 563054 999512 563060 999524
rect 558052 999484 563060 999512
rect 558052 999472 558058 999484
rect 563054 999472 563060 999484
rect 563112 999472 563118 999524
rect 556798 999404 556804 999456
rect 556856 999444 556862 999456
rect 561766 999444 561772 999456
rect 556856 999416 561772 999444
rect 556856 999404 556862 999416
rect 561766 999404 561772 999416
rect 561824 999404 561830 999456
rect 590746 999404 590752 999456
rect 590804 999444 590810 999456
rect 625430 999444 625436 999456
rect 590804 999416 625436 999444
rect 590804 999404 590810 999416
rect 625430 999404 625436 999416
rect 625488 999404 625494 999456
rect 557166 999336 557172 999388
rect 557224 999376 557230 999388
rect 561950 999376 561956 999388
rect 557224 999348 561956 999376
rect 557224 999336 557230 999348
rect 561950 999336 561956 999348
rect 562008 999336 562014 999388
rect 540388 999280 554774 999308
rect 540388 999268 540394 999280
rect 558822 999268 558828 999320
rect 558880 999308 558886 999320
rect 563146 999308 563152 999320
rect 558880 999280 563152 999308
rect 558880 999268 558886 999280
rect 563146 999268 563152 999280
rect 563204 999268 563210 999320
rect 607122 999268 607128 999320
rect 607180 999308 607186 999320
rect 625614 999308 625620 999320
rect 607180 999280 625620 999308
rect 607180 999268 607186 999280
rect 625614 999268 625620 999280
rect 625672 999268 625678 999320
rect 95326 999200 95332 999252
rect 95384 999240 95390 999252
rect 100294 999240 100300 999252
rect 95384 999212 100300 999240
rect 95384 999200 95390 999212
rect 100294 999200 100300 999212
rect 100352 999200 100358 999252
rect 198642 999200 198648 999252
rect 198700 999240 198706 999252
rect 202690 999240 202696 999252
rect 198700 999212 202696 999240
rect 198700 999200 198706 999212
rect 202690 999200 202696 999212
rect 202748 999200 202754 999252
rect 211706 999200 211712 999252
rect 211764 999240 211770 999252
rect 216582 999240 216588 999252
rect 211764 999212 216588 999240
rect 211764 999200 211770 999212
rect 216582 999200 216588 999212
rect 216640 999200 216646 999252
rect 252462 999200 252468 999252
rect 252520 999240 252526 999252
rect 256510 999240 256516 999252
rect 252520 999212 256516 999240
rect 252520 999200 252526 999212
rect 256510 999200 256516 999212
rect 256568 999200 256574 999252
rect 364242 999200 364248 999252
rect 364300 999240 364306 999252
rect 368382 999240 368388 999252
rect 364300 999212 368388 999240
rect 364300 999200 364306 999212
rect 368382 999200 368388 999212
rect 368440 999200 368446 999252
rect 432046 999200 432052 999252
rect 432104 999240 432110 999252
rect 436094 999240 436100 999252
rect 432104 999212 436100 999240
rect 432104 999200 432110 999212
rect 436094 999200 436100 999212
rect 436152 999200 436158 999252
rect 500862 999200 500868 999252
rect 500920 999240 500926 999252
rect 507854 999240 507860 999252
rect 500920 999212 507860 999240
rect 500920 999200 500926 999212
rect 507854 999200 507860 999212
rect 507912 999200 507918 999252
rect 509510 999200 509516 999252
rect 509568 999240 509574 999252
rect 514662 999240 514668 999252
rect 509568 999212 514668 999240
rect 509568 999200 509574 999212
rect 514662 999200 514668 999212
rect 514720 999200 514726 999252
rect 548886 999200 548892 999252
rect 548944 999240 548950 999252
rect 554314 999240 554320 999252
rect 548944 999212 554320 999240
rect 548944 999200 548950 999212
rect 554314 999200 554320 999212
rect 554372 999200 554378 999252
rect 559650 999200 559656 999252
rect 559708 999240 559714 999252
rect 563238 999240 563244 999252
rect 559708 999212 563244 999240
rect 559708 999200 559714 999212
rect 563238 999200 563244 999212
rect 563296 999200 563302 999252
rect 602246 999200 602252 999252
rect 602304 999240 602310 999252
rect 625706 999240 625712 999252
rect 602304 999212 625712 999240
rect 602304 999200 602310 999212
rect 625706 999200 625712 999212
rect 625764 999200 625770 999252
rect 92310 999132 92316 999184
rect 92368 999172 92374 999184
rect 93046 999172 93052 999184
rect 92368 999144 93052 999172
rect 92368 999132 92374 999144
rect 93046 999132 93052 999144
rect 93104 999132 93110 999184
rect 95510 999132 95516 999184
rect 95568 999172 95574 999184
rect 99926 999172 99932 999184
rect 95568 999144 99932 999172
rect 95568 999132 95574 999144
rect 99926 999132 99932 999144
rect 99984 999132 99990 999184
rect 143810 999132 143816 999184
rect 143868 999172 143874 999184
rect 148962 999172 148968 999184
rect 143868 999144 148968 999172
rect 143868 999132 143874 999144
rect 148962 999132 148968 999144
rect 149020 999132 149026 999184
rect 154114 999132 154120 999184
rect 154172 999172 154178 999184
rect 155770 999172 155776 999184
rect 154172 999144 155776 999172
rect 154172 999132 154178 999144
rect 155770 999132 155776 999144
rect 155828 999132 155834 999184
rect 198550 999132 198556 999184
rect 198608 999172 198614 999184
rect 203058 999172 203064 999184
rect 198608 999144 203064 999172
rect 198608 999132 198614 999144
rect 203058 999132 203064 999144
rect 203116 999132 203122 999184
rect 211246 999132 211252 999184
rect 211304 999172 211310 999184
rect 215294 999172 215300 999184
rect 211304 999144 215300 999172
rect 211304 999132 211310 999144
rect 215294 999132 215300 999144
rect 215352 999132 215358 999184
rect 250622 999132 250628 999184
rect 250680 999172 250686 999184
rect 254118 999172 254124 999184
rect 250680 999144 254124 999172
rect 250680 999132 250686 999144
rect 254118 999132 254124 999144
rect 254176 999132 254182 999184
rect 258534 999132 258540 999184
rect 258592 999172 258598 999184
rect 262214 999172 262220 999184
rect 258592 999144 262220 999172
rect 258592 999132 258598 999144
rect 262214 999132 262220 999144
rect 262272 999132 262278 999184
rect 355962 999132 355968 999184
rect 356020 999172 356026 999184
rect 358906 999172 358912 999184
rect 356020 999144 358912 999172
rect 356020 999132 356026 999144
rect 358906 999132 358912 999144
rect 358964 999132 358970 999184
rect 363046 999132 363052 999184
rect 363104 999172 363110 999184
rect 367094 999172 367100 999184
rect 363104 999144 367100 999172
rect 363104 999132 363110 999144
rect 367094 999132 367100 999144
rect 367152 999132 367158 999184
rect 378042 999132 378048 999184
rect 378100 999172 378106 999184
rect 383184 999172 383190 999184
rect 378100 999144 383190 999172
rect 378100 999132 378106 999144
rect 383184 999132 383190 999144
rect 383242 999132 383248 999184
rect 400030 999132 400036 999184
rect 400088 999172 400094 999184
rect 444374 999172 444380 999184
rect 400088 999144 444380 999172
rect 400088 999132 400094 999144
rect 444374 999132 444380 999144
rect 444432 999132 444438 999184
rect 464246 999132 464252 999184
rect 464304 999172 464310 999184
rect 472434 999172 472440 999184
rect 464304 999144 472440 999172
rect 464304 999132 464310 999144
rect 472434 999132 472440 999144
rect 472492 999132 472498 999184
rect 499482 999132 499488 999184
rect 499540 999172 499546 999184
rect 503346 999172 503352 999184
rect 499540 999144 503352 999172
rect 499540 999132 499546 999144
rect 503346 999132 503352 999144
rect 503404 999132 503410 999184
rect 509878 999132 509884 999184
rect 509936 999172 509942 999184
rect 514846 999172 514852 999184
rect 509936 999144 514852 999172
rect 509936 999132 509942 999144
rect 514846 999132 514852 999144
rect 514904 999132 514910 999184
rect 549070 999132 549076 999184
rect 549128 999172 549134 999184
rect 551922 999172 551928 999184
rect 549128 999144 551928 999172
rect 549128 999132 549134 999144
rect 551922 999132 551928 999144
rect 551980 999132 551986 999184
rect 557626 999132 557632 999184
rect 557684 999172 557690 999184
rect 561582 999172 561588 999184
rect 557684 999144 561588 999172
rect 557684 999132 557690 999144
rect 561582 999132 561588 999144
rect 561640 999132 561646 999184
rect 561674 999132 561680 999184
rect 561732 999172 561738 999184
rect 567102 999172 567108 999184
rect 561732 999144 567108 999172
rect 561732 999132 561738 999144
rect 567102 999132 567108 999144
rect 567160 999132 567166 999184
rect 612734 999132 612740 999184
rect 612792 999172 612798 999184
rect 625798 999172 625804 999184
rect 612792 999144 625804 999172
rect 612792 999132 612798 999144
rect 625798 999132 625804 999144
rect 625856 999132 625862 999184
rect 118694 999064 118700 999116
rect 118752 999104 118758 999116
rect 122098 999104 122104 999116
rect 118752 999076 122104 999104
rect 118752 999064 118758 999076
rect 122098 999064 122104 999076
rect 122156 999064 122162 999116
rect 143994 999064 144000 999116
rect 144052 999104 144058 999116
rect 158254 999104 158260 999116
rect 144052 999076 158260 999104
rect 144052 999064 144058 999076
rect 158254 999064 158260 999076
rect 158312 999064 158318 999116
rect 247954 999064 247960 999116
rect 248012 999104 248018 999116
rect 265158 999104 265164 999116
rect 248012 999076 265164 999104
rect 248012 999064 248018 999076
rect 265158 999064 265164 999076
rect 265216 999064 265222 999116
rect 298738 999064 298744 999116
rect 298796 999104 298802 999116
rect 312630 999104 312636 999116
rect 298796 999076 312636 999104
rect 298796 999064 298802 999076
rect 312630 999064 312636 999076
rect 312688 999064 312694 999116
rect 399938 999064 399944 999116
rect 399996 999104 400002 999116
rect 436186 999104 436192 999116
rect 399996 999076 436192 999104
rect 399996 999064 400002 999076
rect 436186 999064 436192 999076
rect 436244 999064 436250 999116
rect 453942 999064 453948 999116
rect 454000 999104 454006 999116
rect 462774 999104 462780 999116
rect 454000 999076 462780 999104
rect 454000 999064 454006 999076
rect 462774 999064 462780 999076
rect 462832 999064 462838 999116
rect 488902 999064 488908 999116
rect 488960 999104 488966 999116
rect 513466 999104 513472 999116
rect 488960 999076 513472 999104
rect 488960 999064 488966 999076
rect 513466 999064 513472 999076
rect 513524 999064 513530 999116
rect 509326 998996 509332 999048
rect 509384 999036 509390 999048
rect 521286 999036 521292 999048
rect 509384 999008 521292 999036
rect 509384 998996 509390 999008
rect 521286 998996 521292 999008
rect 521344 998996 521350 999048
rect 509234 998928 509240 998980
rect 509292 998968 509298 998980
rect 521470 998968 521476 998980
rect 509292 998940 521476 998968
rect 509292 998928 509298 998940
rect 521470 998928 521476 998940
rect 521528 998928 521534 998980
rect 509142 998860 509148 998912
rect 509200 998900 509206 998912
rect 521378 998900 521384 998912
rect 509200 998872 521384 998900
rect 509200 998860 509206 998872
rect 521378 998860 521384 998872
rect 521436 998860 521442 998912
rect 507854 998792 507860 998844
rect 507912 998832 507918 998844
rect 521562 998832 521568 998844
rect 507912 998804 521568 998832
rect 507912 998792 507918 998804
rect 521562 998792 521568 998804
rect 521620 998792 521626 998844
rect 467742 998316 467748 998368
rect 467800 998356 467806 998368
rect 470870 998356 470876 998368
rect 467800 998328 470876 998356
rect 467800 998316 467806 998328
rect 470870 998316 470876 998328
rect 470928 998316 470934 998368
rect 364334 998180 364340 998232
rect 364392 998220 364398 998232
rect 375190 998220 375196 998232
rect 364392 998192 375196 998220
rect 364392 998180 364398 998192
rect 375190 998180 375196 998192
rect 375248 998180 375254 998232
rect 467834 998112 467840 998164
rect 467892 998152 467898 998164
rect 469398 998152 469404 998164
rect 467892 998124 469404 998152
rect 467892 998112 467898 998124
rect 469398 998112 469404 998124
rect 469456 998112 469462 998164
rect 364426 997908 364432 997960
rect 364484 997948 364490 997960
rect 374454 997948 374460 997960
rect 364484 997920 374460 997948
rect 364484 997908 364490 997920
rect 374454 997908 374460 997920
rect 374512 997908 374518 997960
rect 549070 997772 549076 997824
rect 549128 997812 549134 997824
rect 575566 997812 575572 997824
rect 549128 997784 575572 997812
rect 549128 997772 549134 997784
rect 575566 997772 575572 997784
rect 575624 997772 575630 997824
rect 144086 997704 144092 997756
rect 144144 997744 144150 997756
rect 156138 997744 156144 997756
rect 144144 997716 156144 997744
rect 144144 997704 144150 997716
rect 156138 997704 156144 997716
rect 156196 997704 156202 997756
rect 571518 997704 571524 997756
rect 571576 997744 571582 997756
rect 623774 997744 623780 997756
rect 571576 997716 623780 997744
rect 571576 997704 571582 997716
rect 623774 997704 623780 997716
rect 623832 997704 623838 997756
rect 561950 997636 561956 997688
rect 562008 997676 562014 997688
rect 590654 997676 590660 997688
rect 562008 997648 590660 997676
rect 562008 997636 562014 997648
rect 590654 997636 590660 997648
rect 590712 997636 590718 997688
rect 548886 997568 548892 997620
rect 548944 997608 548950 997620
rect 612734 997608 612740 997620
rect 548944 997580 612740 997608
rect 548944 997568 548950 997580
rect 612734 997568 612740 997580
rect 612792 997568 612798 997620
rect 571334 997500 571340 997552
rect 571392 997540 571398 997552
rect 590746 997540 590752 997552
rect 571392 997512 590752 997540
rect 571392 997500 571398 997512
rect 590746 997500 590752 997512
rect 590804 997500 590810 997552
rect 569862 997432 569868 997484
rect 569920 997472 569926 997484
rect 607122 997472 607128 997484
rect 569920 997444 607128 997472
rect 569920 997432 569926 997444
rect 607122 997432 607128 997444
rect 607180 997432 607186 997484
rect 571426 997364 571432 997416
rect 571484 997404 571490 997416
rect 602246 997404 602252 997416
rect 571484 997376 602252 997404
rect 571484 997364 571490 997376
rect 602246 997364 602252 997376
rect 602304 997364 602310 997416
rect 562134 997296 562140 997348
rect 562192 997336 562198 997348
rect 623682 997336 623688 997348
rect 562192 997308 623688 997336
rect 562192 997296 562198 997308
rect 623682 997296 623688 997308
rect 623740 997296 623746 997348
rect 107654 997160 107660 997212
rect 107712 997200 107718 997212
rect 115934 997200 115940 997212
rect 107712 997172 115940 997200
rect 107712 997160 107718 997172
rect 115934 997160 115940 997172
rect 115992 997160 115998 997212
rect 143994 997092 144000 997144
rect 144052 997132 144058 997144
rect 147766 997132 147772 997144
rect 144052 997104 147772 997132
rect 144052 997092 144058 997104
rect 147766 997092 147772 997104
rect 147824 997092 147830 997144
rect 301774 996276 301780 996328
rect 301832 996316 301838 996328
rect 308122 996316 308128 996328
rect 301832 996288 308128 996316
rect 301832 996276 301838 996288
rect 308122 996276 308128 996288
rect 308180 996276 308186 996328
rect 300210 996208 300216 996260
rect 300268 996248 300274 996260
rect 305730 996248 305736 996260
rect 300268 996220 305736 996248
rect 300268 996208 300274 996220
rect 305730 996208 305736 996220
rect 305788 996208 305794 996260
rect 125594 996135 125600 996187
rect 125652 996175 125658 996187
rect 157794 996175 157800 996187
rect 125652 996147 157800 996175
rect 125652 996135 125658 996147
rect 157794 996135 157800 996147
rect 157852 996135 157858 996187
rect 173894 996135 173900 996187
rect 173952 996175 173958 996187
rect 215294 996175 215300 996187
rect 173952 996147 215300 996175
rect 173952 996135 173958 996147
rect 215294 996135 215300 996147
rect 215352 996135 215358 996187
rect 227898 996135 227904 996187
rect 227956 996175 227962 996187
rect 267826 996175 267832 996187
rect 227956 996147 267832 996175
rect 227956 996135 227962 996147
rect 267826 996135 267832 996147
rect 267884 996175 267890 996187
rect 270402 996175 270408 996187
rect 267884 996147 270408 996175
rect 267884 996135 267890 996147
rect 270402 996135 270408 996147
rect 270460 996135 270466 996187
rect 280246 996130 280252 996182
rect 280304 996170 280310 996182
rect 314286 996170 314292 996192
rect 280304 996142 314292 996170
rect 280304 996130 280310 996142
rect 314286 996140 314292 996142
rect 314344 996140 314350 996192
rect 512270 996130 512276 996182
rect 512328 996170 512334 996182
rect 563238 996170 563244 996182
rect 512328 996142 563244 996170
rect 512328 996130 512334 996142
rect 563238 996130 563244 996142
rect 563296 996130 563302 996182
rect 108482 996072 108488 996124
rect 108540 996112 108546 996124
rect 113358 996112 113364 996124
rect 108540 996084 113364 996112
rect 108540 996072 108546 996084
rect 113358 996072 113364 996084
rect 113416 996072 113422 996124
rect 125686 996067 125692 996119
rect 125744 996107 125750 996119
rect 159450 996107 159456 996119
rect 125744 996079 159456 996107
rect 125744 996067 125750 996079
rect 159450 996067 159456 996079
rect 159508 996067 159514 996119
rect 173986 996067 173992 996119
rect 174044 996107 174050 996119
rect 212626 996107 212632 996119
rect 174044 996079 212632 996107
rect 174044 996067 174050 996079
rect 212626 996067 212632 996079
rect 212684 996067 212690 996119
rect 227806 996067 227812 996119
rect 227864 996107 227870 996119
rect 265250 996107 265256 996119
rect 227864 996079 265256 996107
rect 227864 996067 227870 996079
rect 265250 996067 265256 996079
rect 265308 996107 265314 996119
rect 267642 996107 267648 996119
rect 265308 996079 267648 996107
rect 265308 996067 265314 996079
rect 267642 996067 267648 996079
rect 267700 996067 267706 996119
rect 280154 996062 280160 996114
rect 280212 996102 280218 996114
rect 315114 996102 315120 996124
rect 280212 996074 315120 996102
rect 280212 996062 280218 996074
rect 315114 996072 315120 996074
rect 315172 996112 315178 996124
rect 317506 996112 317512 996124
rect 315172 996084 317512 996112
rect 315172 996072 315178 996084
rect 317506 996072 317512 996084
rect 317564 996072 317570 996124
rect 125778 995999 125784 996051
rect 125836 996039 125842 996051
rect 156966 996039 156972 996051
rect 125836 996011 156972 996039
rect 125836 995999 125842 996011
rect 156966 995999 156972 996011
rect 157024 996039 157030 996051
rect 160462 996039 160468 996051
rect 157024 996011 160468 996039
rect 157024 995999 157030 996011
rect 160462 995999 160468 996011
rect 160520 995999 160526 996051
rect 174078 995999 174084 996051
rect 174136 996039 174142 996051
rect 212718 996039 212724 996051
rect 174136 996011 212724 996039
rect 174136 995999 174142 996011
rect 212718 995999 212724 996011
rect 212776 995999 212782 996051
rect 227714 995999 227720 996051
rect 227772 996039 227778 996051
rect 265066 996039 265072 996051
rect 227772 996011 265072 996039
rect 227772 995999 227778 996011
rect 265066 995999 265072 996011
rect 265124 996039 265130 996051
rect 267550 996039 267556 996051
rect 265124 996011 267556 996039
rect 265124 995999 265130 996011
rect 267550 995999 267556 996011
rect 267608 995999 267614 996051
rect 280338 995994 280344 996046
rect 280396 996034 280402 996046
rect 311802 996034 311808 996046
rect 280396 996006 311808 996034
rect 280396 995994 280402 996006
rect 311802 995994 311808 996006
rect 311860 995994 311866 996046
rect 92678 995976 92684 995988
rect 86604 995948 92684 995976
rect 86604 995852 86632 995948
rect 92678 995936 92684 995948
rect 92736 995936 92742 995988
rect 145190 995971 145196 995983
rect 136468 995943 145196 995971
rect 92402 995908 92408 995920
rect 91066 995880 92408 995908
rect 86586 995800 86592 995852
rect 86644 995800 86650 995852
rect 88978 995800 88984 995852
rect 89036 995840 89042 995852
rect 91066 995840 91094 995880
rect 92402 995868 92408 995880
rect 92460 995868 92466 995920
rect 92228 995840 92234 995852
rect 89036 995812 91094 995840
rect 91204 995812 92234 995840
rect 89036 995800 89042 995812
rect 86034 995732 86040 995784
rect 86092 995772 86098 995784
rect 91204 995772 91232 995812
rect 92228 995800 92234 995812
rect 92286 995800 92292 995852
rect 136266 995800 136272 995852
rect 136324 995840 136330 995852
rect 136468 995840 136496 995943
rect 145190 995931 145196 995943
rect 145248 995931 145254 995983
rect 195698 995971 195704 995983
rect 188724 995943 195704 995971
rect 143718 995908 143724 995914
rect 136836 995880 143724 995908
rect 136836 995852 136864 995880
rect 143718 995862 143724 995880
rect 143776 995862 143782 995914
rect 136324 995812 136496 995840
rect 136324 995800 136330 995812
rect 136818 995800 136824 995852
rect 136876 995800 136882 995852
rect 137922 995800 137928 995852
rect 137980 995840 137986 995852
rect 143626 995840 143632 995852
rect 137980 995812 143632 995840
rect 137980 995800 137986 995812
rect 143626 995800 143632 995812
rect 143684 995800 143690 995852
rect 86092 995744 91232 995772
rect 86092 995732 86098 995744
rect 91554 995732 91560 995784
rect 91612 995772 91618 995784
rect 92320 995772 92326 995784
rect 91612 995744 92326 995772
rect 91612 995732 91618 995744
rect 92320 995732 92326 995744
rect 92378 995732 92384 995784
rect 139210 995732 139216 995784
rect 139268 995772 139274 995784
rect 143810 995772 143816 995784
rect 139268 995744 143816 995772
rect 139268 995732 139274 995744
rect 143810 995732 143816 995744
rect 143868 995732 143874 995784
rect 183278 995732 183284 995784
rect 183336 995772 183342 995784
rect 188724 995772 188752 995943
rect 195698 995931 195704 995943
rect 195756 995931 195762 995983
rect 307754 995966 307760 995978
rect 286796 995938 307760 995966
rect 195606 995903 195612 995915
rect 188816 995875 195612 995903
rect 188816 995838 188844 995875
rect 195606 995863 195612 995875
rect 195664 995863 195670 995915
rect 246942 995908 246948 995920
rect 240888 995880 246948 995908
rect 240888 995852 240916 995880
rect 246942 995868 246948 995880
rect 247000 995868 247006 995920
rect 286796 995852 286824 995938
rect 307754 995926 307760 995938
rect 307812 995926 307818 995978
rect 383460 995936 383466 995988
rect 383518 995976 383524 995988
rect 383518 995948 391980 995976
rect 383518 995936 383524 995948
rect 306926 995898 306932 995910
rect 293604 995870 306932 995898
rect 188798 995786 188804 995838
rect 188856 995786 188862 995838
rect 189442 995790 189448 995842
rect 189500 995840 189506 995842
rect 195238 995840 195244 995847
rect 189500 995812 195244 995840
rect 189500 995790 189506 995812
rect 195238 995795 195244 995812
rect 195296 995795 195302 995847
rect 240870 995800 240876 995852
rect 240928 995800 240934 995852
rect 245562 995800 245568 995852
rect 245620 995840 245626 995852
rect 246482 995840 246488 995852
rect 245620 995812 246488 995840
rect 245620 995800 245626 995812
rect 246482 995800 246488 995812
rect 246540 995800 246546 995852
rect 286778 995800 286784 995852
rect 286836 995800 286842 995852
rect 293604 995842 293632 995870
rect 306926 995858 306932 995870
rect 306984 995858 306990 995910
rect 383368 995868 383374 995920
rect 383426 995908 383432 995920
rect 383426 995880 385724 995908
rect 383426 995868 383432 995880
rect 385696 995852 385724 995880
rect 391952 995852 391980 995948
rect 472158 995936 472164 995988
rect 472216 995976 472222 995988
rect 472216 995948 477494 995976
rect 472216 995936 472222 995948
rect 472710 995868 472716 995920
rect 472768 995908 472774 995920
rect 472768 995880 476436 995908
rect 472768 995868 472774 995880
rect 476408 995852 476436 995880
rect 293586 995790 293592 995842
rect 293644 995790 293650 995842
rect 295058 995790 295064 995842
rect 295116 995830 295122 995842
rect 310146 995830 310152 995852
rect 295116 995802 310152 995830
rect 295116 995790 295122 995802
rect 310146 995800 310152 995802
rect 310204 995800 310210 995852
rect 383736 995800 383742 995852
rect 383794 995840 383800 995852
rect 384390 995840 384396 995852
rect 383794 995812 384396 995840
rect 383794 995800 383800 995812
rect 384390 995800 384396 995812
rect 384448 995800 384454 995852
rect 385678 995800 385684 995852
rect 385736 995800 385742 995852
rect 391934 995800 391940 995852
rect 391992 995800 391998 995852
rect 396626 995800 396632 995852
rect 396684 995840 396690 995852
rect 400030 995840 400036 995852
rect 396684 995812 400036 995840
rect 396684 995800 396690 995812
rect 400030 995800 400036 995812
rect 400088 995800 400094 995852
rect 472526 995800 472532 995852
rect 472584 995840 472590 995852
rect 473998 995840 474004 995852
rect 472584 995812 474004 995840
rect 472584 995800 472590 995812
rect 473998 995800 474004 995812
rect 474056 995800 474062 995852
rect 476390 995800 476396 995852
rect 476448 995800 476454 995852
rect 477466 995840 477494 995948
rect 625614 995936 625620 995988
rect 625672 995976 625678 995988
rect 625672 995948 630628 995976
rect 625672 995936 625678 995948
rect 523586 995868 523592 995920
rect 523644 995908 523650 995920
rect 523644 995880 530164 995908
rect 523644 995868 523650 995880
rect 530136 995852 530164 995880
rect 625890 995868 625896 995920
rect 625948 995908 625954 995920
rect 625948 995880 627868 995908
rect 625948 995868 625954 995880
rect 627840 995852 627868 995880
rect 477678 995840 477684 995852
rect 477466 995812 477684 995840
rect 477678 995800 477684 995812
rect 477736 995800 477742 995852
rect 522942 995800 522948 995852
rect 523000 995840 523006 995852
rect 524782 995840 524788 995852
rect 523000 995812 524788 995840
rect 523000 995800 523006 995812
rect 524782 995800 524788 995812
rect 524840 995800 524846 995852
rect 530118 995800 530124 995852
rect 530176 995800 530182 995852
rect 537018 995800 537024 995852
rect 537076 995840 537082 995852
rect 540330 995840 540336 995852
rect 537076 995812 540336 995840
rect 537076 995800 537082 995812
rect 540330 995800 540336 995812
rect 540388 995800 540394 995852
rect 623682 995800 623688 995852
rect 623740 995840 623746 995852
rect 626534 995840 626540 995852
rect 623740 995812 626540 995840
rect 623740 995800 623746 995812
rect 626534 995800 626540 995812
rect 626592 995800 626598 995852
rect 627822 995800 627828 995852
rect 627880 995800 627886 995852
rect 630600 995840 630628 995948
rect 630858 995840 630864 995852
rect 630600 995812 630864 995840
rect 630858 995800 630864 995812
rect 630916 995800 630922 995852
rect 183336 995744 188752 995772
rect 183336 995732 183342 995744
rect 194318 995732 194324 995784
rect 194376 995772 194382 995784
rect 194376 995762 195082 995772
rect 195422 995762 195428 995784
rect 194376 995744 195428 995762
rect 194376 995732 194382 995744
rect 195046 995734 195428 995744
rect 195422 995732 195428 995734
rect 195480 995732 195486 995784
rect 239030 995732 239036 995784
rect 239088 995772 239094 995784
rect 246666 995772 246672 995784
rect 239088 995744 246672 995772
rect 239088 995732 239094 995744
rect 246666 995732 246672 995744
rect 246724 995732 246730 995784
rect 383644 995732 383650 995784
rect 383702 995772 383708 995784
rect 384942 995772 384948 995784
rect 383702 995744 384948 995772
rect 383702 995732 383708 995744
rect 384942 995732 384948 995744
rect 385000 995732 385006 995784
rect 472618 995732 472624 995784
rect 472676 995772 472682 995784
rect 473262 995772 473268 995784
rect 472676 995744 473268 995772
rect 472676 995732 472682 995744
rect 473262 995732 473268 995744
rect 473320 995732 473326 995784
rect 523770 995732 523776 995784
rect 523828 995772 523834 995784
rect 529014 995772 529020 995784
rect 523828 995744 529020 995772
rect 523828 995732 523834 995744
rect 529014 995732 529020 995744
rect 529072 995732 529078 995784
rect 625798 995732 625804 995784
rect 625856 995772 625862 995784
rect 627178 995772 627184 995784
rect 625856 995744 627184 995772
rect 625856 995732 625862 995744
rect 627178 995732 627184 995744
rect 627236 995732 627242 995784
rect 89714 995664 89720 995716
rect 89772 995704 89778 995716
rect 92586 995704 92592 995716
rect 89772 995676 92592 995704
rect 89772 995664 89778 995676
rect 92586 995664 92592 995676
rect 92644 995664 92650 995716
rect 141050 995664 141056 995716
rect 141108 995704 141114 995716
rect 154114 995704 154120 995716
rect 141108 995676 154120 995704
rect 141108 995664 141114 995676
rect 154114 995664 154120 995676
rect 154172 995664 154178 995716
rect 188154 995664 188160 995716
rect 188212 995704 188218 995716
rect 198642 995704 198648 995716
rect 188212 995676 198648 995704
rect 188212 995664 188218 995676
rect 198642 995664 198648 995676
rect 198700 995664 198706 995716
rect 243906 995664 243912 995716
rect 243964 995704 243970 995716
rect 246758 995704 246764 995716
rect 243964 995676 246764 995704
rect 243964 995664 243970 995676
rect 246758 995664 246764 995676
rect 246816 995664 246822 995716
rect 291746 995664 291752 995716
rect 291804 995704 291810 995716
rect 306466 995704 306472 995716
rect 291804 995676 306472 995704
rect 291804 995664 291810 995676
rect 306466 995664 306472 995676
rect 306524 995664 306530 995716
rect 383276 995664 383282 995716
rect 383334 995704 383340 995716
rect 388622 995704 388628 995716
rect 383334 995676 388628 995704
rect 383334 995664 383340 995676
rect 388622 995664 388628 995676
rect 388680 995664 388686 995716
rect 472434 995664 472440 995716
rect 472492 995704 472498 995716
rect 474734 995704 474740 995716
rect 472492 995676 474740 995704
rect 472492 995664 472498 995676
rect 474734 995664 474740 995676
rect 474792 995664 474798 995716
rect 521562 995664 521568 995716
rect 521620 995704 521626 995716
rect 532694 995704 532700 995716
rect 521620 995676 532700 995704
rect 521620 995664 521626 995676
rect 532694 995664 532700 995676
rect 532752 995664 532758 995716
rect 625706 995664 625712 995716
rect 625764 995704 625770 995716
rect 630214 995704 630220 995716
rect 625764 995676 630220 995704
rect 625764 995664 625770 995676
rect 630214 995664 630220 995676
rect 630272 995664 630278 995716
rect 77938 995596 77944 995648
rect 77996 995636 78002 995648
rect 92862 995636 92868 995648
rect 77996 995608 92868 995636
rect 77996 995596 78002 995608
rect 92862 995596 92868 995608
rect 92920 995596 92926 995648
rect 133138 995596 133144 995648
rect 133196 995636 133202 995648
rect 143902 995636 143908 995648
rect 133196 995608 143908 995636
rect 133196 995596 133202 995608
rect 143902 995596 143908 995608
rect 143960 995596 143966 995648
rect 184658 995596 184664 995648
rect 184716 995636 184722 995648
rect 198550 995636 198556 995648
rect 184716 995608 198556 995636
rect 184716 995596 184722 995608
rect 198550 995596 198556 995608
rect 198608 995596 198614 995648
rect 239582 995596 239588 995648
rect 239640 995636 239646 995648
rect 250622 995636 250628 995648
rect 239640 995608 250628 995636
rect 239640 995596 239646 995608
rect 250622 995596 250628 995608
rect 250680 995596 250686 995648
rect 287514 995596 287520 995648
rect 287572 995636 287578 995648
rect 307294 995636 307300 995648
rect 287572 995608 307300 995636
rect 287572 995596 287578 995608
rect 307294 995596 307300 995608
rect 307352 995596 307358 995648
rect 383552 995596 383558 995648
rect 383610 995636 383616 995648
rect 387518 995636 387524 995648
rect 383610 995608 387524 995636
rect 383610 995596 383616 995608
rect 387518 995596 387524 995608
rect 387576 995596 387582 995648
rect 472250 995596 472256 995648
rect 472308 995636 472314 995648
rect 481910 995636 481916 995648
rect 472308 995608 481916 995636
rect 472308 995596 472314 995608
rect 481910 995596 481916 995608
rect 481968 995596 481974 995648
rect 521470 995596 521476 995648
rect 521528 995636 521534 995648
rect 533430 995636 533436 995648
rect 521528 995608 533436 995636
rect 521528 995596 521534 995608
rect 533430 995596 533436 995608
rect 533488 995596 533494 995648
rect 625430 995596 625436 995648
rect 625488 995636 625494 995648
rect 631502 995636 631508 995648
rect 625488 995608 631508 995636
rect 625488 995596 625494 995608
rect 631502 995596 631508 995608
rect 631560 995596 631566 995648
rect 132402 995528 132408 995580
rect 132460 995568 132466 995580
rect 144914 995568 144920 995580
rect 132460 995540 144920 995568
rect 132460 995528 132466 995540
rect 144914 995528 144920 995540
rect 144972 995528 144978 995580
rect 190638 995528 190644 995580
rect 190696 995568 190702 995580
rect 195514 995568 195520 995580
rect 190696 995540 195520 995568
rect 190696 995528 190702 995540
rect 195514 995528 195520 995540
rect 195572 995528 195578 995580
rect 383184 995528 383190 995580
rect 383242 995568 383248 995580
rect 389358 995568 389364 995580
rect 383242 995540 389364 995568
rect 383242 995528 383248 995540
rect 389358 995528 389364 995540
rect 389416 995528 389422 995580
rect 472342 995528 472348 995580
rect 472400 995568 472406 995580
rect 476942 995568 476948 995580
rect 472400 995540 476948 995568
rect 472400 995528 472406 995540
rect 476942 995528 476948 995540
rect 477000 995528 477006 995580
rect 482646 995568 482652 995580
rect 477144 995540 482652 995568
rect 130010 995460 130016 995512
rect 130068 995500 130074 995512
rect 144086 995500 144092 995512
rect 130068 995472 144092 995500
rect 130068 995460 130074 995472
rect 144086 995460 144092 995472
rect 144144 995460 144150 995512
rect 184474 995460 184480 995512
rect 184532 995500 184538 995512
rect 198458 995500 198464 995512
rect 184532 995472 198464 995500
rect 184532 995460 184538 995472
rect 198458 995460 198464 995472
rect 198516 995460 198522 995512
rect 380986 995460 380992 995512
rect 381044 995500 381050 995512
rect 393590 995500 393596 995512
rect 381044 995472 393596 995500
rect 381044 995460 381050 995472
rect 393590 995460 393596 995472
rect 393648 995460 393654 995512
rect 131850 995392 131856 995444
rect 131908 995432 131914 995444
rect 145098 995432 145104 995444
rect 131908 995404 145104 995432
rect 131908 995392 131914 995404
rect 145098 995392 145104 995404
rect 145156 995392 145162 995444
rect 183830 995392 183836 995444
rect 183888 995432 183894 995444
rect 198366 995432 198372 995444
rect 183888 995404 198372 995432
rect 183888 995392 183894 995404
rect 198366 995392 198372 995404
rect 198424 995392 198430 995444
rect 469398 995392 469404 995444
rect 469456 995432 469462 995444
rect 477144 995432 477172 995540
rect 482646 995528 482652 995540
rect 482704 995528 482710 995580
rect 521286 995528 521292 995580
rect 521344 995568 521350 995580
rect 533982 995568 533988 995580
rect 521344 995540 533988 995568
rect 521344 995528 521350 995540
rect 533982 995528 533988 995540
rect 534040 995528 534046 995580
rect 623774 995528 623780 995580
rect 623832 995568 623838 995580
rect 635826 995568 635832 995580
rect 623832 995540 635832 995568
rect 623832 995528 623838 995540
rect 635826 995528 635832 995540
rect 635884 995528 635890 995580
rect 469456 995404 477172 995432
rect 469456 995392 469462 995404
rect 469214 995324 469220 995376
rect 469272 995364 469278 995376
rect 480806 995364 480812 995376
rect 469272 995336 480812 995364
rect 469272 995324 469278 995336
rect 480806 995324 480812 995336
rect 480864 995324 480870 995376
rect 303522 994720 303528 994772
rect 303580 994720 303586 994772
rect 283466 993828 283472 993880
rect 283524 993868 283530 993880
rect 301774 993868 301780 993880
rect 283524 993840 301780 993868
rect 283524 993828 283530 993840
rect 301774 993828 301780 993840
rect 301832 993828 301838 993880
rect 378318 993828 378324 993880
rect 378376 993868 378382 993880
rect 392670 993868 392676 993880
rect 378376 993840 392676 993868
rect 378376 993828 378382 993840
rect 392670 993828 392676 993840
rect 392728 993828 392734 993880
rect 145006 993800 145012 993812
rect 129706 993772 145012 993800
rect 129090 993692 129096 993744
rect 129148 993732 129154 993744
rect 129706 993732 129734 993772
rect 145006 993760 145012 993772
rect 145064 993760 145070 993812
rect 180150 993760 180156 993812
rect 180208 993800 180214 993812
rect 200022 993800 200028 993812
rect 180208 993772 200028 993800
rect 180208 993760 180214 993772
rect 200022 993760 200028 993772
rect 200080 993760 200086 993812
rect 285950 993760 285956 993812
rect 286008 993800 286014 993812
rect 309318 993800 309324 993812
rect 286008 993772 309324 993800
rect 286008 993760 286014 993772
rect 309318 993760 309324 993772
rect 309376 993760 309382 993812
rect 469306 993760 469312 993812
rect 469364 993800 469370 993812
rect 487798 993800 487804 993812
rect 469364 993772 487804 993800
rect 469364 993760 469370 993772
rect 487798 993760 487804 993772
rect 487856 993760 487862 993812
rect 521378 993760 521384 993812
rect 521436 993800 521442 993812
rect 535546 993800 535552 993812
rect 521436 993772 535552 993800
rect 521436 993760 521442 993772
rect 535546 993760 535552 993772
rect 535604 993760 535610 993812
rect 129148 993704 129734 993732
rect 129148 993692 129154 993704
rect 140498 993692 140504 993744
rect 140556 993732 140562 993744
rect 151814 993732 151820 993744
rect 140556 993704 151820 993732
rect 140556 993692 140562 993704
rect 151814 993692 151820 993704
rect 151872 993692 151878 993744
rect 180794 993692 180800 993744
rect 180852 993732 180858 993744
rect 200114 993732 200120 993744
rect 180852 993704 200120 993732
rect 180852 993692 180858 993704
rect 200114 993692 200120 993704
rect 200172 993692 200178 993744
rect 282822 993692 282828 993744
rect 282880 993732 282886 993744
rect 314930 993732 314936 993744
rect 282880 993704 314936 993732
rect 282880 993692 282886 993704
rect 314930 993692 314936 993704
rect 314988 993692 314994 993744
rect 374454 993692 374460 993744
rect 374512 993732 374518 993744
rect 393314 993732 393320 993744
rect 374512 993704 393320 993732
rect 374512 993692 374518 993704
rect 393314 993692 393320 993704
rect 393372 993692 393378 993744
rect 470870 993692 470876 993744
rect 470928 993732 470934 993744
rect 484118 993732 484124 993744
rect 470928 993704 484124 993732
rect 470928 993692 470934 993704
rect 484118 993692 484124 993704
rect 484176 993692 484182 993744
rect 571610 993692 571616 993744
rect 571668 993732 571674 993744
rect 633986 993732 633992 993744
rect 571668 993704 633992 993732
rect 571668 993692 571674 993704
rect 633986 993692 633992 993704
rect 634044 993692 634050 993744
rect 77018 993624 77024 993676
rect 77076 993664 77082 993676
rect 104158 993664 104164 993676
rect 77076 993636 104164 993664
rect 77076 993624 77082 993636
rect 104158 993624 104164 993636
rect 104216 993624 104222 993676
rect 128446 993624 128452 993676
rect 128504 993664 128510 993676
rect 160278 993664 160284 993676
rect 128504 993636 160284 993664
rect 128504 993624 128510 993636
rect 160278 993624 160284 993636
rect 160336 993624 160342 993676
rect 181438 993624 181444 993676
rect 181496 993664 181502 993676
rect 207566 993664 207572 993676
rect 181496 993636 207572 993664
rect 181496 993624 181502 993636
rect 207566 993624 207572 993636
rect 207624 993624 207630 993676
rect 231578 993624 231584 993676
rect 231636 993664 231642 993676
rect 262214 993664 262220 993676
rect 231636 993636 262220 993664
rect 231636 993624 231642 993636
rect 262214 993624 262220 993636
rect 262272 993624 262278 993676
rect 284110 993624 284116 993676
rect 284168 993664 284174 993676
rect 310606 993664 310612 993676
rect 284168 993636 310612 993664
rect 284168 993624 284174 993636
rect 310606 993624 310612 993636
rect 310664 993624 310670 993676
rect 355962 993624 355968 993676
rect 356020 993664 356026 993676
rect 398834 993664 398840 993676
rect 356020 993636 398840 993664
rect 356020 993624 356026 993636
rect 398834 993624 398840 993636
rect 398892 993624 398898 993676
rect 462774 993624 462780 993676
rect 462832 993664 462838 993676
rect 485958 993664 485964 993676
rect 462832 993636 485964 993664
rect 462832 993624 462838 993636
rect 485958 993624 485964 993636
rect 486016 993624 486022 993676
rect 499482 993624 499488 993676
rect 499540 993664 499546 993676
rect 539226 993664 539232 993676
rect 499540 993636 539232 993664
rect 499540 993624 499546 993636
rect 539226 993624 539232 993636
rect 539284 993624 539290 993676
rect 551646 993624 551652 993676
rect 551704 993664 551710 993676
rect 640702 993664 640708 993676
rect 551704 993636 640708 993664
rect 551704 993624 551710 993636
rect 640702 993624 640708 993636
rect 640760 993624 640766 993676
rect 433518 993556 433524 993608
rect 433576 993596 433582 993608
rect 434622 993596 434628 993608
rect 433576 993568 434628 993596
rect 433576 993556 433582 993568
rect 434622 993556 434628 993568
rect 434680 993596 434686 993608
rect 510706 993596 510712 993608
rect 434680 993568 510712 993596
rect 434680 993556 434686 993568
rect 510706 993556 510712 993568
rect 510764 993556 510770 993608
rect 510890 993556 510896 993608
rect 510948 993596 510954 993608
rect 511902 993596 511908 993608
rect 510948 993568 511908 993596
rect 510948 993556 510954 993568
rect 511902 993556 511908 993568
rect 511960 993596 511966 993608
rect 563146 993596 563152 993608
rect 511960 993568 563152 993596
rect 511960 993556 511966 993568
rect 563146 993556 563152 993568
rect 563204 993556 563210 993608
rect 368566 993488 368572 993540
rect 368624 993528 368630 993540
rect 433426 993528 433432 993540
rect 368624 993500 433432 993528
rect 368624 993488 368630 993500
rect 433426 993488 433432 993500
rect 433484 993488 433490 993540
rect 433610 993488 433616 993540
rect 433668 993528 433674 993540
rect 434806 993528 434812 993540
rect 433668 993500 434812 993528
rect 433668 993488 433674 993500
rect 434806 993488 434812 993500
rect 434864 993528 434870 993540
rect 510614 993528 510620 993540
rect 434864 993500 510620 993528
rect 434864 993488 434870 993500
rect 510614 993488 510620 993500
rect 510672 993488 510678 993540
rect 510798 993488 510804 993540
rect 510856 993528 510862 993540
rect 512086 993528 512092 993540
rect 510856 993500 512092 993528
rect 510856 993488 510862 993500
rect 512086 993488 512092 993500
rect 512144 993528 512150 993540
rect 563054 993528 563060 993540
rect 512144 993500 563060 993528
rect 512144 993488 512150 993500
rect 563054 993488 563060 993500
rect 563112 993488 563118 993540
rect 368750 993420 368756 993472
rect 368808 993460 368814 993472
rect 433334 993460 433340 993472
rect 368808 993432 433340 993460
rect 368808 993420 368814 993432
rect 433334 993420 433340 993432
rect 433392 993420 433398 993472
rect 436186 993420 436192 993472
rect 436244 993460 436250 993472
rect 437934 993460 437940 993472
rect 436244 993432 437940 993460
rect 436244 993420 436250 993432
rect 437934 993420 437940 993432
rect 437992 993460 437998 993472
rect 513374 993460 513380 993472
rect 437992 993432 513380 993460
rect 437992 993420 437998 993432
rect 513374 993420 513380 993432
rect 513432 993420 513438 993472
rect 513466 993420 513472 993472
rect 513524 993460 513530 993472
rect 515214 993460 515220 993472
rect 513524 993432 515220 993460
rect 513524 993420 513530 993432
rect 515214 993420 515220 993432
rect 515272 993460 515278 993472
rect 565814 993460 565820 993472
rect 515272 993432 565820 993460
rect 515272 993420 515278 993432
rect 565814 993420 565820 993432
rect 565872 993420 565878 993472
rect 368382 993352 368388 993404
rect 368440 993392 368446 993404
rect 436094 993392 436100 993404
rect 368440 993364 436100 993392
rect 368440 993352 368446 993364
rect 436094 993352 436100 993364
rect 436152 993352 436158 993404
rect 89622 990768 89628 990820
rect 89680 990808 89686 990820
rect 92494 990808 92500 990820
rect 89680 990780 92500 990808
rect 89680 990768 89686 990780
rect 92494 990768 92500 990780
rect 92552 990768 92558 990820
rect 564250 990768 564256 990820
rect 564308 990808 564314 990820
rect 576302 990808 576308 990820
rect 564308 990780 576308 990808
rect 564308 990768 564314 990780
rect 576302 990768 576308 990780
rect 576360 990768 576366 990820
rect 168374 990632 168380 990684
rect 168432 990672 168438 990684
rect 170398 990672 170404 990684
rect 168432 990644 170404 990672
rect 168432 990632 168438 990644
rect 170398 990632 170404 990644
rect 170456 990632 170462 990684
rect 203150 990632 203156 990684
rect 203208 990672 203214 990684
rect 204162 990672 204168 990684
rect 203208 990644 204168 990672
rect 203208 990632 203214 990644
rect 204162 990632 204168 990644
rect 204220 990632 204226 990684
rect 331214 990632 331220 990684
rect 331272 990672 331278 990684
rect 332686 990672 332692 990684
rect 331272 990644 332692 990672
rect 331272 990632 331278 990644
rect 332686 990632 332692 990644
rect 332744 990632 332750 990684
rect 444374 990632 444380 990684
rect 444432 990672 444438 990684
rect 446214 990672 446220 990684
rect 444432 990644 446220 990672
rect 444432 990632 444438 990644
rect 446214 990632 446220 990644
rect 446272 990632 446278 990684
rect 366174 989680 366180 989732
rect 366232 989720 366238 989732
rect 381630 989720 381636 989732
rect 366232 989692 381636 989720
rect 366232 989680 366238 989692
rect 381630 989680 381636 989692
rect 381688 989680 381694 989732
rect 371142 989612 371148 989664
rect 371200 989652 371206 989664
rect 397822 989652 397828 989664
rect 371200 989624 397828 989652
rect 371200 989612 371206 989624
rect 397822 989612 397828 989624
rect 397880 989612 397886 989664
rect 437750 989612 437756 989664
rect 437808 989652 437814 989664
rect 462774 989652 462780 989664
rect 437808 989624 462780 989652
rect 437808 989612 437814 989624
rect 462774 989612 462780 989624
rect 462832 989612 462838 989664
rect 514846 989612 514852 989664
rect 514904 989652 514910 989664
rect 527634 989652 527640 989664
rect 514904 989624 527640 989652
rect 514904 989612 514910 989624
rect 527634 989612 527640 989624
rect 527692 989612 527698 989664
rect 567102 989612 567108 989664
rect 567160 989652 567166 989664
rect 592494 989652 592500 989664
rect 567160 989624 592500 989652
rect 567160 989612 567166 989624
rect 592494 989612 592500 989624
rect 592552 989612 592558 989664
rect 321462 989544 321468 989596
rect 321520 989584 321526 989596
rect 349154 989584 349160 989596
rect 321520 989556 349160 989584
rect 321520 989544 321526 989556
rect 349154 989544 349160 989556
rect 349212 989544 349218 989596
rect 371326 989544 371332 989596
rect 371384 989584 371390 989596
rect 414106 989584 414112 989596
rect 371384 989556 414112 989584
rect 371384 989544 371390 989556
rect 414106 989544 414112 989556
rect 414164 989544 414170 989596
rect 437382 989544 437388 989596
rect 437440 989584 437446 989596
rect 478966 989584 478972 989596
rect 437440 989556 478972 989584
rect 437440 989544 437446 989556
rect 478966 989544 478972 989556
rect 479024 989544 479030 989596
rect 515030 989544 515036 989596
rect 515088 989584 515094 989596
rect 543826 989584 543832 989596
rect 515088 989556 543832 989584
rect 515088 989544 515094 989556
rect 543826 989544 543832 989556
rect 543884 989544 543890 989596
rect 567470 989544 567476 989596
rect 567528 989584 567534 989596
rect 608778 989584 608784 989596
rect 567528 989556 608784 989584
rect 567528 989544 567534 989556
rect 608778 989544 608784 989556
rect 608836 989544 608842 989596
rect 269206 989476 269212 989528
rect 269264 989516 269270 989528
rect 300486 989516 300492 989528
rect 269264 989488 300492 989516
rect 269264 989476 269270 989488
rect 300486 989476 300492 989488
rect 300544 989476 300550 989528
rect 319070 989476 319076 989528
rect 319128 989516 319134 989528
rect 365438 989516 365444 989528
rect 319128 989488 365444 989516
rect 319128 989476 319134 989488
rect 365438 989476 365444 989488
rect 365496 989476 365502 989528
rect 371510 989476 371516 989528
rect 371568 989516 371574 989528
rect 430298 989516 430304 989528
rect 371568 989488 430304 989516
rect 371568 989476 371574 989488
rect 430298 989476 430304 989488
rect 430356 989476 430362 989528
rect 437566 989476 437572 989528
rect 437624 989516 437630 989528
rect 495158 989516 495164 989528
rect 437624 989488 495164 989516
rect 437624 989476 437630 989488
rect 495158 989476 495164 989488
rect 495216 989476 495222 989528
rect 514662 989476 514668 989528
rect 514720 989516 514726 989528
rect 560110 989516 560116 989528
rect 514720 989488 560116 989516
rect 514720 989476 514726 989488
rect 560110 989476 560116 989488
rect 560168 989476 560174 989528
rect 567286 989476 567292 989528
rect 567344 989516 567350 989528
rect 624970 989516 624976 989528
rect 567344 989488 624976 989516
rect 567344 989476 567350 989488
rect 624970 989476 624976 989488
rect 625028 989476 625034 989528
rect 73430 989408 73436 989460
rect 73488 989448 73494 989460
rect 92954 989448 92960 989460
rect 73488 989420 92960 989448
rect 73488 989408 73494 989420
rect 92954 989408 92960 989420
rect 93012 989408 93018 989460
rect 105814 989408 105820 989460
rect 105872 989448 105878 989460
rect 113266 989448 113272 989460
rect 105872 989420 113272 989448
rect 105872 989408 105878 989420
rect 113266 989408 113272 989420
rect 113324 989408 113330 989460
rect 151814 989408 151820 989460
rect 151872 989448 151878 989460
rect 186958 989448 186964 989460
rect 151872 989420 186964 989448
rect 151872 989408 151878 989420
rect 186958 989408 186964 989420
rect 187016 989408 187022 989460
rect 216582 989408 216588 989460
rect 216640 989448 216646 989460
rect 235626 989448 235632 989460
rect 216640 989420 235632 989448
rect 216640 989408 216646 989420
rect 235626 989408 235632 989420
rect 235684 989408 235690 989460
rect 269022 989408 269028 989460
rect 269080 989448 269086 989460
rect 284294 989448 284300 989460
rect 269080 989420 284300 989448
rect 269080 989408 269086 989420
rect 284294 989408 284300 989420
rect 284352 989408 284358 989460
rect 303522 989408 303528 989460
rect 303580 989448 303586 989460
rect 666554 989448 666560 989460
rect 303580 989420 666560 989448
rect 303580 989408 303586 989420
rect 666554 989408 666560 989420
rect 666612 989408 666618 989460
rect 138290 988728 138296 988780
rect 138348 988768 138354 988780
rect 144822 988768 144828 988780
rect 138348 988740 144828 988768
rect 138348 988728 138354 988740
rect 144822 988728 144828 988740
rect 144880 988728 144886 988780
rect 248322 988116 248328 988168
rect 248380 988156 248386 988168
rect 251818 988156 251824 988168
rect 248380 988128 251824 988156
rect 248380 988116 248386 988128
rect 251818 988116 251824 988128
rect 251876 988116 251882 988168
rect 45462 988048 45468 988100
rect 45520 988088 45526 988100
rect 367186 988088 367192 988100
rect 45520 988060 367192 988088
rect 45520 988048 45526 988060
rect 367186 988048 367192 988060
rect 367244 988048 367250 988100
rect 45738 987980 45744 988032
rect 45796 988020 45802 988032
rect 368750 988020 368756 988032
rect 45796 987992 368756 988020
rect 45796 987980 45802 987992
rect 368750 987980 368756 987992
rect 368808 987980 368814 988032
rect 45554 987912 45560 987964
rect 45612 987952 45618 987964
rect 369854 987952 369860 987964
rect 45612 987924 369860 987952
rect 45612 987912 45618 987924
rect 369854 987912 369860 987924
rect 369912 987912 369918 987964
rect 314286 987844 314292 987896
rect 314344 987884 314350 987896
rect 666830 987884 666836 987896
rect 314344 987856 666836 987884
rect 314344 987844 314350 987856
rect 666830 987844 666836 987856
rect 666888 987844 666894 987896
rect 318886 987776 318892 987828
rect 318944 987816 318950 987828
rect 669222 987816 669228 987828
rect 318944 987788 669228 987816
rect 318944 987776 318950 987788
rect 669222 987776 669228 987788
rect 669280 987776 669286 987828
rect 311802 987708 311808 987760
rect 311860 987748 311866 987760
rect 666646 987748 666652 987760
rect 311860 987720 666652 987748
rect 311860 987708 311866 987720
rect 666646 987708 666652 987720
rect 666704 987708 666710 987760
rect 318702 987640 318708 987692
rect 318760 987680 318766 987692
rect 669314 987680 669320 987692
rect 318760 987652 669320 987680
rect 318760 987640 318766 987652
rect 669314 987640 669320 987652
rect 669372 987640 669378 987692
rect 280062 987572 280068 987624
rect 280120 987612 280126 987624
rect 651374 987612 651380 987624
rect 280120 987584 651380 987612
rect 280120 987572 280126 987584
rect 651374 987572 651380 987584
rect 651432 987572 651438 987624
rect 270402 987504 270408 987556
rect 270460 987544 270466 987556
rect 652846 987544 652852 987556
rect 270460 987516 652852 987544
rect 270460 987504 270466 987516
rect 652846 987504 652852 987516
rect 652904 987504 652910 987556
rect 267642 987436 267648 987488
rect 267700 987476 267706 987488
rect 652662 987476 652668 987488
rect 267700 987448 652668 987476
rect 267700 987436 267706 987448
rect 652662 987436 652668 987448
rect 652720 987436 652726 987488
rect 48222 987368 48228 987420
rect 48280 987408 48286 987420
rect 433518 987408 433524 987420
rect 48280 987380 433524 987408
rect 48280 987368 48286 987380
rect 433518 987368 433524 987380
rect 433576 987368 433582 987420
rect 267550 987300 267556 987352
rect 267608 987340 267614 987352
rect 652754 987340 652760 987352
rect 267608 987312 652760 987340
rect 267608 987300 267614 987312
rect 652754 987300 652760 987312
rect 652812 987300 652818 987352
rect 227622 987232 227628 987284
rect 227680 987272 227686 987284
rect 651466 987272 651472 987284
rect 227680 987244 651472 987272
rect 227680 987232 227686 987244
rect 651466 987232 651472 987244
rect 651524 987232 651530 987284
rect 212626 987164 212632 987216
rect 212684 987204 212690 987216
rect 652938 987204 652944 987216
rect 212684 987176 652944 987204
rect 212684 987164 212690 987176
rect 652938 987164 652944 987176
rect 652996 987164 653002 987216
rect 215294 987096 215300 987148
rect 215352 987136 215358 987148
rect 658274 987136 658280 987148
rect 215352 987108 658280 987136
rect 215352 987096 215358 987108
rect 658274 987096 658280 987108
rect 658332 987096 658338 987148
rect 212718 987028 212724 987080
rect 212776 987068 212782 987080
rect 658182 987068 658188 987080
rect 212776 987040 658188 987068
rect 212776 987028 212782 987040
rect 658182 987028 658188 987040
rect 658240 987028 658246 987080
rect 175182 986960 175188 987012
rect 175240 987000 175246 987012
rect 651558 987000 651564 987012
rect 175240 986972 651564 987000
rect 175240 986960 175246 986972
rect 651558 986960 651564 986972
rect 651616 986960 651622 987012
rect 125502 986892 125508 986944
rect 125560 986932 125566 986944
rect 651650 986932 651656 986944
rect 125560 986904 651656 986932
rect 125560 986892 125566 986904
rect 651650 986892 651656 986904
rect 651708 986892 651714 986944
rect 62666 986824 62672 986876
rect 62724 986864 62730 986876
rect 113358 986864 113364 986876
rect 62724 986836 113364 986864
rect 62724 986824 62730 986836
rect 113358 986824 113364 986836
rect 113416 986864 113422 986876
rect 669590 986864 669596 986876
rect 113416 986836 669596 986864
rect 113416 986824 113422 986836
rect 669590 986824 669596 986836
rect 669648 986824 669654 986876
rect 62482 986756 62488 986808
rect 62540 986796 62546 986808
rect 110506 986796 110512 986808
rect 62540 986768 110512 986796
rect 62540 986756 62546 986768
rect 110506 986756 110512 986768
rect 110564 986796 110570 986808
rect 669406 986796 669412 986808
rect 110564 986768 669412 986796
rect 110564 986756 110570 986768
rect 669406 986756 669412 986768
rect 669464 986756 669470 986808
rect 62298 986688 62304 986740
rect 62356 986728 62362 986740
rect 110598 986728 110604 986740
rect 62356 986700 110604 986728
rect 62356 986688 62362 986700
rect 110598 986688 110604 986700
rect 110656 986728 110662 986740
rect 669498 986728 669504 986740
rect 110656 986700 669504 986728
rect 110656 986688 110662 986700
rect 669498 986688 669504 986700
rect 669556 986688 669562 986740
rect 564526 985464 564532 985516
rect 564584 985504 564590 985516
rect 564710 985504 564716 985516
rect 564584 985476 564716 985504
rect 564584 985464 564590 985476
rect 564710 985464 564716 985476
rect 564768 985504 564774 985516
rect 675662 985504 675668 985516
rect 564768 985476 675668 985504
rect 564768 985464 564774 985476
rect 675662 985464 675668 985476
rect 675720 985464 675726 985516
rect 62850 985396 62856 985448
rect 62908 985436 62914 985448
rect 669682 985436 669688 985448
rect 62908 985408 669688 985436
rect 62908 985396 62914 985408
rect 669682 985396 669688 985408
rect 669740 985396 669746 985448
rect 62390 985328 62396 985380
rect 62448 985368 62454 985380
rect 670050 985368 670056 985380
rect 62448 985340 670056 985368
rect 62448 985328 62454 985340
rect 670050 985328 670056 985340
rect 670108 985328 670114 985380
rect 350442 985056 350448 985108
rect 350500 985096 350506 985108
rect 670970 985096 670976 985108
rect 350500 985068 670976 985096
rect 350500 985056 350506 985068
rect 670970 985056 670976 985068
rect 671028 985056 671034 985108
rect 45646 984988 45652 985040
rect 45704 985028 45710 985040
rect 367094 985028 367100 985040
rect 45704 985000 367100 985028
rect 45704 984988 45710 985000
rect 367094 984988 367100 985000
rect 367152 984988 367158 985040
rect 45922 984920 45928 984972
rect 45980 984960 45986 984972
rect 368566 984960 368572 984972
rect 45980 984932 368572 984960
rect 45980 984920 45986 984932
rect 368566 984920 368572 984932
rect 368624 984920 368630 984972
rect 45830 984852 45836 984904
rect 45888 984892 45894 984904
rect 368382 984892 368388 984904
rect 45888 984864 368388 984892
rect 45888 984852 45894 984864
rect 368382 984852 368388 984864
rect 368440 984852 368446 984904
rect 419074 984852 419080 984904
rect 419132 984892 419138 984904
rect 670878 984892 670884 984904
rect 419132 984864 670884 984892
rect 419132 984852 419138 984864
rect 670878 984852 670884 984864
rect 670936 984852 670942 984904
rect 317506 984784 317512 984836
rect 317564 984824 317570 984836
rect 666738 984824 666744 984836
rect 317564 984796 666744 984824
rect 317564 984784 317570 984796
rect 666738 984784 666744 984796
rect 666796 984784 666802 984836
rect 315942 984716 315948 984768
rect 316000 984756 316006 984768
rect 671982 984756 671988 984768
rect 316000 984728 671988 984756
rect 316000 984716 316006 984728
rect 671982 984716 671988 984728
rect 672040 984716 672046 984768
rect 300762 984648 300768 984700
rect 300820 984688 300826 984700
rect 671062 984688 671068 984700
rect 300820 984660 671068 984688
rect 300820 984648 300826 984660
rect 671062 984648 671068 984660
rect 671120 984648 671126 984700
rect 46106 984580 46112 984632
rect 46164 984620 46170 984632
rect 433610 984620 433616 984632
rect 46164 984592 433616 984620
rect 46164 984580 46170 984592
rect 433610 984580 433616 984592
rect 433668 984580 433674 984632
rect 48314 984512 48320 984564
rect 48372 984552 48378 984564
rect 436186 984552 436192 984564
rect 48372 984524 436192 984552
rect 48372 984512 48378 984524
rect 436186 984512 436192 984524
rect 436244 984512 436250 984564
rect 496630 984512 496636 984564
rect 496688 984552 496694 984564
rect 670786 984552 670792 984564
rect 496688 984524 670792 984552
rect 496688 984512 496694 984524
rect 670786 984512 670792 984524
rect 670844 984512 670850 984564
rect 46382 984444 46388 984496
rect 46440 984484 46446 984496
rect 510798 984484 510804 984496
rect 46440 984456 510804 984484
rect 46440 984444 46446 984456
rect 510798 984444 510804 984456
rect 510856 984444 510862 984496
rect 46198 984376 46204 984428
rect 46256 984416 46262 984428
rect 510890 984416 510896 984428
rect 46256 984388 510896 984416
rect 46256 984376 46262 984388
rect 510890 984376 510896 984388
rect 510948 984376 510954 984428
rect 48406 984308 48412 984360
rect 48464 984348 48470 984360
rect 513466 984348 513472 984360
rect 48464 984320 513472 984348
rect 48464 984308 48470 984320
rect 513466 984308 513472 984320
rect 513524 984308 513530 984360
rect 546402 984308 546408 984360
rect 546460 984348 546466 984360
rect 670694 984348 670700 984360
rect 546460 984320 670700 984348
rect 546460 984308 546466 984320
rect 670694 984308 670700 984320
rect 670752 984308 670758 984360
rect 162854 984240 162860 984292
rect 162912 984280 162918 984292
rect 655422 984280 655428 984292
rect 162912 984252 655428 984280
rect 162912 984240 162918 984252
rect 655422 984240 655428 984252
rect 655480 984240 655486 984292
rect 162946 984172 162952 984224
rect 163004 984212 163010 984224
rect 658458 984212 658464 984224
rect 163004 984184 658464 984212
rect 163004 984172 163010 984184
rect 658458 984172 658464 984184
rect 658516 984172 658522 984224
rect 46014 984104 46020 984156
rect 46072 984144 46078 984156
rect 110414 984144 110420 984156
rect 46072 984116 110420 984144
rect 46072 984104 46078 984116
rect 110414 984104 110420 984116
rect 110472 984104 110478 984156
rect 160462 984104 160468 984156
rect 160520 984144 160526 984156
rect 658366 984144 658372 984156
rect 160520 984116 658372 984144
rect 160520 984104 160526 984116
rect 658366 984104 658372 984116
rect 658424 984104 658430 984156
rect 62206 984036 62212 984088
rect 62264 984076 62270 984088
rect 561030 984076 561036 984088
rect 62264 984048 561036 984076
rect 62264 984036 62270 984048
rect 561030 984036 561036 984048
rect 561088 984036 561094 984088
rect 564342 984036 564348 984088
rect 564400 984076 564406 984088
rect 649902 984076 649908 984088
rect 564400 984048 649908 984076
rect 564400 984036 564406 984048
rect 649902 984036 649908 984048
rect 649960 984036 649966 984088
rect 62114 983968 62120 984020
rect 62172 984008 62178 984020
rect 564526 984008 564532 984020
rect 62172 983980 564532 984008
rect 62172 983968 62178 983980
rect 564526 983968 564532 983980
rect 564584 983968 564590 984020
rect 62022 983900 62028 983952
rect 62080 983940 62086 983952
rect 564434 983940 564440 983952
rect 62080 983912 564440 983940
rect 62080 983900 62086 983912
rect 564434 983900 564440 983912
rect 564492 983900 564498 983952
rect 62574 983084 62580 983136
rect 62632 983124 62638 983136
rect 668946 983124 668952 983136
rect 62632 983096 668952 983124
rect 62632 983084 62638 983096
rect 668946 983084 668952 983096
rect 669004 983084 669010 983136
rect 62758 983016 62764 983068
rect 62816 983056 62822 983068
rect 670234 983056 670240 983068
rect 62816 983028 670240 983056
rect 62816 983016 62822 983028
rect 670234 983016 670240 983028
rect 670292 983016 670298 983068
rect 63126 982948 63132 983000
rect 63184 982988 63190 983000
rect 668578 982988 668584 983000
rect 63184 982960 668584 982988
rect 63184 982948 63190 982960
rect 668578 982948 668584 982960
rect 668636 982948 668642 983000
rect 62942 982880 62948 982932
rect 63000 982920 63006 982932
rect 668486 982920 668492 982932
rect 63000 982892 668492 982920
rect 63000 982880 63006 982892
rect 668486 982880 668492 982892
rect 668544 982880 668550 982932
rect 42334 972884 42340 972936
rect 42392 972924 42398 972936
rect 58434 972924 58440 972936
rect 42392 972896 58440 972924
rect 42392 972884 42398 972896
rect 58434 972884 58440 972896
rect 58492 972884 58498 972936
rect 674834 970096 674840 970148
rect 674892 970136 674898 970148
rect 675662 970136 675668 970148
rect 674892 970108 675668 970136
rect 674892 970096 674898 970108
rect 675662 970096 675668 970108
rect 675720 970096 675726 970148
rect 42150 967240 42156 967292
rect 42208 967280 42214 967292
rect 42334 967280 42340 967292
rect 42208 967252 42340 967280
rect 42208 967240 42214 967252
rect 42334 967240 42340 967252
rect 42392 967240 42398 967292
rect 42058 967036 42064 967088
rect 42116 967076 42122 967088
rect 42794 967076 42800 967088
rect 42116 967048 42800 967076
rect 42116 967036 42122 967048
rect 42794 967036 42800 967048
rect 42852 967036 42858 967088
rect 673546 966356 673552 966408
rect 673604 966396 673610 966408
rect 675386 966396 675392 966408
rect 673604 966368 675392 966396
rect 673604 966356 673610 966368
rect 675386 966356 675392 966368
rect 675444 966356 675450 966408
rect 674742 965540 674748 965592
rect 674800 965580 674806 965592
rect 675386 965580 675392 965592
rect 674800 965552 675392 965580
rect 674800 965540 674806 965552
rect 675386 965540 675392 965552
rect 675444 965540 675450 965592
rect 673454 964996 673460 965048
rect 673512 965036 673518 965048
rect 675478 965036 675484 965048
rect 673512 965008 675484 965036
rect 673512 964996 673518 965008
rect 675478 964996 675484 965008
rect 675536 964996 675542 965048
rect 42150 963976 42156 964028
rect 42208 964016 42214 964028
rect 42978 964016 42984 964028
rect 42208 963988 42984 964016
rect 42208 963976 42214 963988
rect 42978 963976 42984 963988
rect 43036 963976 43042 964028
rect 673638 963296 673644 963348
rect 673696 963336 673702 963348
rect 675386 963336 675392 963348
rect 673696 963308 675392 963336
rect 673696 963296 673702 963308
rect 675386 963296 675392 963308
rect 675444 963296 675450 963348
rect 673914 962684 673920 962736
rect 673972 962724 673978 962736
rect 675478 962724 675484 962736
rect 673972 962696 675484 962724
rect 673972 962684 673978 962696
rect 675478 962684 675484 962696
rect 675536 962684 675542 962736
rect 42150 962616 42156 962668
rect 42208 962656 42214 962668
rect 42886 962656 42892 962668
rect 42208 962628 42892 962656
rect 42208 962616 42214 962628
rect 42886 962616 42892 962628
rect 42944 962616 42950 962668
rect 42150 962072 42156 962124
rect 42208 962112 42214 962124
rect 43070 962112 43076 962124
rect 42208 962084 43076 962112
rect 42208 962072 42214 962084
rect 43070 962072 43076 962084
rect 43128 962072 43134 962124
rect 673822 962004 673828 962056
rect 673880 962044 673886 962056
rect 675386 962044 675392 962056
rect 673880 962016 675392 962044
rect 673880 962004 673886 962016
rect 675386 962004 675392 962016
rect 675444 962004 675450 962056
rect 673730 961324 673736 961376
rect 673788 961364 673794 961376
rect 675386 961364 675392 961376
rect 673788 961336 675392 961364
rect 673788 961324 673794 961336
rect 675386 961324 675392 961336
rect 675444 961324 675450 961376
rect 48498 960508 48504 960560
rect 48556 960548 48562 960560
rect 57974 960548 57980 960560
rect 48556 960520 57980 960548
rect 48556 960508 48562 960520
rect 57974 960508 57980 960520
rect 58032 960508 58038 960560
rect 655606 960508 655612 960560
rect 655664 960548 655670 960560
rect 675018 960548 675024 960560
rect 655664 960520 675024 960548
rect 655664 960508 655670 960520
rect 675018 960508 675024 960520
rect 675076 960508 675082 960560
rect 42886 959624 42892 959676
rect 42944 959664 42950 959676
rect 43622 959664 43628 959676
rect 42944 959636 43628 959664
rect 42944 959624 42950 959636
rect 43622 959624 43628 959636
rect 43680 959624 43686 959676
rect 42058 959488 42064 959540
rect 42116 959528 42122 959540
rect 42886 959528 42892 959540
rect 42116 959500 42892 959528
rect 42116 959488 42122 959500
rect 42886 959488 42892 959500
rect 42944 959488 42950 959540
rect 42150 958876 42156 958928
rect 42208 958916 42214 958928
rect 43254 958916 43260 958928
rect 42208 958888 43260 958916
rect 42208 958876 42214 958888
rect 43254 958876 43260 958888
rect 43312 958876 43318 958928
rect 674466 958808 674472 958860
rect 674524 958848 674530 958860
rect 675386 958848 675392 958860
rect 674524 958820 675392 958848
rect 674524 958808 674530 958820
rect 675386 958808 675392 958820
rect 675444 958808 675450 958860
rect 42058 958468 42064 958520
rect 42116 958508 42122 958520
rect 43346 958508 43352 958520
rect 42116 958480 43352 958508
rect 42116 958468 42122 958480
rect 43346 958468 43352 958480
rect 43404 958468 43410 958520
rect 674282 958332 674288 958384
rect 674340 958372 674346 958384
rect 675386 958372 675392 958384
rect 674340 958344 675392 958372
rect 674340 958332 674346 958344
rect 675386 958332 675392 958344
rect 675444 958332 675450 958384
rect 42058 957720 42064 957772
rect 42116 957760 42122 957772
rect 43162 957760 43168 957772
rect 42116 957732 43168 957760
rect 42116 957720 42122 957732
rect 43162 957720 43168 957732
rect 43220 957720 43226 957772
rect 674374 957720 674380 957772
rect 674432 957760 674438 957772
rect 675478 957760 675484 957772
rect 674432 957732 675484 957760
rect 674432 957720 674438 957732
rect 675478 957720 675484 957732
rect 675536 957720 675542 957772
rect 674558 956972 674564 957024
rect 674616 957012 674622 957024
rect 675386 957012 675392 957024
rect 674616 956984 675392 957012
rect 674616 956972 674622 956984
rect 675386 956972 675392 956984
rect 675444 956972 675450 957024
rect 674650 955680 674656 955732
rect 674708 955720 674714 955732
rect 675478 955720 675484 955732
rect 674708 955692 675484 955720
rect 674708 955680 674714 955692
rect 675478 955680 675484 955692
rect 675536 955680 675542 955732
rect 675018 955476 675024 955528
rect 675076 955516 675082 955528
rect 675478 955516 675484 955528
rect 675076 955488 675484 955516
rect 675076 955476 675082 955488
rect 675478 955476 675484 955488
rect 675536 955476 675542 955528
rect 42150 955340 42156 955392
rect 42208 955380 42214 955392
rect 42702 955380 42708 955392
rect 42208 955352 42708 955380
rect 42208 955340 42214 955352
rect 42702 955340 42708 955352
rect 42760 955340 42766 955392
rect 673914 953980 673920 954032
rect 673972 954020 673978 954032
rect 674742 954020 674748 954032
rect 673972 953992 674748 954020
rect 673972 953980 673978 953992
rect 674742 953980 674748 953992
rect 674800 953980 674806 954032
rect 674742 953844 674748 953896
rect 674800 953884 674806 953896
rect 675386 953884 675392 953896
rect 674800 953856 675392 953884
rect 674800 953844 674806 953856
rect 675386 953844 675392 953856
rect 675444 953844 675450 953896
rect 674834 952144 674840 952196
rect 674892 952184 674898 952196
rect 674892 952156 675708 952184
rect 674892 952144 674898 952156
rect 674834 952008 674840 952060
rect 674892 952048 674898 952060
rect 675386 952048 675392 952060
rect 674892 952020 675392 952048
rect 674892 952008 674898 952020
rect 675386 952008 675392 952020
rect 675444 952008 675450 952060
rect 675680 951788 675708 952156
rect 675662 951736 675668 951788
rect 675720 951736 675726 951788
rect 673914 951056 673920 951108
rect 673972 951096 673978 951108
rect 675754 951096 675760 951108
rect 673972 951068 675760 951096
rect 673972 951056 673978 951068
rect 675754 951056 675760 951068
rect 675812 951056 675818 951108
rect 41966 950784 41972 950836
rect 42024 950824 42030 950836
rect 62666 950824 62672 950836
rect 42024 950796 62672 950824
rect 42024 950784 42030 950796
rect 62666 950784 62672 950796
rect 62724 950784 62730 950836
rect 673454 950580 673460 950632
rect 673512 950620 673518 950632
rect 673638 950620 673644 950632
rect 673512 950592 673644 950620
rect 673512 950580 673518 950592
rect 673638 950580 673644 950592
rect 673696 950580 673702 950632
rect 35618 949560 35624 949612
rect 35676 949600 35682 949612
rect 43622 949600 43628 949612
rect 35676 949572 43628 949600
rect 35676 949560 35682 949572
rect 43622 949560 43628 949572
rect 43680 949560 43686 949612
rect 35710 949492 35716 949544
rect 35768 949532 35774 949544
rect 42886 949532 42892 949544
rect 35768 949504 42892 949532
rect 35768 949492 35774 949504
rect 42886 949492 42892 949504
rect 42944 949492 42950 949544
rect 41506 949424 41512 949476
rect 41564 949464 41570 949476
rect 58434 949464 58440 949476
rect 41564 949436 58440 949464
rect 41564 949424 41570 949436
rect 58434 949424 58440 949436
rect 58492 949424 58498 949476
rect 41782 943032 41788 943084
rect 41840 943072 41846 943084
rect 49694 943072 49700 943084
rect 41840 943044 49700 943072
rect 41840 943032 41846 943044
rect 49694 943032 49700 943044
rect 49752 943032 49758 943084
rect 41782 942692 41788 942744
rect 41840 942732 41846 942744
rect 48498 942732 48504 942744
rect 41840 942704 48504 942732
rect 41840 942692 41846 942704
rect 48498 942692 48504 942704
rect 48556 942692 48562 942744
rect 41782 941468 41788 941520
rect 41840 941508 41846 941520
rect 46014 941508 46020 941520
rect 41840 941480 46020 941508
rect 41840 941468 41846 941480
rect 46014 941468 46020 941480
rect 46072 941468 46078 941520
rect 41782 941332 41788 941384
rect 41840 941372 41846 941384
rect 42702 941372 42708 941384
rect 41840 941344 42708 941372
rect 41840 941332 41846 941344
rect 42702 941332 42708 941344
rect 42760 941332 42766 941384
rect 41874 941196 41880 941248
rect 41932 941236 41938 941248
rect 42702 941236 42708 941248
rect 41932 941208 42708 941236
rect 41932 941196 41938 941208
rect 42702 941196 42708 941208
rect 42760 941196 42766 941248
rect 655790 938816 655796 938868
rect 655848 938856 655854 938868
rect 676214 938856 676220 938868
rect 655848 938828 676220 938856
rect 655848 938816 655854 938828
rect 676214 938816 676220 938828
rect 676272 938816 676278 938868
rect 655698 938680 655704 938732
rect 655756 938720 655762 938732
rect 676306 938720 676312 938732
rect 655756 938692 676312 938720
rect 655756 938680 655762 938692
rect 676306 938680 676312 938692
rect 676364 938680 676370 938732
rect 655514 938544 655520 938596
rect 655572 938584 655578 938596
rect 676122 938584 676128 938596
rect 655572 938556 676128 938584
rect 655572 938544 655578 938556
rect 676122 938544 676128 938556
rect 676180 938544 676186 938596
rect 49694 938340 49700 938392
rect 49752 938380 49758 938392
rect 58434 938380 58440 938392
rect 49752 938352 58440 938380
rect 49752 938340 49758 938352
rect 58434 938340 58440 938352
rect 58492 938340 58498 938392
rect 41148 936504 41154 936556
rect 41206 936544 41212 936556
rect 41690 936544 41696 936556
rect 41206 936516 41696 936544
rect 41206 936504 41212 936516
rect 41690 936504 41696 936516
rect 41748 936504 41754 936556
rect 670326 935756 670332 935808
rect 670384 935796 670390 935808
rect 676214 935796 676220 935808
rect 670384 935768 676220 935796
rect 670384 935756 670390 935768
rect 676214 935756 676220 935768
rect 676272 935756 676278 935808
rect 670142 935688 670148 935740
rect 670200 935728 670206 935740
rect 676030 935728 676036 935740
rect 670200 935700 676036 935728
rect 670200 935688 670206 935700
rect 676030 935688 676036 935700
rect 676088 935688 676094 935740
rect 649902 935620 649908 935672
rect 649960 935660 649966 935672
rect 678974 935660 678980 935672
rect 649960 935632 678980 935660
rect 649960 935620 649966 935632
rect 678974 935620 678980 935632
rect 679032 935620 679038 935672
rect 674742 935552 674748 935604
rect 674800 935592 674806 935604
rect 676030 935592 676036 935604
rect 674800 935564 676036 935592
rect 674800 935552 674806 935564
rect 676030 935552 676036 935564
rect 676088 935552 676094 935604
rect 674466 935484 674472 935536
rect 674524 935524 674530 935536
rect 676122 935524 676128 935536
rect 674524 935496 676128 935524
rect 674524 935484 674530 935496
rect 676122 935484 676128 935496
rect 676180 935484 676186 935536
rect 673638 935416 673644 935468
rect 673696 935456 673702 935468
rect 675938 935456 675944 935468
rect 673696 935428 675944 935456
rect 673696 935416 673702 935428
rect 675938 935416 675944 935428
rect 675996 935416 676002 935468
rect 673546 935348 673552 935400
rect 673604 935388 673610 935400
rect 675846 935388 675852 935400
rect 673604 935360 675852 935388
rect 673604 935348 673610 935360
rect 675846 935348 675852 935360
rect 675904 935348 675910 935400
rect 673730 935280 673736 935332
rect 673788 935320 673794 935332
rect 675938 935320 675944 935332
rect 673788 935292 675944 935320
rect 673788 935280 673794 935292
rect 675938 935280 675944 935292
rect 675996 935280 676002 935332
rect 674834 934940 674840 934992
rect 674892 934980 674898 934992
rect 676030 934980 676036 934992
rect 674892 934952 676036 934980
rect 674892 934940 674898 934952
rect 676030 934940 676036 934952
rect 676088 934940 676094 934992
rect 674650 932832 674656 932884
rect 674708 932872 674714 932884
rect 676030 932872 676036 932884
rect 674708 932844 676036 932872
rect 674708 932832 674714 932844
rect 676030 932832 676036 932844
rect 676088 932832 676094 932884
rect 674006 932764 674012 932816
rect 674064 932804 674070 932816
rect 676122 932804 676128 932816
rect 674064 932776 676128 932804
rect 674064 932764 674070 932776
rect 676122 932764 676128 932776
rect 676180 932764 676186 932816
rect 673822 932696 673828 932748
rect 673880 932736 673886 932748
rect 675938 932736 675944 932748
rect 673880 932708 675944 932736
rect 673880 932696 673886 932708
rect 675938 932696 675944 932708
rect 675996 932696 676002 932748
rect 673914 932628 673920 932680
rect 673972 932668 673978 932680
rect 676122 932668 676128 932680
rect 673972 932640 676128 932668
rect 673972 932628 673978 932640
rect 676122 932628 676128 932640
rect 676180 932628 676186 932680
rect 674282 932220 674288 932272
rect 674340 932260 674346 932272
rect 676122 932260 676128 932272
rect 674340 932232 676128 932260
rect 674340 932220 674346 932232
rect 676122 932220 676128 932232
rect 676180 932220 676186 932272
rect 41782 932016 41788 932068
rect 41840 932056 41846 932068
rect 46014 932056 46020 932068
rect 41840 932028 46020 932056
rect 41840 932016 41846 932028
rect 46014 932016 46020 932028
rect 46072 932016 46078 932068
rect 674374 931676 674380 931728
rect 674432 931716 674438 931728
rect 676030 931716 676036 931728
rect 674432 931688 676036 931716
rect 674432 931676 674438 931688
rect 676030 931676 676036 931688
rect 676088 931676 676094 931728
rect 674558 931268 674564 931320
rect 674616 931308 674622 931320
rect 676030 931308 676036 931320
rect 674616 931280 676036 931308
rect 674616 931268 674622 931280
rect 676030 931268 676036 931280
rect 676088 931268 676094 931320
rect 672074 927392 672080 927444
rect 672132 927432 672138 927444
rect 678974 927432 678980 927444
rect 672132 927404 678980 927432
rect 672132 927392 672138 927404
rect 678974 927392 678980 927404
rect 679032 927392 679038 927444
rect 654870 922224 654876 922276
rect 654928 922264 654934 922276
rect 669866 922264 669872 922276
rect 654928 922236 669872 922264
rect 654928 922224 654934 922236
rect 669866 922224 669872 922236
rect 669924 922224 669930 922276
rect 48590 921816 48596 921868
rect 48648 921856 48654 921868
rect 58434 921856 58440 921868
rect 48648 921828 58440 921856
rect 48648 921816 48654 921828
rect 58434 921816 58440 921828
rect 58492 921816 58498 921868
rect 53834 908080 53840 908132
rect 53892 908120 53898 908132
rect 59170 908120 59176 908132
rect 53892 908092 59176 908120
rect 53892 908080 53898 908092
rect 59170 908080 59176 908092
rect 59228 908080 59234 908132
rect 654870 908080 654876 908132
rect 654928 908120 654934 908132
rect 663794 908120 663800 908132
rect 654928 908092 663800 908120
rect 654928 908080 654934 908092
rect 663794 908080 663800 908092
rect 663852 908080 663858 908132
rect 53926 896996 53932 897048
rect 53984 897036 53990 897048
rect 58434 897036 58440 897048
rect 53984 897008 58440 897036
rect 53984 896996 53990 897008
rect 58434 896996 58440 897008
rect 58492 896996 58498 897048
rect 654870 895500 654876 895552
rect 654928 895540 654934 895552
rect 661126 895540 661132 895552
rect 654928 895512 661132 895540
rect 654928 895500 654934 895512
rect 661126 895500 661132 895512
rect 661184 895500 661190 895552
rect 51074 883192 51080 883244
rect 51132 883232 51138 883244
rect 58434 883232 58440 883244
rect 51132 883204 58440 883232
rect 51132 883192 51138 883204
rect 58434 883192 58440 883204
rect 58492 883192 58498 883244
rect 674650 873468 674656 873520
rect 674708 873508 674714 873520
rect 675386 873508 675392 873520
rect 674708 873480 675392 873508
rect 674708 873468 674714 873480
rect 675386 873468 675392 873480
rect 675444 873468 675450 873520
rect 674742 872652 674748 872704
rect 674800 872692 674806 872704
rect 675386 872692 675392 872704
rect 674800 872664 675392 872692
rect 674800 872652 674806 872664
rect 675386 872652 675392 872664
rect 675444 872652 675450 872704
rect 655146 870748 655152 870800
rect 655204 870788 655210 870800
rect 674926 870788 674932 870800
rect 655204 870760 674932 870788
rect 655204 870748 655210 870760
rect 674926 870748 674932 870760
rect 674984 870748 674990 870800
rect 673638 869796 673644 869848
rect 673696 869836 673702 869848
rect 675386 869836 675392 869848
rect 673696 869808 675392 869836
rect 673696 869796 673702 869808
rect 675386 869796 675392 869808
rect 675444 869796 675450 869848
rect 656802 869592 656808 869644
rect 656860 869632 656866 869644
rect 663702 869632 663708 869644
rect 656860 869604 663708 869632
rect 656860 869592 656866 869604
rect 663702 869592 663708 869604
rect 663760 869592 663766 869644
rect 50982 869388 50988 869440
rect 51040 869428 51046 869440
rect 58434 869428 58440 869440
rect 51040 869400 58440 869428
rect 51040 869388 51046 869400
rect 58434 869388 58440 869400
rect 58492 869388 58498 869440
rect 674190 868980 674196 869032
rect 674248 869020 674254 869032
rect 675386 869020 675392 869032
rect 674248 868992 675392 869020
rect 674248 868980 674254 868992
rect 675386 868980 675392 868992
rect 675444 868980 675450 869032
rect 673730 868504 673736 868556
rect 673788 868544 673794 868556
rect 675386 868544 675392 868556
rect 673788 868516 675392 868544
rect 673788 868504 673794 868516
rect 675386 868504 675392 868516
rect 675444 868504 675450 868556
rect 674282 867756 674288 867808
rect 674340 867796 674346 867808
rect 675386 867796 675392 867808
rect 674340 867768 675392 867796
rect 674340 867756 674346 867768
rect 675386 867756 675392 867768
rect 675444 867756 675450 867808
rect 673822 866464 673828 866516
rect 673880 866504 673886 866516
rect 675386 866504 675392 866516
rect 673880 866476 675392 866504
rect 673880 866464 673886 866476
rect 675386 866464 675392 866476
rect 675444 866464 675450 866516
rect 674926 866260 674932 866312
rect 674984 866300 674990 866312
rect 675386 866300 675392 866312
rect 674984 866272 675392 866300
rect 674984 866260 674990 866272
rect 675386 866260 675392 866272
rect 675444 866260 675450 866312
rect 674006 864628 674012 864680
rect 674064 864668 674070 864680
rect 675386 864668 675392 864680
rect 674064 864640 675392 864668
rect 674064 864628 674070 864640
rect 675386 864628 675392 864640
rect 675444 864628 675450 864680
rect 673914 862792 673920 862844
rect 673972 862832 673978 862844
rect 675478 862832 675484 862844
rect 673972 862804 675484 862832
rect 673972 862792 673978 862804
rect 675478 862792 675484 862804
rect 675536 862792 675542 862844
rect 48682 858372 48688 858424
rect 48740 858412 48746 858424
rect 58434 858412 58440 858424
rect 48740 858384 58440 858412
rect 48740 858372 48746 858384
rect 58434 858372 58440 858384
rect 58492 858372 58498 858424
rect 654686 855652 654692 855704
rect 654744 855692 654750 855704
rect 661034 855692 661040 855704
rect 654744 855664 661040 855692
rect 654744 855652 654750 855664
rect 661034 855652 661040 855664
rect 661092 855652 661098 855704
rect 674650 854224 674656 854276
rect 674708 854264 674714 854276
rect 675570 854264 675576 854276
rect 674708 854236 675576 854264
rect 674708 854224 674714 854236
rect 675570 854224 675576 854236
rect 675628 854224 675634 854276
rect 674742 854156 674748 854208
rect 674800 854196 674806 854208
rect 675754 854196 675760 854208
rect 674800 854168 675760 854196
rect 674800 854156 674806 854168
rect 675754 854156 675760 854168
rect 675812 854156 675818 854208
rect 48774 844568 48780 844620
rect 48832 844608 48838 844620
rect 58434 844608 58440 844620
rect 48832 844580 58440 844608
rect 48832 844568 48838 844580
rect 58434 844568 58440 844580
rect 58492 844568 58498 844620
rect 655054 841916 655060 841968
rect 655112 841956 655118 841968
rect 668762 841956 668768 841968
rect 655112 841928 668768 841956
rect 655112 841916 655118 841928
rect 668762 841916 668768 841928
rect 668820 841916 668826 841968
rect 54018 830764 54024 830816
rect 54076 830804 54082 830816
rect 57974 830804 57980 830816
rect 54076 830776 57980 830804
rect 54076 830764 54082 830776
rect 57974 830764 57980 830776
rect 58032 830764 58038 830816
rect 41782 817640 41788 817692
rect 41840 817680 41846 817692
rect 53926 817680 53932 817692
rect 41840 817652 53932 817680
rect 41840 817640 41846 817652
rect 53926 817640 53932 817652
rect 53984 817640 53990 817692
rect 41782 817300 41788 817352
rect 41840 817340 41846 817352
rect 51074 817340 51080 817352
rect 41840 817312 51080 817340
rect 41840 817300 41846 817312
rect 51074 817300 51080 817312
rect 51132 817300 51138 817352
rect 53742 817096 53748 817148
rect 53800 817136 53806 817148
rect 59170 817136 59176 817148
rect 53800 817108 59176 817136
rect 53800 817096 53806 817108
rect 59170 817096 59176 817108
rect 59228 817096 59234 817148
rect 42702 817028 42708 817080
rect 42760 817068 42766 817080
rect 62298 817068 62304 817080
rect 42760 817040 62304 817068
rect 42760 817028 42766 817040
rect 62298 817028 62304 817040
rect 62356 817028 62362 817080
rect 41148 816960 41154 817012
rect 41206 817000 41212 817012
rect 41782 817000 41788 817012
rect 41206 816972 41788 817000
rect 41206 816960 41212 816972
rect 41782 816960 41788 816972
rect 41840 817000 41846 817012
rect 62482 817000 62488 817012
rect 41840 816972 62488 817000
rect 41840 816960 41846 816972
rect 62482 816960 62488 816972
rect 62540 816960 62546 817012
rect 654134 814716 654140 814768
rect 654192 814756 654198 814768
rect 660942 814756 660948 814768
rect 654192 814728 660948 814756
rect 654192 814716 654198 814728
rect 660942 814716 660948 814728
rect 661000 814716 661006 814768
rect 41782 814240 41788 814292
rect 41840 814280 41846 814292
rect 42886 814280 42892 814292
rect 41840 814252 42892 814280
rect 41840 814240 41846 814252
rect 42886 814240 42892 814252
rect 42944 814280 42950 814292
rect 62666 814280 62672 814292
rect 42944 814252 62672 814280
rect 42944 814240 42950 814252
rect 62666 814240 62672 814252
rect 62724 814240 62730 814292
rect 41782 808664 41788 808716
rect 41840 808704 41846 808716
rect 44082 808704 44088 808716
rect 41840 808676 44088 808704
rect 41840 808664 41846 808676
rect 44082 808664 44088 808676
rect 44140 808664 44146 808716
rect 41782 808256 41788 808308
rect 41840 808296 41846 808308
rect 42610 808296 42616 808308
rect 41840 808268 42616 808296
rect 41840 808256 41846 808268
rect 42610 808256 42616 808268
rect 42668 808256 42674 808308
rect 41782 806012 41788 806064
rect 41840 806052 41846 806064
rect 42702 806052 42708 806064
rect 41840 806024 42708 806052
rect 41840 806012 41846 806024
rect 42702 806012 42708 806024
rect 42760 806012 42766 806064
rect 41966 805944 41972 805996
rect 42024 805984 42030 805996
rect 48498 805984 48504 805996
rect 42024 805956 48504 805984
rect 42024 805944 42030 805956
rect 48498 805944 48504 805956
rect 48556 805944 48562 805996
rect 51074 805944 51080 805996
rect 51132 805984 51138 805996
rect 58434 805984 58440 805996
rect 51132 805956 58440 805984
rect 51132 805944 51138 805956
rect 58434 805944 58440 805956
rect 58492 805944 58498 805996
rect 656802 803224 656808 803276
rect 656860 803264 656866 803276
rect 666462 803264 666468 803276
rect 656860 803236 666468 803264
rect 656860 803224 656866 803236
rect 666462 803224 666468 803236
rect 666520 803224 666526 803276
rect 44266 800436 44272 800488
rect 44324 800476 44330 800488
rect 48590 800476 48596 800488
rect 44324 800448 48596 800476
rect 44324 800436 44330 800448
rect 48590 800436 48596 800448
rect 48648 800436 48654 800488
rect 41874 800164 41880 800216
rect 41932 800164 41938 800216
rect 43898 800164 43904 800216
rect 43956 800204 43962 800216
rect 44082 800204 44088 800216
rect 43956 800176 44088 800204
rect 43956 800164 43962 800176
rect 44082 800164 44088 800176
rect 44140 800164 44146 800216
rect 41892 800012 41920 800164
rect 42334 800028 42340 800080
rect 42392 800068 42398 800080
rect 43898 800068 43904 800080
rect 42392 800040 43904 800068
rect 42392 800028 42398 800040
rect 43898 800028 43904 800040
rect 43956 800028 43962 800080
rect 41874 799960 41880 800012
rect 41932 799960 41938 800012
rect 42150 798124 42156 798176
rect 42208 798164 42214 798176
rect 42886 798164 42892 798176
rect 42208 798136 42892 798164
rect 42208 798124 42214 798136
rect 42886 798124 42892 798136
rect 42944 798124 42950 798176
rect 43898 798164 43904 798176
rect 43824 798136 43904 798164
rect 42886 797988 42892 798040
rect 42944 798028 42950 798040
rect 43346 798028 43352 798040
rect 42944 798000 43352 798028
rect 42944 797988 42950 798000
rect 43346 797988 43352 798000
rect 43404 797988 43410 798040
rect 42610 797852 42616 797904
rect 42668 797892 42674 797904
rect 42668 797864 42748 797892
rect 42668 797852 42674 797864
rect 42426 797580 42432 797632
rect 42484 797620 42490 797632
rect 42720 797620 42748 797864
rect 43346 797852 43352 797904
rect 43404 797892 43410 797904
rect 43714 797892 43720 797904
rect 43404 797864 43720 797892
rect 43404 797852 43410 797864
rect 43714 797852 43720 797864
rect 43772 797852 43778 797904
rect 43714 797716 43720 797768
rect 43772 797756 43778 797768
rect 43824 797756 43852 798136
rect 43898 798124 43904 798136
rect 43956 798124 43962 798176
rect 43898 797988 43904 798040
rect 43956 798028 43962 798040
rect 44174 798028 44180 798040
rect 43956 798000 44180 798028
rect 43956 797988 43962 798000
rect 44174 797988 44180 798000
rect 44232 797988 44238 798040
rect 43772 797728 43852 797756
rect 43772 797716 43778 797728
rect 42484 797592 42748 797620
rect 42484 797580 42490 797592
rect 42150 797240 42156 797292
rect 42208 797280 42214 797292
rect 44266 797280 44272 797292
rect 42208 797252 44272 797280
rect 42208 797240 42214 797252
rect 44266 797240 44272 797252
rect 44324 797240 44330 797292
rect 42150 796288 42156 796340
rect 42208 796328 42214 796340
rect 43070 796328 43076 796340
rect 42208 796300 43076 796328
rect 42208 796288 42214 796300
rect 43070 796288 43076 796300
rect 43128 796288 43134 796340
rect 674742 796288 674748 796340
rect 674800 796328 674806 796340
rect 675754 796328 675760 796340
rect 674800 796300 675760 796328
rect 674800 796288 674806 796300
rect 675754 796288 675760 796300
rect 675812 796288 675818 796340
rect 674558 796220 674564 796272
rect 674616 796260 674622 796272
rect 675570 796260 675576 796272
rect 674616 796232 675576 796260
rect 674616 796220 674622 796232
rect 675570 796220 675576 796232
rect 675628 796220 675634 796272
rect 43070 796152 43076 796204
rect 43128 796192 43134 796204
rect 44082 796192 44088 796204
rect 43128 796164 44088 796192
rect 43128 796152 43134 796164
rect 44082 796152 44088 796164
rect 44140 796152 44146 796204
rect 42150 794996 42156 795048
rect 42208 795036 42214 795048
rect 42702 795036 42708 795048
rect 42208 795008 42708 795036
rect 42208 794996 42214 795008
rect 42702 794996 42708 795008
rect 42760 794996 42766 795048
rect 42150 794248 42156 794300
rect 42208 794288 42214 794300
rect 43254 794288 43260 794300
rect 42208 794260 43260 794288
rect 42208 794248 42214 794260
rect 43254 794248 43260 794260
rect 43312 794248 43318 794300
rect 42150 793772 42156 793824
rect 42208 793812 42214 793824
rect 42426 793812 42432 793824
rect 42208 793784 42432 793812
rect 42208 793772 42214 793784
rect 42426 793772 42432 793784
rect 42484 793772 42490 793824
rect 42150 792956 42156 793008
rect 42208 792996 42214 793008
rect 43898 792996 43904 793008
rect 42208 792968 43904 792996
rect 42208 792956 42214 792968
rect 43898 792956 43904 792968
rect 43956 792956 43962 793008
rect 51258 792140 51264 792192
rect 51316 792180 51322 792192
rect 58066 792180 58072 792192
rect 51316 792152 58072 792180
rect 51316 792140 51322 792152
rect 58066 792140 58072 792152
rect 58124 792140 58130 792192
rect 42150 790644 42156 790696
rect 42208 790684 42214 790696
rect 43622 790684 43628 790696
rect 42208 790656 43628 790684
rect 42208 790644 42214 790656
rect 43622 790644 43628 790656
rect 43680 790644 43686 790696
rect 42150 790100 42156 790152
rect 42208 790140 42214 790152
rect 43990 790140 43996 790152
rect 42208 790112 43996 790140
rect 42208 790100 42214 790112
rect 43990 790100 43996 790112
rect 44048 790100 44054 790152
rect 42150 789420 42156 789472
rect 42208 789460 42214 789472
rect 43162 789460 43168 789472
rect 42208 789432 43168 789460
rect 42208 789420 42214 789432
rect 43162 789420 43168 789432
rect 43220 789420 43226 789472
rect 655054 789352 655060 789404
rect 655112 789392 655118 789404
rect 663886 789392 663892 789404
rect 655112 789364 663892 789392
rect 655112 789352 655118 789364
rect 663886 789352 663892 789364
rect 663944 789352 663950 789404
rect 42150 788808 42156 788860
rect 42208 788848 42214 788860
rect 43530 788848 43536 788860
rect 42208 788820 43536 788848
rect 42208 788808 42214 788820
rect 43530 788808 43536 788820
rect 43588 788808 43594 788860
rect 42150 786972 42156 787024
rect 42208 787012 42214 787024
rect 42978 787012 42984 787024
rect 42208 786984 42984 787012
rect 42208 786972 42214 786984
rect 42978 786972 42984 786984
rect 43036 786972 43042 787024
rect 42058 786224 42064 786276
rect 42116 786264 42122 786276
rect 43070 786264 43076 786276
rect 42116 786236 43076 786264
rect 42116 786224 42122 786236
rect 43070 786224 43076 786236
rect 43128 786224 43134 786276
rect 42150 785612 42156 785664
rect 42208 785652 42214 785664
rect 43438 785652 43444 785664
rect 42208 785624 43444 785652
rect 42208 785612 42214 785624
rect 43438 785612 43444 785624
rect 43496 785612 43502 785664
rect 673454 784932 673460 784984
rect 673512 784972 673518 784984
rect 675386 784972 675392 784984
rect 673512 784944 675392 784972
rect 673512 784932 673518 784944
rect 675386 784932 675392 784944
rect 675444 784932 675450 784984
rect 673546 782892 673552 782944
rect 673604 782932 673610 782944
rect 675478 782932 675484 782944
rect 673604 782904 675484 782932
rect 673604 782892 673610 782904
rect 675478 782892 675484 782904
rect 675536 782892 675542 782944
rect 655514 782416 655520 782468
rect 655572 782456 655578 782468
rect 674650 782456 674656 782468
rect 655572 782428 674656 782456
rect 655572 782416 655578 782428
rect 674650 782416 674656 782428
rect 674708 782416 674714 782468
rect 674282 780580 674288 780632
rect 674340 780620 674346 780632
rect 675478 780620 675484 780632
rect 674340 780592 675484 780620
rect 674340 780580 674346 780592
rect 675478 780580 675484 780592
rect 675536 780580 675542 780632
rect 674466 779764 674472 779816
rect 674524 779804 674530 779816
rect 675478 779804 675484 779816
rect 674524 779776 675484 779804
rect 674524 779764 674530 779776
rect 675478 779764 675484 779776
rect 675536 779764 675542 779816
rect 674190 779288 674196 779340
rect 674248 779328 674254 779340
rect 675386 779328 675392 779340
rect 674248 779300 675392 779328
rect 674248 779288 674254 779300
rect 675386 779288 675392 779300
rect 675444 779288 675450 779340
rect 674374 778744 674380 778796
rect 674432 778784 674438 778796
rect 674742 778784 674748 778796
rect 674432 778756 674748 778784
rect 674432 778744 674438 778756
rect 674742 778744 674748 778756
rect 674800 778744 674806 778796
rect 674742 778608 674748 778660
rect 674800 778648 674806 778660
rect 675478 778648 675484 778660
rect 674800 778620 675484 778648
rect 674800 778608 674806 778620
rect 675478 778608 675484 778620
rect 675536 778608 675542 778660
rect 48590 778336 48596 778388
rect 48648 778376 48654 778388
rect 58434 778376 58440 778388
rect 48648 778348 58440 778376
rect 48648 778336 48654 778348
rect 58434 778336 58440 778348
rect 58492 778336 58498 778388
rect 674374 777316 674380 777368
rect 674432 777356 674438 777368
rect 675386 777356 675392 777368
rect 674432 777328 675392 777356
rect 674432 777316 674438 777328
rect 675386 777316 675392 777328
rect 675444 777316 675450 777368
rect 674650 777044 674656 777096
rect 674708 777084 674714 777096
rect 675386 777084 675392 777096
rect 674708 777056 675392 777084
rect 674708 777044 674714 777056
rect 675386 777044 675392 777056
rect 675444 777044 675450 777096
rect 674558 775480 674564 775532
rect 674616 775520 674622 775532
rect 675386 775520 675392 775532
rect 674616 775492 675392 775520
rect 674616 775480 674622 775492
rect 675386 775480 675392 775492
rect 675444 775480 675450 775532
rect 41506 774732 41512 774784
rect 41564 774772 41570 774784
rect 48774 774772 48780 774784
rect 41564 774744 48780 774772
rect 41564 774732 41570 774744
rect 48774 774732 48780 774744
rect 48832 774732 48838 774784
rect 41506 774392 41512 774444
rect 41564 774432 41570 774444
rect 54018 774432 54024 774444
rect 41564 774404 54024 774432
rect 41564 774392 41570 774404
rect 54018 774392 54024 774404
rect 54076 774392 54082 774444
rect 41506 773916 41512 773968
rect 41564 773956 41570 773968
rect 48682 773956 48688 773968
rect 41564 773928 48688 773956
rect 41564 773916 41570 773928
rect 48682 773916 48688 773928
rect 48740 773916 48746 773968
rect 674650 773848 674656 773900
rect 674708 773888 674714 773900
rect 675202 773888 675208 773900
rect 674708 773860 675208 773888
rect 674708 773848 674714 773860
rect 675202 773848 675208 773860
rect 675260 773848 675266 773900
rect 674650 773576 674656 773628
rect 674708 773616 674714 773628
rect 675478 773616 675484 773628
rect 674708 773588 675484 773616
rect 674708 773576 674714 773588
rect 675478 773576 675484 773588
rect 675536 773576 675542 773628
rect 674466 773372 674472 773424
rect 674524 773412 674530 773424
rect 675662 773412 675668 773424
rect 674524 773384 675668 773412
rect 674524 773372 674530 773384
rect 675662 773372 675668 773384
rect 675720 773372 675726 773424
rect 675202 773304 675208 773356
rect 675260 773344 675266 773356
rect 675570 773344 675576 773356
rect 675260 773316 675576 773344
rect 675260 773304 675266 773316
rect 675570 773304 675576 773316
rect 675628 773304 675634 773356
rect 674742 773100 674748 773152
rect 674800 773140 674806 773152
rect 675478 773140 675484 773152
rect 674800 773112 675484 773140
rect 674800 773100 674806 773112
rect 675478 773100 675484 773112
rect 675536 773100 675542 773152
rect 42886 772828 42892 772880
rect 42944 772868 42950 772880
rect 62850 772868 62856 772880
rect 42944 772840 62856 772868
rect 42944 772828 42950 772840
rect 62850 772828 62856 772840
rect 62908 772828 62914 772880
rect 42058 772760 42064 772812
rect 42116 772800 42122 772812
rect 62390 772800 62396 772812
rect 42116 772772 62396 772800
rect 42116 772760 42122 772772
rect 62390 772760 62396 772772
rect 62448 772760 62454 772812
rect 674282 770516 674288 770568
rect 674340 770556 674346 770568
rect 674558 770556 674564 770568
rect 674340 770528 674564 770556
rect 674340 770516 674346 770528
rect 674558 770516 674564 770528
rect 674616 770516 674622 770568
rect 673546 770244 673552 770296
rect 673604 770284 673610 770296
rect 674190 770284 674196 770296
rect 673604 770256 674196 770284
rect 673604 770244 673610 770256
rect 674190 770244 674196 770256
rect 674248 770244 674254 770296
rect 673454 770176 673460 770228
rect 673512 770216 673518 770228
rect 674282 770216 674288 770228
rect 673512 770188 674288 770216
rect 673512 770176 673518 770188
rect 674282 770176 674288 770188
rect 674340 770176 674346 770228
rect 48774 767320 48780 767372
rect 48832 767360 48838 767372
rect 58434 767360 58440 767372
rect 48832 767332 58440 767360
rect 48832 767320 48838 767332
rect 58434 767320 58440 767332
rect 58492 767320 58498 767372
rect 43622 766368 43628 766420
rect 43680 766408 43686 766420
rect 43898 766408 43904 766420
rect 43680 766380 43904 766408
rect 43680 766368 43686 766380
rect 43898 766368 43904 766380
rect 43956 766368 43962 766420
rect 43622 766232 43628 766284
rect 43680 766272 43686 766284
rect 44082 766272 44088 766284
rect 43680 766244 44088 766272
rect 43680 766232 43686 766244
rect 44082 766232 44088 766244
rect 44140 766232 44146 766284
rect 43254 766096 43260 766148
rect 43312 766136 43318 766148
rect 44082 766136 44088 766148
rect 43312 766108 44088 766136
rect 43312 766096 43318 766108
rect 44082 766096 44088 766108
rect 44140 766096 44146 766148
rect 41506 762832 41512 762884
rect 41564 762872 41570 762884
rect 46290 762872 46296 762884
rect 41564 762844 46296 762872
rect 41564 762832 41570 762844
rect 46290 762832 46296 762844
rect 46348 762832 46354 762884
rect 654778 762764 654784 762816
rect 654836 762804 654842 762816
rect 668854 762804 668860 762816
rect 654836 762776 668860 762804
rect 654836 762764 654842 762776
rect 668854 762764 668860 762776
rect 668912 762764 668918 762816
rect 41782 760520 41788 760572
rect 41840 760560 41846 760572
rect 50982 760560 50988 760572
rect 41840 760532 50988 760560
rect 41840 760520 41846 760532
rect 50982 760520 50988 760532
rect 51040 760520 51046 760572
rect 669866 759568 669872 759620
rect 669924 759608 669930 759620
rect 676214 759608 676220 759620
rect 669924 759580 676220 759608
rect 669924 759568 669930 759580
rect 676214 759568 676220 759580
rect 676272 759568 676278 759620
rect 663794 759432 663800 759484
rect 663852 759472 663858 759484
rect 678974 759472 678980 759484
rect 663852 759444 678980 759472
rect 663852 759432 663858 759444
rect 678974 759432 678980 759444
rect 679032 759432 679038 759484
rect 661126 759296 661132 759348
rect 661184 759336 661190 759348
rect 676122 759336 676128 759348
rect 661184 759308 676128 759336
rect 661184 759296 661190 759308
rect 676122 759296 676128 759308
rect 676180 759296 676186 759348
rect 673362 759092 673368 759144
rect 673420 759132 673426 759144
rect 676030 759132 676036 759144
rect 673420 759104 676036 759132
rect 673420 759092 673426 759104
rect 676030 759092 676036 759104
rect 676088 759092 676094 759144
rect 670510 759024 670516 759076
rect 670568 759064 670574 759076
rect 676306 759064 676312 759076
rect 670568 759036 676312 759064
rect 670568 759024 670574 759036
rect 676306 759024 676312 759036
rect 676364 759024 676370 759076
rect 674006 758956 674012 759008
rect 674064 758996 674070 759008
rect 676030 758996 676036 759008
rect 674064 758968 676036 758996
rect 674064 758956 674070 758968
rect 676030 758956 676036 758968
rect 676088 758956 676094 759008
rect 42058 757596 42064 757648
rect 42116 757636 42122 757648
rect 42978 757636 42984 757648
rect 42116 757608 42984 757636
rect 42116 757596 42122 757608
rect 42978 757596 42984 757608
rect 43036 757596 43042 757648
rect 43438 757460 43444 757512
rect 43496 757500 43502 757512
rect 43990 757500 43996 757512
rect 43496 757472 43996 757500
rect 43496 757460 43502 757472
rect 43990 757460 43996 757472
rect 44048 757460 44054 757512
rect 42150 757392 42156 757444
rect 42208 757432 42214 757444
rect 43530 757432 43536 757444
rect 42208 757404 43536 757432
rect 42208 757392 42214 757404
rect 43530 757392 43536 757404
rect 43588 757392 43594 757444
rect 42702 757324 42708 757376
rect 42760 757364 42766 757376
rect 43990 757364 43996 757376
rect 42760 757336 43996 757364
rect 42760 757324 42766 757336
rect 43990 757324 43996 757336
rect 44048 757324 44054 757376
rect 41874 756984 41880 757036
rect 41932 756984 41938 757036
rect 41892 756764 41920 756984
rect 41874 756712 41880 756764
rect 41932 756712 41938 756764
rect 670602 756440 670608 756492
rect 670660 756480 670666 756492
rect 676214 756480 676220 756492
rect 670660 756452 676220 756480
rect 670660 756440 670666 756452
rect 676214 756440 676220 756452
rect 676272 756440 676278 756492
rect 668394 756372 668400 756424
rect 668452 756412 668458 756424
rect 676306 756412 676312 756424
rect 668452 756384 676312 756412
rect 668452 756372 668458 756384
rect 676306 756372 676312 756384
rect 676364 756372 676370 756424
rect 669958 756304 669964 756356
rect 670016 756344 670022 756356
rect 670142 756344 670148 756356
rect 670016 756316 670148 756344
rect 670016 756304 670022 756316
rect 670142 756304 670148 756316
rect 670200 756344 670206 756356
rect 676122 756344 676128 756356
rect 670200 756316 676128 756344
rect 670200 756304 670206 756316
rect 676122 756304 676128 756316
rect 676180 756304 676186 756356
rect 669866 756236 669872 756288
rect 669924 756276 669930 756288
rect 670326 756276 670332 756288
rect 669924 756248 670332 756276
rect 669924 756236 669930 756248
rect 670326 756236 670332 756248
rect 670384 756276 670390 756288
rect 678974 756276 678980 756288
rect 670384 756248 678980 756276
rect 670384 756236 670390 756248
rect 678974 756236 678980 756248
rect 679032 756236 679038 756288
rect 673914 756168 673920 756220
rect 673972 756208 673978 756220
rect 676030 756208 676036 756220
rect 673972 756180 676036 756208
rect 673972 756168 673978 756180
rect 676030 756168 676036 756180
rect 676088 756168 676094 756220
rect 673638 756100 673644 756152
rect 673696 756140 673702 756152
rect 676122 756140 676128 756152
rect 673696 756112 676128 756140
rect 673696 756100 673702 756112
rect 676122 756100 676128 756112
rect 676180 756100 676186 756152
rect 42426 755528 42432 755540
rect 42168 755500 42432 755528
rect 42168 755472 42196 755500
rect 42426 755488 42432 755500
rect 42484 755488 42490 755540
rect 42150 755420 42156 755472
rect 42208 755420 42214 755472
rect 42150 755148 42156 755200
rect 42208 755148 42214 755200
rect 42168 754928 42196 755148
rect 42150 754876 42156 754928
rect 42208 754876 42214 754928
rect 53834 753516 53840 753568
rect 53892 753556 53898 753568
rect 58342 753556 58348 753568
rect 53892 753528 58348 753556
rect 53892 753516 53898 753528
rect 58342 753516 58348 753528
rect 58400 753516 58406 753568
rect 673822 753448 673828 753500
rect 673880 753488 673886 753500
rect 676030 753488 676036 753500
rect 673880 753460 676036 753488
rect 673880 753448 673886 753460
rect 676030 753448 676036 753460
rect 676088 753448 676094 753500
rect 673730 753244 673736 753296
rect 673788 753284 673794 753296
rect 676030 753284 676036 753296
rect 673788 753256 676036 753284
rect 673788 753244 673794 753256
rect 676030 753244 676036 753256
rect 676088 753244 676094 753296
rect 42150 753040 42156 753092
rect 42208 753080 42214 753092
rect 43070 753080 43076 753092
rect 42208 753052 43076 753080
rect 42208 753040 42214 753052
rect 43070 753040 43076 753052
rect 43128 753040 43134 753092
rect 42150 751748 42156 751800
rect 42208 751788 42214 751800
rect 42886 751788 42892 751800
rect 42208 751760 42892 751788
rect 42208 751748 42214 751760
rect 42886 751748 42892 751760
rect 42944 751748 42950 751800
rect 42150 751068 42156 751120
rect 42208 751108 42214 751120
rect 43254 751108 43260 751120
rect 42208 751080 43260 751108
rect 42208 751068 42214 751080
rect 43254 751068 43260 751080
rect 43312 751068 43318 751120
rect 43254 750932 43260 750984
rect 43312 750972 43318 750984
rect 43714 750972 43720 750984
rect 43312 750944 43720 750972
rect 43312 750932 43318 750944
rect 43714 750932 43720 750944
rect 43772 750932 43778 750984
rect 42058 750592 42064 750644
rect 42116 750632 42122 750644
rect 43162 750632 43168 750644
rect 42116 750604 43168 750632
rect 42116 750592 42122 750604
rect 43162 750592 43168 750604
rect 43220 750592 43226 750644
rect 43162 750456 43168 750508
rect 43220 750496 43226 750508
rect 43990 750496 43996 750508
rect 43220 750468 43996 750496
rect 43220 750456 43226 750468
rect 43990 750456 43996 750468
rect 44048 750456 44054 750508
rect 42150 749776 42156 749828
rect 42208 749816 42214 749828
rect 43346 749816 43352 749828
rect 42208 749788 43352 749816
rect 42208 749776 42214 749788
rect 43346 749776 43352 749788
rect 43404 749776 43410 749828
rect 672166 749776 672172 749828
rect 672224 749816 672230 749828
rect 678974 749816 678980 749828
rect 672224 749788 678980 749816
rect 672224 749776 672230 749788
rect 678974 749776 678980 749788
rect 679032 749776 679038 749828
rect 42610 749640 42616 749692
rect 42668 749680 42674 749692
rect 43346 749680 43352 749692
rect 42668 749652 43352 749680
rect 42668 749640 42674 749652
rect 43346 749640 43352 749652
rect 43404 749640 43410 749692
rect 654870 748960 654876 749012
rect 654928 749000 654934 749012
rect 668670 749000 668676 749012
rect 654928 748972 668676 749000
rect 654928 748960 654934 748972
rect 668670 748960 668676 748972
rect 668728 748960 668734 749012
rect 42150 746920 42156 746972
rect 42208 746960 42214 746972
rect 43254 746960 43260 746972
rect 42208 746932 43260 746960
rect 42208 746920 42214 746932
rect 43254 746920 43260 746932
rect 43312 746920 43318 746972
rect 42150 746716 42156 746768
rect 42208 746756 42214 746768
rect 43346 746756 43352 746768
rect 42208 746728 43352 746756
rect 42208 746716 42214 746728
rect 43346 746716 43352 746728
rect 43404 746716 43410 746768
rect 42150 746240 42156 746292
rect 42208 746280 42214 746292
rect 43162 746280 43168 746292
rect 42208 746252 43168 746280
rect 42208 746240 42214 746252
rect 43162 746240 43168 746252
rect 43220 746240 43226 746292
rect 42150 745424 42156 745476
rect 42208 745464 42214 745476
rect 43622 745464 43628 745476
rect 42208 745436 43628 745464
rect 42208 745424 42214 745436
rect 43622 745424 43628 745436
rect 43680 745424 43686 745476
rect 42150 743724 42156 743776
rect 42208 743764 42214 743776
rect 43438 743764 43444 743776
rect 42208 743736 43444 743764
rect 42208 743724 42214 743736
rect 43438 743724 43444 743736
rect 43496 743724 43502 743776
rect 42150 743044 42156 743096
rect 42208 743084 42214 743096
rect 43898 743084 43904 743096
rect 42208 743056 43904 743084
rect 42208 743044 42214 743056
rect 43898 743044 43904 743056
rect 43956 743044 43962 743096
rect 42150 742568 42156 742620
rect 42208 742608 42214 742620
rect 43990 742608 43996 742620
rect 42208 742580 43996 742608
rect 42208 742568 42214 742580
rect 43990 742568 43996 742580
rect 44048 742568 44054 742620
rect 48682 739712 48688 739764
rect 48740 739752 48746 739764
rect 58434 739752 58440 739764
rect 48740 739724 58440 739752
rect 48740 739712 48746 739724
rect 58434 739712 58440 739724
rect 58492 739712 58498 739764
rect 673914 738420 673920 738472
rect 673972 738460 673978 738472
rect 674650 738460 674656 738472
rect 673972 738432 674656 738460
rect 673972 738420 673978 738432
rect 674650 738420 674656 738432
rect 674708 738420 674714 738472
rect 655514 738284 655520 738336
rect 655572 738324 655578 738336
rect 674650 738324 674656 738336
rect 655572 738296 674656 738324
rect 655572 738284 655578 738296
rect 674650 738284 674656 738296
rect 674708 738284 674714 738336
rect 654778 735972 654784 736024
rect 654836 736012 654842 736024
rect 661126 736012 661132 736024
rect 654836 735984 661132 736012
rect 654836 735972 654842 735984
rect 661126 735972 661132 735984
rect 661184 735972 661190 736024
rect 674006 735428 674012 735480
rect 674064 735468 674070 735480
rect 675386 735468 675392 735480
rect 674064 735440 675392 735468
rect 674064 735428 674070 735440
rect 675386 735428 675392 735440
rect 675444 735428 675450 735480
rect 673638 734952 673644 735004
rect 673696 734992 673702 735004
rect 675386 734992 675392 735004
rect 673696 734964 675392 734992
rect 673696 734952 673702 734964
rect 675386 734952 675392 734964
rect 675444 734952 675450 735004
rect 673822 734340 673828 734392
rect 673880 734380 673886 734392
rect 675386 734380 675392 734392
rect 673880 734352 675392 734380
rect 673880 734340 673886 734352
rect 675386 734340 675392 734352
rect 675444 734340 675450 734392
rect 673546 733592 673552 733644
rect 673604 733632 673610 733644
rect 675386 733632 675392 733644
rect 673604 733604 675392 733632
rect 673604 733592 673610 733604
rect 675386 733592 675392 733604
rect 675444 733592 675450 733644
rect 673730 732300 673736 732352
rect 673788 732340 673794 732352
rect 675386 732340 675392 732352
rect 673788 732312 675392 732340
rect 673788 732300 673794 732312
rect 675386 732300 675392 732312
rect 675444 732300 675450 732352
rect 674650 732028 674656 732080
rect 674708 732068 674714 732080
rect 675386 732068 675392 732080
rect 674708 732040 675392 732068
rect 674708 732028 674714 732040
rect 675386 732028 675392 732040
rect 675444 732028 675450 732080
rect 674006 731892 674012 731944
rect 674064 731932 674070 731944
rect 674650 731932 674656 731944
rect 674064 731904 674656 731932
rect 674064 731892 674070 731904
rect 674650 731892 674656 731904
rect 674708 731892 674714 731944
rect 673914 731824 673920 731876
rect 673972 731824 673978 731876
rect 673932 731604 673960 731824
rect 673914 731552 673920 731604
rect 673972 731552 673978 731604
rect 673638 730464 673644 730516
rect 673696 730504 673702 730516
rect 675386 730504 675392 730516
rect 673696 730476 675392 730504
rect 673696 730464 673702 730476
rect 675386 730464 675392 730476
rect 675444 730464 675450 730516
rect 41506 729648 41512 729700
rect 41564 729688 41570 729700
rect 43530 729688 43536 729700
rect 41564 729660 43536 729688
rect 41564 729648 41570 729660
rect 43530 729648 43536 729660
rect 43588 729648 43594 729700
rect 42518 729512 42524 729564
rect 42576 729552 42582 729564
rect 43070 729552 43076 729564
rect 42576 729524 43076 729552
rect 42576 729512 42582 729524
rect 43070 729512 43076 729524
rect 43128 729512 43134 729564
rect 41782 728832 41788 728884
rect 41840 728872 41846 728884
rect 44358 728872 44364 728884
rect 41840 728844 44364 728872
rect 41840 728832 41846 728844
rect 44358 728832 44364 728844
rect 44416 728832 44422 728884
rect 42518 728696 42524 728748
rect 42576 728736 42582 728748
rect 62390 728736 62396 728748
rect 42576 728708 62396 728736
rect 42576 728696 42582 728708
rect 62390 728696 62396 728708
rect 62448 728696 62454 728748
rect 675662 728628 675668 728680
rect 675720 728628 675726 728680
rect 675680 728408 675708 728628
rect 675662 728356 675668 728408
rect 675720 728356 675726 728408
rect 51166 725908 51172 725960
rect 51224 725948 51230 725960
rect 58434 725948 58440 725960
rect 51224 725920 58440 725948
rect 51224 725908 51230 725920
rect 58434 725908 58440 725920
rect 58492 725908 58498 725960
rect 673362 723120 673368 723172
rect 673420 723160 673426 723172
rect 678974 723160 678980 723172
rect 673420 723132 678980 723160
rect 673420 723120 673426 723132
rect 678974 723120 678980 723132
rect 679032 723120 679038 723172
rect 41506 719584 41512 719636
rect 41564 719624 41570 719636
rect 48590 719624 48596 719636
rect 41564 719596 48596 719624
rect 41564 719584 41570 719596
rect 48590 719584 48596 719596
rect 48648 719584 48654 719636
rect 674190 718088 674196 718140
rect 674248 718128 674254 718140
rect 674834 718128 674840 718140
rect 674248 718100 674840 718128
rect 674248 718088 674254 718100
rect 674834 718088 674840 718100
rect 674892 718088 674898 718140
rect 673914 717952 673920 718004
rect 673972 717992 673978 718004
rect 674190 717992 674196 718004
rect 673972 717964 674196 717992
rect 673972 717952 673978 717964
rect 674190 717952 674196 717964
rect 674248 717952 674254 718004
rect 673638 717612 673644 717664
rect 673696 717652 673702 717664
rect 673914 717652 673920 717664
rect 673696 717624 673920 717652
rect 673696 717612 673702 717624
rect 673914 717612 673920 717624
rect 673972 717612 673978 717664
rect 41322 717544 41328 717596
rect 41380 717584 41386 717596
rect 43714 717584 43720 717596
rect 41380 717556 43720 717584
rect 41380 717544 41386 717556
rect 43714 717544 43720 717556
rect 43772 717544 43778 717596
rect 42518 716592 42524 716644
rect 42576 716632 42582 716644
rect 53742 716632 53748 716644
rect 42576 716604 53748 716632
rect 42576 716592 42582 716604
rect 53742 716592 53748 716604
rect 53800 716592 53806 716644
rect 663702 716116 663708 716168
rect 663760 716156 663766 716168
rect 675938 716156 675944 716168
rect 663760 716128 675944 716156
rect 663760 716116 663766 716128
rect 675938 716116 675944 716128
rect 675996 716116 676002 716168
rect 668762 715708 668768 715760
rect 668820 715748 668826 715760
rect 675938 715748 675944 715760
rect 668820 715720 675944 715748
rect 668820 715708 668826 715720
rect 675938 715708 675944 715720
rect 675996 715708 676002 715760
rect 670510 715300 670516 715352
rect 670568 715340 670574 715352
rect 675938 715340 675944 715352
rect 670568 715312 675944 715340
rect 670568 715300 670574 715312
rect 675938 715300 675944 715312
rect 675996 715300 676002 715352
rect 661034 714960 661040 715012
rect 661092 715000 661098 715012
rect 676030 715000 676036 715012
rect 661092 714972 676036 715000
rect 661092 714960 661098 714972
rect 676030 714960 676036 714972
rect 676088 714960 676094 715012
rect 670142 714892 670148 714944
rect 670200 714932 670206 714944
rect 670510 714932 670516 714944
rect 670200 714904 670516 714932
rect 670200 714892 670206 714904
rect 670510 714892 670516 714904
rect 670568 714892 670574 714944
rect 50982 714824 50988 714876
rect 51040 714864 51046 714876
rect 58434 714864 58440 714876
rect 51040 714836 58440 714864
rect 51040 714824 51046 714836
rect 58434 714824 58440 714836
rect 58492 714824 58498 714876
rect 670234 714824 670240 714876
rect 670292 714864 670298 714876
rect 676030 714864 676036 714876
rect 670292 714836 676036 714864
rect 670292 714824 670298 714836
rect 676030 714824 676036 714836
rect 676088 714824 676094 714876
rect 673086 714008 673092 714060
rect 673144 714048 673150 714060
rect 676030 714048 676036 714060
rect 673144 714020 676036 714048
rect 673144 714008 673150 714020
rect 676030 714008 676036 714020
rect 676088 714008 676094 714060
rect 41874 713804 41880 713856
rect 41932 713804 41938 713856
rect 41892 713584 41920 713804
rect 668394 713668 668400 713720
rect 668452 713708 668458 713720
rect 670326 713708 670332 713720
rect 668452 713680 670332 713708
rect 668452 713668 668458 713680
rect 670326 713668 670332 713680
rect 670384 713708 670390 713720
rect 676030 713708 676036 713720
rect 670384 713680 676036 713708
rect 670384 713668 670390 713680
rect 676030 713668 676036 713680
rect 676088 713668 676094 713720
rect 41874 713532 41880 713584
rect 41932 713532 41938 713584
rect 668946 713192 668952 713244
rect 669004 713232 669010 713244
rect 670510 713232 670516 713244
rect 669004 713204 670516 713232
rect 669004 713192 669010 713204
rect 670510 713192 670516 713204
rect 670568 713232 670574 713244
rect 676030 713232 676036 713244
rect 670568 713204 676036 713232
rect 670568 713192 670574 713204
rect 676030 713192 676036 713204
rect 676088 713192 676094 713244
rect 668762 712784 668768 712836
rect 668820 712824 668826 712836
rect 670602 712824 670608 712836
rect 668820 712796 670608 712824
rect 668820 712784 668826 712796
rect 670602 712784 670608 712796
rect 670660 712824 670666 712836
rect 676030 712824 676036 712836
rect 670660 712796 676036 712824
rect 670660 712784 670666 712796
rect 676030 712784 676036 712796
rect 676088 712784 676094 712836
rect 669038 712376 669044 712428
rect 669096 712416 669102 712428
rect 676030 712416 676036 712428
rect 669096 712388 676036 712416
rect 669096 712376 669102 712388
rect 676030 712376 676036 712388
rect 676088 712376 676094 712428
rect 674742 712036 674748 712088
rect 674800 712076 674806 712088
rect 676030 712076 676036 712088
rect 674800 712048 676036 712076
rect 674800 712036 674806 712048
rect 676030 712036 676036 712048
rect 676088 712036 676094 712088
rect 674558 711968 674564 712020
rect 674616 712008 674622 712020
rect 675938 712008 675944 712020
rect 674616 711980 675944 712008
rect 674616 711968 674622 711980
rect 675938 711968 675944 711980
rect 675996 711968 676002 712020
rect 674282 711900 674288 711952
rect 674340 711940 674346 711952
rect 675846 711940 675852 711952
rect 674340 711912 675852 711940
rect 674340 711900 674346 711912
rect 675846 711900 675852 711912
rect 675904 711900 675910 711952
rect 674190 711832 674196 711884
rect 674248 711872 674254 711884
rect 675754 711872 675760 711884
rect 674248 711844 675760 711872
rect 674248 711832 674254 711844
rect 675754 711832 675760 711844
rect 675812 711832 675818 711884
rect 42150 711628 42156 711680
rect 42208 711668 42214 711680
rect 42886 711668 42892 711680
rect 42208 711640 42892 711668
rect 42208 711628 42214 711640
rect 42886 711628 42892 711640
rect 42944 711628 42950 711680
rect 42978 711356 42984 711408
rect 43036 711396 43042 711408
rect 43622 711396 43628 711408
rect 43036 711368 43628 711396
rect 43036 711356 43042 711368
rect 43622 711356 43628 711368
rect 43680 711356 43686 711408
rect 42150 711084 42156 711136
rect 42208 711124 42214 711136
rect 42518 711124 42524 711136
rect 42208 711096 42524 711124
rect 42208 711084 42214 711096
rect 42518 711084 42524 711096
rect 42576 711084 42582 711136
rect 673822 710812 673828 710864
rect 673880 710852 673886 710864
rect 675478 710852 675484 710864
rect 673880 710824 675484 710852
rect 673880 710812 673886 710824
rect 675478 710812 675484 710824
rect 675536 710812 675542 710864
rect 673546 710676 673552 710728
rect 673604 710716 673610 710728
rect 673822 710716 673828 710728
rect 673604 710688 673828 710716
rect 673604 710676 673610 710688
rect 673822 710676 673828 710688
rect 673880 710676 673886 710728
rect 674650 710676 674656 710728
rect 674708 710716 674714 710728
rect 675570 710716 675576 710728
rect 674708 710688 675576 710716
rect 674708 710676 674714 710688
rect 675570 710676 675576 710688
rect 675628 710676 675634 710728
rect 42150 709860 42156 709912
rect 42208 709900 42214 709912
rect 42794 709900 42800 709912
rect 42208 709872 42800 709900
rect 42208 709860 42214 709872
rect 42794 709860 42800 709872
rect 42852 709860 42858 709912
rect 42794 709724 42800 709776
rect 42852 709764 42858 709776
rect 43254 709764 43260 709776
rect 42852 709736 43260 709764
rect 42852 709724 42858 709736
rect 43254 709724 43260 709736
rect 43312 709724 43318 709776
rect 655974 709724 655980 709776
rect 656032 709764 656038 709776
rect 666922 709764 666928 709776
rect 656032 709736 666928 709764
rect 656032 709724 656038 709736
rect 666922 709724 666928 709736
rect 666980 709724 666986 709776
rect 674466 709248 674472 709300
rect 674524 709288 674530 709300
rect 676030 709288 676036 709300
rect 674524 709260 676036 709288
rect 674524 709248 674530 709260
rect 676030 709248 676036 709260
rect 676088 709248 676094 709300
rect 42150 708568 42156 708620
rect 42208 708608 42214 708620
rect 43162 708608 43168 708620
rect 42208 708580 43168 708608
rect 42208 708568 42214 708580
rect 43162 708568 43168 708580
rect 43220 708568 43226 708620
rect 674374 708228 674380 708280
rect 674432 708268 674438 708280
rect 676030 708268 676036 708280
rect 674432 708240 676036 708268
rect 674432 708228 674438 708240
rect 676030 708228 676036 708240
rect 676088 708228 676094 708280
rect 42150 708024 42156 708076
rect 42208 708064 42214 708076
rect 43898 708064 43904 708076
rect 42208 708036 43904 708064
rect 42208 708024 42214 708036
rect 43898 708024 43904 708036
rect 43956 708024 43962 708076
rect 674834 707820 674840 707872
rect 674892 707860 674898 707872
rect 676030 707860 676036 707872
rect 674892 707832 676036 707860
rect 674892 707820 674898 707832
rect 676030 707820 676036 707832
rect 676088 707820 676094 707872
rect 676030 707412 676036 707464
rect 676088 707452 676094 707464
rect 676950 707452 676956 707464
rect 676088 707424 676956 707452
rect 676088 707412 676094 707424
rect 676950 707412 676956 707424
rect 677008 707412 677014 707464
rect 42150 707344 42156 707396
rect 42208 707384 42214 707396
rect 43806 707384 43812 707396
rect 42208 707356 43812 707384
rect 42208 707344 42214 707356
rect 43806 707344 43812 707356
rect 43864 707344 43870 707396
rect 42150 706732 42156 706784
rect 42208 706772 42214 706784
rect 43254 706772 43260 706784
rect 42208 706744 43260 706772
rect 42208 706732 42214 706744
rect 43254 706732 43260 706744
rect 43312 706732 43318 706784
rect 671798 705100 671804 705152
rect 671856 705140 671862 705152
rect 676030 705140 676036 705152
rect 671856 705112 676036 705140
rect 671856 705100 671862 705112
rect 676030 705100 676036 705112
rect 676088 705100 676094 705152
rect 42242 704828 42248 704880
rect 42300 704868 42306 704880
rect 43070 704868 43076 704880
rect 42300 704840 43076 704868
rect 42300 704828 42306 704840
rect 43070 704828 43076 704840
rect 43128 704828 43134 704880
rect 42058 704216 42064 704268
rect 42116 704256 42122 704268
rect 43990 704256 43996 704268
rect 42116 704228 43996 704256
rect 42116 704216 42122 704228
rect 43990 704216 43996 704228
rect 44048 704216 44054 704268
rect 42058 702856 42064 702908
rect 42116 702896 42122 702908
rect 43714 702896 43720 702908
rect 42116 702868 43720 702896
rect 42116 702856 42122 702868
rect 43714 702856 43720 702868
rect 43772 702856 43778 702908
rect 42058 702380 42064 702432
rect 42116 702420 42122 702432
rect 43438 702420 43444 702432
rect 42116 702392 43444 702420
rect 42116 702380 42122 702392
rect 43438 702380 43444 702392
rect 43496 702380 43502 702432
rect 53742 701020 53748 701072
rect 53800 701060 53806 701072
rect 58618 701060 58624 701072
rect 53800 701032 58624 701060
rect 53800 701020 53806 701032
rect 58618 701020 58624 701032
rect 58676 701020 58682 701072
rect 42150 700408 42156 700460
rect 42208 700448 42214 700460
rect 43530 700448 43536 700460
rect 42208 700420 43536 700448
rect 42208 700408 42214 700420
rect 43530 700408 43536 700420
rect 43588 700408 43594 700460
rect 42150 700000 42156 700052
rect 42208 700040 42214 700052
rect 42886 700040 42892 700052
rect 42208 700012 42892 700040
rect 42208 700000 42214 700012
rect 42886 700000 42892 700012
rect 42944 700000 42950 700052
rect 674558 699728 674564 699780
rect 674616 699768 674622 699780
rect 675570 699768 675576 699780
rect 674616 699740 675576 699768
rect 674616 699728 674622 699740
rect 675570 699728 675576 699740
rect 675628 699728 675634 699780
rect 674742 699660 674748 699712
rect 674800 699700 674806 699712
rect 675478 699700 675484 699712
rect 674800 699672 675484 699700
rect 674800 699660 674806 699672
rect 675478 699660 675484 699672
rect 675536 699660 675542 699712
rect 674650 699592 674656 699644
rect 674708 699632 674714 699644
rect 675662 699632 675668 699644
rect 674708 699604 675668 699632
rect 674708 699592 674714 699604
rect 675662 699592 675668 699604
rect 675720 699592 675726 699644
rect 42058 699388 42064 699440
rect 42116 699428 42122 699440
rect 42794 699428 42800 699440
rect 42116 699400 42800 699428
rect 42116 699388 42122 699400
rect 42794 699388 42800 699400
rect 42852 699388 42858 699440
rect 654686 695512 654692 695564
rect 654744 695552 654750 695564
rect 663702 695552 663708 695564
rect 654744 695524 663708 695552
rect 654744 695512 654750 695524
rect 663702 695512 663708 695524
rect 663760 695512 663766 695564
rect 655514 691364 655520 691416
rect 655572 691404 655578 691416
rect 674466 691404 674472 691416
rect 655572 691376 674472 691404
rect 655572 691364 655578 691376
rect 674466 691364 674472 691376
rect 674524 691364 674530 691416
rect 673730 690412 673736 690464
rect 673788 690452 673794 690464
rect 675386 690452 675392 690464
rect 673788 690424 675392 690452
rect 673788 690412 673794 690424
rect 675386 690412 675392 690424
rect 675444 690412 675450 690464
rect 673178 689120 673184 689172
rect 673236 689160 673242 689172
rect 675478 689160 675484 689172
rect 673236 689132 675484 689160
rect 673236 689120 673242 689132
rect 675478 689120 675484 689132
rect 675536 689120 675542 689172
rect 672994 688576 673000 688628
rect 673052 688616 673058 688628
rect 675386 688616 675392 688628
rect 673052 688588 675392 688616
rect 673052 688576 673058 688588
rect 675386 688576 675392 688588
rect 675444 688576 675450 688628
rect 41506 688372 41512 688424
rect 41564 688412 41570 688424
rect 48682 688412 48688 688424
rect 41564 688384 48688 688412
rect 41564 688372 41570 688384
rect 48682 688372 48688 688384
rect 48740 688372 48746 688424
rect 41690 688032 41696 688084
rect 41748 688072 41754 688084
rect 53834 688072 53840 688084
rect 41748 688044 53840 688072
rect 41748 688032 41754 688044
rect 53834 688032 53840 688044
rect 53892 688032 53898 688084
rect 41782 687692 41788 687744
rect 41840 687732 41846 687744
rect 51166 687732 51172 687744
rect 41840 687704 51172 687732
rect 41840 687692 41846 687704
rect 51166 687692 51172 687704
rect 51224 687692 51230 687744
rect 673270 687284 673276 687336
rect 673328 687324 673334 687336
rect 675386 687324 675392 687336
rect 673328 687296 675392 687324
rect 673328 687284 673334 687296
rect 675386 687284 675392 687296
rect 675444 687284 675450 687336
rect 51074 687216 51080 687268
rect 51132 687256 51138 687268
rect 58434 687256 58440 687268
rect 51132 687228 58440 687256
rect 51132 687216 51138 687228
rect 58434 687216 58440 687228
rect 58492 687216 58498 687268
rect 674466 687012 674472 687064
rect 674524 687052 674530 687064
rect 675478 687052 675484 687064
rect 674524 687024 675484 687052
rect 674524 687012 674530 687024
rect 675478 687012 675484 687024
rect 675536 687012 675542 687064
rect 673822 685448 673828 685500
rect 673880 685488 673886 685500
rect 675386 685488 675392 685500
rect 673880 685460 675392 685488
rect 673880 685448 673886 685460
rect 675386 685448 675392 685460
rect 675444 685448 675450 685500
rect 674282 683612 674288 683664
rect 674340 683652 674346 683664
rect 675478 683652 675484 683664
rect 674340 683624 675484 683652
rect 674340 683612 674346 683624
rect 675478 683612 675484 683624
rect 675536 683612 675542 683664
rect 654870 682932 654876 682984
rect 654928 682972 654934 682984
rect 663794 682972 663800 682984
rect 654928 682944 663800 682972
rect 654928 682932 654934 682944
rect 663794 682932 663800 682944
rect 663852 682932 663858 682984
rect 42794 681640 42800 681692
rect 42852 681680 42858 681692
rect 62942 681680 62948 681692
rect 42852 681652 62948 681680
rect 42852 681640 42858 681652
rect 62942 681640 62948 681652
rect 63000 681640 63006 681692
rect 673086 678988 673092 679040
rect 673144 679028 673150 679040
rect 678974 679028 678980 679040
rect 673144 679000 678980 679028
rect 673144 678988 673150 679000
rect 678974 678988 678980 679000
rect 679032 678988 679038 679040
rect 41782 678308 41788 678360
rect 41840 678348 41846 678360
rect 44082 678348 44088 678360
rect 41840 678320 44088 678348
rect 41840 678308 41846 678320
rect 44082 678308 44088 678320
rect 44140 678308 44146 678360
rect 41782 676608 41788 676660
rect 41840 676648 41846 676660
rect 48682 676648 48688 676660
rect 41840 676620 48688 676648
rect 41840 676608 41846 676620
rect 48682 676608 48688 676620
rect 48740 676608 48746 676660
rect 48866 673480 48872 673532
rect 48924 673520 48930 673532
rect 58434 673520 58440 673532
rect 48924 673492 58440 673520
rect 48924 673480 48930 673492
rect 58434 673480 58440 673492
rect 58492 673480 58498 673532
rect 41322 673412 41328 673464
rect 41380 673452 41386 673464
rect 42886 673452 42892 673464
rect 41380 673424 42892 673452
rect 41380 673412 41386 673424
rect 42886 673412 42892 673424
rect 42944 673412 42950 673464
rect 666462 671508 666468 671560
rect 666520 671548 666526 671560
rect 676214 671548 676220 671560
rect 666520 671520 676220 671548
rect 666520 671508 666526 671520
rect 676214 671508 676220 671520
rect 676272 671508 676278 671560
rect 674742 671236 674748 671288
rect 674800 671276 674806 671288
rect 675202 671276 675208 671288
rect 674800 671248 675208 671276
rect 674800 671236 674806 671248
rect 675202 671236 675208 671248
rect 675260 671236 675266 671288
rect 660942 670760 660948 670812
rect 661000 670800 661006 670812
rect 676030 670800 676036 670812
rect 661000 670772 676036 670800
rect 661000 670760 661006 670772
rect 676030 670760 676036 670772
rect 676088 670760 676094 670812
rect 44174 670692 44180 670744
rect 44232 670732 44238 670744
rect 48774 670732 48780 670744
rect 44232 670704 48780 670732
rect 44232 670692 44238 670704
rect 48774 670692 48780 670704
rect 48832 670692 48838 670744
rect 43806 670624 43812 670676
rect 43864 670624 43870 670676
rect 43990 670624 43996 670676
rect 44048 670624 44054 670676
rect 44082 670624 44088 670676
rect 44140 670624 44146 670676
rect 41874 670556 41880 670608
rect 41932 670556 41938 670608
rect 41966 670556 41972 670608
rect 42024 670596 42030 670608
rect 42702 670596 42708 670608
rect 42024 670568 42708 670596
rect 42024 670556 42030 670568
rect 42702 670556 42708 670568
rect 42760 670556 42766 670608
rect 43824 670596 43852 670624
rect 43732 670568 43852 670596
rect 41892 670404 41920 670556
rect 41874 670352 41880 670404
rect 41932 670352 41938 670404
rect 43732 670392 43760 670568
rect 44008 670528 44036 670624
rect 43824 670500 44036 670528
rect 43824 670472 43852 670500
rect 43806 670420 43812 670472
rect 43864 670420 43870 670472
rect 43990 670420 43996 670472
rect 44048 670460 44054 670472
rect 44100 670460 44128 670624
rect 663886 670556 663892 670608
rect 663944 670596 663950 670608
rect 676030 670596 676036 670608
rect 663944 670568 676036 670596
rect 663944 670556 663950 670568
rect 676030 670556 676036 670568
rect 676088 670556 676094 670608
rect 44048 670432 44128 670460
rect 44048 670420 44054 670432
rect 43732 670364 44128 670392
rect 44100 670256 44128 670364
rect 670234 670284 670240 670336
rect 670292 670324 670298 670336
rect 676214 670324 676220 670336
rect 670292 670296 676220 670324
rect 670292 670284 670298 670296
rect 676214 670284 676220 670296
rect 676272 670284 676278 670336
rect 44100 670228 44220 670256
rect 44192 670200 44220 670228
rect 44174 670148 44180 670200
rect 44232 670148 44238 670200
rect 669130 669740 669136 669792
rect 669188 669780 669194 669792
rect 674466 669780 674472 669792
rect 669188 669752 674472 669780
rect 669188 669740 669194 669752
rect 674466 669740 674472 669752
rect 674524 669780 674530 669792
rect 676030 669780 676036 669792
rect 674524 669752 676036 669780
rect 674524 669740 674530 669752
rect 676030 669740 676036 669752
rect 676088 669740 676094 669792
rect 670510 668652 670516 668704
rect 670568 668692 670574 668704
rect 676214 668692 676220 668704
rect 670568 668664 676220 668692
rect 670568 668652 670574 668664
rect 676214 668652 676220 668664
rect 676272 668652 676278 668704
rect 42058 668448 42064 668500
rect 42116 668488 42122 668500
rect 43898 668488 43904 668500
rect 42116 668460 43904 668488
rect 42116 668448 42122 668460
rect 43898 668448 43904 668460
rect 43956 668448 43962 668500
rect 673086 668040 673092 668092
rect 673144 668080 673150 668092
rect 675938 668080 675944 668092
rect 673144 668052 675944 668080
rect 673144 668040 673150 668052
rect 675938 668040 675944 668052
rect 675996 668040 676002 668092
rect 674742 667904 674748 667956
rect 674800 667944 674806 667956
rect 676030 667944 676036 667956
rect 674800 667916 676036 667944
rect 674800 667904 674806 667916
rect 676030 667904 676036 667916
rect 676088 667904 676094 667956
rect 673914 667836 673920 667888
rect 673972 667876 673978 667888
rect 676122 667876 676128 667888
rect 673972 667848 676128 667876
rect 673972 667836 673978 667848
rect 676122 667836 676128 667848
rect 676180 667836 676186 667888
rect 674558 667768 674564 667820
rect 674616 667808 674622 667820
rect 676030 667808 676036 667820
rect 674616 667780 676036 667808
rect 674616 667768 674622 667780
rect 676030 667768 676036 667780
rect 676088 667768 676094 667820
rect 42150 667700 42156 667752
rect 42208 667740 42214 667752
rect 44082 667740 44088 667752
rect 42208 667712 44088 667740
rect 42208 667700 42214 667712
rect 44082 667700 44088 667712
rect 44140 667700 44146 667752
rect 669038 667700 669044 667752
rect 669096 667740 669102 667752
rect 675938 667740 675944 667752
rect 669096 667712 675944 667740
rect 669096 667700 669102 667712
rect 675938 667700 675944 667712
rect 675996 667700 676002 667752
rect 42150 666680 42156 666732
rect 42208 666720 42214 666732
rect 43714 666720 43720 666732
rect 42208 666692 43720 666720
rect 42208 666680 42214 666692
rect 43714 666680 43720 666692
rect 43772 666680 43778 666732
rect 42150 665388 42156 665440
rect 42208 665428 42214 665440
rect 42702 665428 42708 665440
rect 42208 665400 42708 665428
rect 42208 665388 42214 665400
rect 42702 665388 42708 665400
rect 42760 665388 42766 665440
rect 674650 665116 674656 665168
rect 674708 665156 674714 665168
rect 676030 665156 676036 665168
rect 674708 665128 676036 665156
rect 674708 665116 674714 665128
rect 676030 665116 676036 665128
rect 676088 665116 676094 665168
rect 675202 664708 675208 664760
rect 675260 664748 675266 664760
rect 676030 664748 676036 664760
rect 675260 664720 676036 664748
rect 675260 664708 675266 664720
rect 676030 664708 676036 664720
rect 676088 664708 676094 664760
rect 42150 664640 42156 664692
rect 42208 664680 42214 664692
rect 43530 664680 43536 664692
rect 42208 664652 43536 664680
rect 42208 664640 42214 664652
rect 43530 664640 43536 664652
rect 43588 664640 43594 664692
rect 42150 663960 42156 664012
rect 42208 664000 42214 664012
rect 43990 664000 43996 664012
rect 42208 663972 43996 664000
rect 42208 663960 42214 663972
rect 43990 663960 43996 663972
rect 44048 663960 44054 664012
rect 42150 663552 42156 663604
rect 42208 663592 42214 663604
rect 42886 663592 42892 663604
rect 42208 663564 42892 663592
rect 42208 663552 42214 663564
rect 42886 663552 42892 663564
rect 42944 663552 42950 663604
rect 48958 662396 48964 662448
rect 49016 662436 49022 662448
rect 58434 662436 58440 662448
rect 49016 662408 58440 662436
rect 49016 662396 49022 662408
rect 58434 662396 58440 662408
rect 58492 662396 58498 662448
rect 42150 661036 42156 661088
rect 42208 661076 42214 661088
rect 43806 661076 43812 661088
rect 42208 661048 43812 661076
rect 42208 661036 42214 661048
rect 43806 661036 43812 661048
rect 43864 661036 43870 661088
rect 42150 660492 42156 660544
rect 42208 660532 42214 660544
rect 43438 660532 43444 660544
rect 42208 660504 43444 660532
rect 42208 660492 42214 660504
rect 43438 660492 43444 660504
rect 43496 660492 43502 660544
rect 42150 659880 42156 659932
rect 42208 659920 42214 659932
rect 43254 659920 43260 659932
rect 42208 659892 43260 659920
rect 42208 659880 42214 659892
rect 43254 659880 43260 659892
rect 43312 659880 43318 659932
rect 672350 659676 672356 659728
rect 672408 659716 672414 659728
rect 678974 659716 678980 659728
rect 672408 659688 678980 659716
rect 672408 659676 672414 659688
rect 678974 659676 678980 659688
rect 679032 659676 679038 659728
rect 42150 659200 42156 659252
rect 42208 659240 42214 659252
rect 42978 659240 42984 659252
rect 42208 659212 42984 659240
rect 42208 659200 42214 659212
rect 42978 659200 42984 659212
rect 43036 659200 43042 659252
rect 42150 657228 42156 657280
rect 42208 657268 42214 657280
rect 43622 657268 43628 657280
rect 42208 657240 43628 657268
rect 42208 657228 42214 657240
rect 43622 657228 43628 657240
rect 43680 657228 43686 657280
rect 656158 657024 656164 657076
rect 656216 657064 656222 657076
rect 660942 657064 660948 657076
rect 656216 657036 660948 657064
rect 656216 657024 656222 657036
rect 660942 657024 660948 657036
rect 661000 657024 661006 657076
rect 42150 656820 42156 656872
rect 42208 656860 42214 656872
rect 44082 656860 44088 656872
rect 42208 656832 44088 656860
rect 42208 656820 42214 656832
rect 44082 656820 44088 656832
rect 44140 656820 44146 656872
rect 42150 656140 42156 656192
rect 42208 656180 42214 656192
rect 43070 656180 43076 656192
rect 42208 656152 43076 656180
rect 42208 656140 42214 656152
rect 43070 656140 43076 656152
rect 43128 656140 43134 656192
rect 673546 649544 673552 649596
rect 673604 649584 673610 649596
rect 675386 649584 675392 649596
rect 673604 649556 675392 649584
rect 673604 649544 673610 649556
rect 675386 649544 675392 649556
rect 675444 649544 675450 649596
rect 53834 648592 53840 648644
rect 53892 648632 53898 648644
rect 59170 648632 59176 648644
rect 53892 648604 59176 648632
rect 53892 648592 53898 648604
rect 59170 648592 59176 648604
rect 59228 648592 59234 648644
rect 674650 647708 674656 647760
rect 674708 647748 674714 647760
rect 675478 647748 675484 647760
rect 674708 647720 675484 647748
rect 674708 647708 674714 647720
rect 675478 647708 675484 647720
rect 675536 647708 675542 647760
rect 673454 647300 673460 647352
rect 673512 647340 673518 647352
rect 674742 647340 674748 647352
rect 673512 647312 674748 647340
rect 673512 647300 673518 647312
rect 674742 647300 674748 647312
rect 674800 647300 674806 647352
rect 655514 647164 655520 647216
rect 655572 647204 655578 647216
rect 674742 647204 674748 647216
rect 655572 647176 674748 647204
rect 655572 647164 655578 647176
rect 674742 647164 674748 647176
rect 674800 647164 674806 647216
rect 673914 645396 673920 645448
rect 673972 645436 673978 645448
rect 675386 645436 675392 645448
rect 673972 645408 675392 645436
rect 673972 645396 673978 645408
rect 675386 645396 675392 645408
rect 675444 645396 675450 645448
rect 41506 645124 41512 645176
rect 41564 645164 41570 645176
rect 51074 645164 51080 645176
rect 41564 645136 51080 645164
rect 41564 645124 41570 645136
rect 51074 645124 51080 645136
rect 51132 645124 51138 645176
rect 41506 644784 41512 644836
rect 41564 644824 41570 644836
rect 53742 644824 53748 644836
rect 41564 644796 53748 644824
rect 41564 644784 41570 644796
rect 53742 644784 53748 644796
rect 53800 644784 53806 644836
rect 674558 644784 674564 644836
rect 674616 644824 674622 644836
rect 675386 644824 675392 644836
rect 674616 644796 675392 644824
rect 674616 644784 674622 644796
rect 675386 644784 675392 644796
rect 675444 644784 675450 644836
rect 41782 644512 41788 644564
rect 41840 644552 41846 644564
rect 48866 644552 48872 644564
rect 41840 644524 48872 644552
rect 41840 644512 41846 644524
rect 48866 644512 48872 644524
rect 48924 644512 48930 644564
rect 673638 644104 673644 644156
rect 673696 644144 673702 644156
rect 675386 644144 675392 644156
rect 673696 644116 675392 644144
rect 673696 644104 673702 644116
rect 675386 644104 675392 644116
rect 675444 644104 675450 644156
rect 674374 643356 674380 643408
rect 674432 643396 674438 643408
rect 675386 643396 675392 643408
rect 674432 643368 675392 643396
rect 674432 643356 674438 643368
rect 675386 643356 675392 643368
rect 675444 643356 675450 643408
rect 654870 643084 654876 643136
rect 654928 643124 654934 643136
rect 663886 643124 663892 643136
rect 654928 643096 663892 643124
rect 654928 643084 654934 643096
rect 663886 643084 663892 643096
rect 663944 643084 663950 643136
rect 674006 642064 674012 642116
rect 674064 642104 674070 642116
rect 675386 642104 675392 642116
rect 674064 642076 675392 642104
rect 674064 642064 674070 642076
rect 675386 642064 675392 642076
rect 675444 642064 675450 642116
rect 674742 641860 674748 641912
rect 674800 641900 674806 641912
rect 675386 641900 675392 641912
rect 674800 641872 675392 641900
rect 674800 641860 674806 641872
rect 675386 641860 675392 641872
rect 675444 641860 675450 641912
rect 674190 640228 674196 640280
rect 674248 640268 674254 640280
rect 675386 640268 675392 640280
rect 674248 640240 675392 640268
rect 674248 640228 674254 640240
rect 675386 640228 675392 640240
rect 675444 640228 675450 640280
rect 674650 638800 674656 638852
rect 674708 638800 674714 638852
rect 674668 638704 674696 638800
rect 675202 638704 675208 638716
rect 674668 638676 675208 638704
rect 675202 638664 675208 638676
rect 675260 638664 675266 638716
rect 674558 638392 674564 638444
rect 674616 638432 674622 638444
rect 675478 638432 675484 638444
rect 674616 638404 675484 638432
rect 674616 638392 674622 638404
rect 675478 638392 675484 638404
rect 675536 638392 675542 638444
rect 675202 638188 675208 638240
rect 675260 638228 675266 638240
rect 675662 638228 675668 638240
rect 675260 638200 675668 638228
rect 675260 638188 675266 638200
rect 675662 638188 675668 638200
rect 675720 638188 675726 638240
rect 673086 637848 673092 637900
rect 673144 637888 673150 637900
rect 679158 637888 679164 637900
rect 673144 637860 679164 637888
rect 673144 637848 673150 637860
rect 679158 637848 679164 637860
rect 679216 637848 679222 637900
rect 673454 637508 673460 637560
rect 673512 637548 673518 637560
rect 679066 637548 679072 637560
rect 673512 637520 679072 637548
rect 673512 637508 673518 637520
rect 679066 637508 679072 637520
rect 679124 637508 679130 637560
rect 48866 634788 48872 634840
rect 48924 634828 48930 634840
rect 58434 634828 58440 634840
rect 48924 634800 58440 634828
rect 48924 634788 48930 634800
rect 58434 634788 58440 634800
rect 58492 634788 58498 634840
rect 41506 633224 41512 633276
rect 41564 633264 41570 633276
rect 48774 633264 48780 633276
rect 41564 633236 48780 633264
rect 41564 633224 41570 633236
rect 48774 633224 48780 633236
rect 48832 633224 48838 633276
rect 43622 629280 43628 629332
rect 43680 629320 43686 629332
rect 50982 629320 50988 629332
rect 43680 629292 50988 629320
rect 43680 629280 43686 629292
rect 50982 629280 50988 629292
rect 51040 629280 51046 629332
rect 655054 629280 655060 629332
rect 655112 629320 655118 629332
rect 669038 629320 669044 629332
rect 655112 629292 669044 629320
rect 655112 629280 655118 629292
rect 669038 629280 669044 629292
rect 669096 629280 669102 629332
rect 30282 627852 30288 627904
rect 30340 627892 30346 627904
rect 42518 627892 42524 627904
rect 30340 627864 42524 627892
rect 30340 627852 30346 627864
rect 42518 627852 42524 627864
rect 42576 627852 42582 627904
rect 41782 627376 41788 627428
rect 41840 627376 41846 627428
rect 41800 627088 41828 627376
rect 41782 627036 41788 627088
rect 41840 627036 41846 627088
rect 674466 626492 674472 626544
rect 674524 626532 674530 626544
rect 676030 626532 676036 626544
rect 674524 626504 676036 626532
rect 674524 626492 674530 626504
rect 676030 626492 676036 626504
rect 676088 626492 676094 626544
rect 42150 625268 42156 625320
rect 42208 625308 42214 625320
rect 43714 625308 43720 625320
rect 42208 625280 43720 625308
rect 42208 625268 42214 625280
rect 43714 625268 43720 625280
rect 43772 625268 43778 625320
rect 42150 624656 42156 624708
rect 42208 624696 42214 624708
rect 43622 624696 43628 624708
rect 42208 624668 43628 624696
rect 42208 624656 42214 624668
rect 43622 624656 43628 624668
rect 43680 624656 43686 624708
rect 668854 624112 668860 624164
rect 668912 624152 668918 624164
rect 676214 624152 676220 624164
rect 668912 624124 676220 624152
rect 668912 624112 668918 624124
rect 676214 624112 676220 624124
rect 676272 624112 676278 624164
rect 668670 623976 668676 624028
rect 668728 624016 668734 624028
rect 678974 624016 678980 624028
rect 668728 623988 678980 624016
rect 668728 623976 668734 623988
rect 678974 623976 678980 623988
rect 679032 623976 679038 624028
rect 673362 623908 673368 623960
rect 673420 623948 673426 623960
rect 676030 623948 676036 623960
rect 673420 623920 676036 623948
rect 673420 623908 673426 623920
rect 676030 623908 676036 623920
rect 676088 623908 676094 623960
rect 661126 623840 661132 623892
rect 661184 623880 661190 623892
rect 676306 623880 676312 623892
rect 661184 623852 676312 623880
rect 661184 623840 661190 623852
rect 676306 623840 676312 623852
rect 676364 623840 676370 623892
rect 51074 623772 51080 623824
rect 51132 623812 51138 623824
rect 58434 623812 58440 623824
rect 51132 623784 58440 623812
rect 51132 623772 51138 623784
rect 58434 623772 58440 623784
rect 58492 623772 58498 623824
rect 668578 623772 668584 623824
rect 668636 623812 668642 623824
rect 670602 623812 670608 623824
rect 668636 623784 670608 623812
rect 668636 623772 668642 623784
rect 670602 623772 670608 623784
rect 670660 623812 670666 623824
rect 676122 623812 676128 623824
rect 670660 623784 676128 623812
rect 670660 623772 670666 623784
rect 676122 623772 676128 623784
rect 676180 623772 676186 623824
rect 673822 623704 673828 623756
rect 673880 623744 673886 623756
rect 676030 623744 676036 623756
rect 673880 623716 676036 623744
rect 673880 623704 673886 623716
rect 676030 623704 676036 623716
rect 676088 623704 676094 623756
rect 42150 623432 42156 623484
rect 42208 623472 42214 623484
rect 43070 623472 43076 623484
rect 42208 623444 43076 623472
rect 42208 623432 42214 623444
rect 43070 623432 43076 623444
rect 43128 623432 43134 623484
rect 42058 622140 42064 622192
rect 42116 622180 42122 622192
rect 42518 622180 42524 622192
rect 42116 622152 42524 622180
rect 42116 622140 42122 622152
rect 42518 622140 42524 622152
rect 42576 622140 42582 622192
rect 42150 621460 42156 621512
rect 42208 621500 42214 621512
rect 43254 621500 43260 621512
rect 42208 621472 43260 621500
rect 42208 621460 42214 621472
rect 43254 621460 43260 621472
rect 43312 621460 43318 621512
rect 670234 621052 670240 621104
rect 670292 621092 670298 621104
rect 678974 621092 678980 621104
rect 670292 621064 678980 621092
rect 670292 621052 670298 621064
rect 678974 621052 678980 621064
rect 679032 621052 679038 621104
rect 42058 620984 42064 621036
rect 42116 621024 42122 621036
rect 43162 621024 43168 621036
rect 42116 620996 43168 621024
rect 42116 620984 42122 620996
rect 43162 620984 43168 620996
rect 43220 620984 43226 621036
rect 668486 620984 668492 621036
rect 668544 621024 668550 621036
rect 670510 621024 670516 621036
rect 668544 620996 670516 621024
rect 668544 620984 668550 620996
rect 670510 620984 670516 620996
rect 670568 621024 670574 621036
rect 676214 621024 676220 621036
rect 670568 620996 676220 621024
rect 670568 620984 670574 620996
rect 676214 620984 676220 620996
rect 676272 620984 676278 621036
rect 674282 620916 674288 620968
rect 674340 620956 674346 620968
rect 676030 620956 676036 620968
rect 674340 620928 676036 620956
rect 674340 620916 674346 620928
rect 676030 620916 676036 620928
rect 676088 620916 676094 620968
rect 673730 620848 673736 620900
rect 673788 620888 673794 620900
rect 676122 620888 676128 620900
rect 673788 620860 676128 620888
rect 673788 620848 673794 620860
rect 676122 620848 676128 620860
rect 676180 620848 676186 620900
rect 42058 620168 42064 620220
rect 42116 620208 42122 620220
rect 43898 620208 43904 620220
rect 42116 620180 43904 620208
rect 42116 620168 42122 620180
rect 43898 620168 43904 620180
rect 43956 620168 43962 620220
rect 42242 619012 42248 619064
rect 42300 619052 42306 619064
rect 42886 619052 42892 619064
rect 42300 619024 42892 619052
rect 42300 619012 42306 619024
rect 42886 619012 42892 619024
rect 42944 619012 42950 619064
rect 673270 618196 673276 618248
rect 673328 618236 673334 618248
rect 676030 618236 676036 618248
rect 673328 618208 676036 618236
rect 673328 618196 673334 618208
rect 676030 618196 676036 618208
rect 676088 618196 676094 618248
rect 673178 617924 673184 617976
rect 673236 617964 673242 617976
rect 676214 617964 676220 617976
rect 673236 617936 676220 617964
rect 673236 617924 673242 617936
rect 676214 617924 676220 617936
rect 676272 617924 676278 617976
rect 42150 617856 42156 617908
rect 42208 617896 42214 617908
rect 43806 617896 43812 617908
rect 42208 617868 43812 617896
rect 42208 617856 42214 617868
rect 43806 617856 43812 617868
rect 43864 617856 43870 617908
rect 42058 617312 42064 617364
rect 42116 617352 42122 617364
rect 43438 617352 43444 617364
rect 42116 617324 43444 617352
rect 42116 617312 42122 617324
rect 43438 617312 43444 617324
rect 43496 617312 43502 617364
rect 672994 616700 673000 616752
rect 673052 616740 673058 616752
rect 676214 616740 676220 616752
rect 673052 616712 676220 616740
rect 673052 616700 673058 616712
rect 676214 616700 676220 616712
rect 676272 616700 676278 616752
rect 42242 616020 42248 616072
rect 42300 616060 42306 616072
rect 43530 616060 43536 616072
rect 42300 616032 43536 616060
rect 42300 616020 42306 616032
rect 43530 616020 43536 616032
rect 43588 616020 43594 616072
rect 672442 614592 672448 614644
rect 672500 614632 672506 614644
rect 678974 614632 678980 614644
rect 672500 614604 678980 614632
rect 672500 614592 672506 614604
rect 678974 614592 678980 614604
rect 679032 614592 679038 614644
rect 42150 614184 42156 614236
rect 42208 614224 42214 614236
rect 43346 614224 43352 614236
rect 42208 614196 43352 614224
rect 42208 614184 42214 614196
rect 43346 614184 43352 614196
rect 43404 614184 43410 614236
rect 42150 613640 42156 613692
rect 42208 613680 42214 613692
rect 42978 613680 42984 613692
rect 42208 613652 42984 613680
rect 42208 613640 42214 613652
rect 42978 613640 42984 613652
rect 43036 613640 43042 613692
rect 42150 612960 42156 613012
rect 42208 613000 42214 613012
rect 42794 613000 42800 613012
rect 42208 612972 42800 613000
rect 42208 612960 42214 612972
rect 42794 612960 42800 612972
rect 42852 612960 42858 613012
rect 50982 609968 50988 610020
rect 51040 610008 51046 610020
rect 58434 610008 58440 610020
rect 51040 609980 58440 610008
rect 51040 609968 51046 609980
rect 58434 609968 58440 609980
rect 58492 609968 58498 610020
rect 674466 608744 674472 608796
rect 674524 608784 674530 608796
rect 675662 608784 675668 608796
rect 674524 608756 675668 608784
rect 674524 608744 674530 608756
rect 675662 608744 675668 608756
rect 675720 608744 675726 608796
rect 654594 603032 654600 603084
rect 654652 603072 654658 603084
rect 674650 603072 674656 603084
rect 654652 603044 674656 603072
rect 654652 603032 654658 603044
rect 674650 603032 674656 603044
rect 674708 603032 674714 603084
rect 654318 602148 654324 602200
rect 654376 602188 654382 602200
rect 661034 602188 661040 602200
rect 654376 602160 661040 602188
rect 654376 602148 654382 602160
rect 661034 602148 661040 602160
rect 661092 602148 661098 602200
rect 41506 601876 41512 601928
rect 41564 601916 41570 601928
rect 48866 601916 48872 601928
rect 41564 601888 48872 601916
rect 41564 601876 41570 601888
rect 48866 601876 48872 601888
rect 48924 601876 48930 601928
rect 674282 600380 674288 600432
rect 674340 600420 674346 600432
rect 675478 600420 675484 600432
rect 674340 600392 675484 600420
rect 674340 600380 674346 600392
rect 675478 600380 675484 600392
rect 675536 600380 675542 600432
rect 674742 599564 674748 599616
rect 674800 599604 674806 599616
rect 675478 599604 675484 599616
rect 674800 599576 675484 599604
rect 674800 599564 674806 599576
rect 675478 599564 675484 599576
rect 675536 599564 675542 599616
rect 673730 598952 673736 599004
rect 673788 598992 673794 599004
rect 675386 598992 675392 599004
rect 673788 598964 675392 598992
rect 673788 598952 673794 598964
rect 675386 598952 675392 598964
rect 675444 598952 675450 599004
rect 42426 598884 42432 598936
rect 42484 598924 42490 598936
rect 62758 598924 62764 598936
rect 42484 598896 62764 598924
rect 42484 598884 42490 598896
rect 62758 598884 62764 598896
rect 62816 598884 62822 598936
rect 673454 598408 673460 598460
rect 673512 598448 673518 598460
rect 675478 598448 675484 598460
rect 673512 598420 675484 598448
rect 673512 598408 673518 598420
rect 675478 598408 675484 598420
rect 675536 598408 675542 598460
rect 673822 597116 673828 597168
rect 673880 597156 673886 597168
rect 675386 597156 675392 597168
rect 673880 597128 675392 597156
rect 673880 597116 673886 597128
rect 675386 597116 675392 597128
rect 675444 597116 675450 597168
rect 674650 596844 674656 596896
rect 674708 596884 674714 596896
rect 675386 596884 675392 596896
rect 674708 596856 675392 596884
rect 674708 596844 674714 596856
rect 675386 596844 675392 596856
rect 675444 596844 675450 596896
rect 674466 596572 674472 596624
rect 674524 596612 674530 596624
rect 674742 596612 674748 596624
rect 674524 596584 674748 596612
rect 674524 596572 674530 596584
rect 674742 596572 674748 596584
rect 674800 596572 674806 596624
rect 53742 596164 53748 596216
rect 53800 596204 53806 596216
rect 59170 596204 59176 596216
rect 53800 596176 59176 596204
rect 53800 596164 53806 596176
rect 59170 596164 59176 596176
rect 59228 596164 59234 596216
rect 674466 595280 674472 595332
rect 674524 595320 674530 595332
rect 675386 595320 675392 595332
rect 674524 595292 675392 595320
rect 674524 595280 674530 595292
rect 675386 595280 675392 595292
rect 675444 595280 675450 595332
rect 674374 593648 674380 593700
rect 674432 593688 674438 593700
rect 675478 593688 675484 593700
rect 674432 593660 675484 593688
rect 674432 593648 674438 593660
rect 675478 593648 675484 593660
rect 675536 593648 675542 593700
rect 656802 590656 656808 590708
rect 656860 590696 656866 590708
rect 669130 590696 669136 590708
rect 656860 590668 669136 590696
rect 656860 590656 656866 590668
rect 669130 590656 669136 590668
rect 669188 590656 669194 590708
rect 41506 589976 41512 590028
rect 41564 590016 41570 590028
rect 48866 590016 48872 590028
rect 41564 589988 48872 590016
rect 41564 589976 41570 589988
rect 48866 589976 48872 589988
rect 48924 589976 48930 590028
rect 673362 587868 673368 587920
rect 673420 587908 673426 587920
rect 678974 587908 678980 587920
rect 673420 587880 678980 587908
rect 673420 587868 673426 587880
rect 678974 587868 678980 587880
rect 679032 587868 679038 587920
rect 43346 586712 43352 586764
rect 43404 586752 43410 586764
rect 44082 586752 44088 586764
rect 43404 586724 44088 586752
rect 43404 586712 43410 586724
rect 44082 586712 44088 586724
rect 44140 586712 44146 586764
rect 42794 586576 42800 586628
rect 42852 586616 42858 586628
rect 43346 586616 43352 586628
rect 42852 586588 43352 586616
rect 42852 586576 42858 586588
rect 43346 586576 43352 586588
rect 43404 586576 43410 586628
rect 41138 585148 41144 585200
rect 41196 585188 41202 585200
rect 44174 585188 44180 585200
rect 41196 585160 44180 585188
rect 41196 585148 41202 585160
rect 44174 585148 44180 585160
rect 44232 585148 44238 585200
rect 44266 585148 44272 585200
rect 44324 585188 44330 585200
rect 48958 585188 48964 585200
rect 44324 585160 48964 585188
rect 44324 585148 44330 585160
rect 48958 585148 48964 585160
rect 49016 585148 49022 585200
rect 673362 584264 673368 584316
rect 673420 584304 673426 584316
rect 673546 584304 673552 584316
rect 673420 584276 673552 584304
rect 673420 584264 673426 584276
rect 673546 584264 673552 584276
rect 673604 584264 673610 584316
rect 41874 584196 41880 584248
rect 41932 584196 41938 584248
rect 41892 583976 41920 584196
rect 673546 584128 673552 584180
rect 673604 584168 673610 584180
rect 673914 584168 673920 584180
rect 673604 584140 673920 584168
rect 673604 584128 673610 584140
rect 673914 584128 673920 584140
rect 673972 584128 673978 584180
rect 674742 583992 674748 584044
rect 674800 584032 674806 584044
rect 675662 584032 675668 584044
rect 674800 584004 675668 584032
rect 674800 583992 674806 584004
rect 675662 583992 675668 584004
rect 675720 583992 675726 584044
rect 41874 583924 41880 583976
rect 41932 583924 41938 583976
rect 674466 583856 674472 583908
rect 674524 583896 674530 583908
rect 674742 583896 674748 583908
rect 674524 583868 674748 583896
rect 674524 583856 674530 583868
rect 674742 583856 674748 583868
rect 674800 583856 674806 583908
rect 42426 583720 42432 583772
rect 42484 583760 42490 583772
rect 42794 583760 42800 583772
rect 42484 583732 42800 583760
rect 42484 583720 42490 583732
rect 42794 583720 42800 583732
rect 42852 583720 42858 583772
rect 42886 583720 42892 583772
rect 42944 583760 42950 583772
rect 43070 583760 43076 583772
rect 42944 583732 43076 583760
rect 42944 583720 42950 583732
rect 43070 583720 43076 583732
rect 43128 583720 43134 583772
rect 673454 583720 673460 583772
rect 673512 583760 673518 583772
rect 673822 583760 673828 583772
rect 673512 583732 673828 583760
rect 673512 583720 673518 583732
rect 673822 583720 673828 583732
rect 673880 583720 673886 583772
rect 673914 583652 673920 583704
rect 673972 583692 673978 583704
rect 674374 583692 674380 583704
rect 673972 583664 674380 583692
rect 673972 583652 673978 583664
rect 674374 583652 674380 583664
rect 674432 583652 674438 583704
rect 43070 583584 43076 583636
rect 43128 583624 43134 583636
rect 43254 583624 43260 583636
rect 43128 583596 43260 583624
rect 43128 583584 43134 583596
rect 43254 583584 43260 583596
rect 43312 583584 43318 583636
rect 43254 583448 43260 583500
rect 43312 583488 43318 583500
rect 43990 583488 43996 583500
rect 43312 583460 43996 583488
rect 43312 583448 43318 583460
rect 43990 583448 43996 583460
rect 44048 583448 44054 583500
rect 44082 583448 44088 583500
rect 44140 583448 44146 583500
rect 44100 583160 44128 583448
rect 44082 583108 44088 583160
rect 44140 583108 44146 583160
rect 48958 582360 48964 582412
rect 49016 582400 49022 582412
rect 58434 582400 58440 582412
rect 49016 582372 58440 582400
rect 49016 582360 49022 582372
rect 58434 582360 58440 582372
rect 58492 582360 58498 582412
rect 42150 582088 42156 582140
rect 42208 582128 42214 582140
rect 42702 582128 42708 582140
rect 42208 582100 42708 582128
rect 42208 582088 42214 582100
rect 42702 582088 42708 582100
rect 42760 582088 42766 582140
rect 42150 581272 42156 581324
rect 42208 581312 42214 581324
rect 44266 581312 44272 581324
rect 42208 581284 44272 581312
rect 42208 581272 42214 581284
rect 44266 581272 44272 581284
rect 44324 581272 44330 581324
rect 42150 580252 42156 580304
rect 42208 580292 42214 580304
rect 43346 580292 43352 580304
rect 42208 580264 43352 580292
rect 42208 580252 42214 580264
rect 43346 580252 43352 580264
rect 43404 580252 43410 580304
rect 670602 580184 670608 580236
rect 670660 580224 670666 580236
rect 676030 580224 676036 580236
rect 670660 580196 676036 580224
rect 670660 580184 670666 580196
rect 676030 580184 676036 580196
rect 676088 580184 676094 580236
rect 666922 580048 666928 580100
rect 666980 580088 666986 580100
rect 676122 580088 676128 580100
rect 666980 580060 676128 580088
rect 666980 580048 666986 580060
rect 676122 580048 676128 580060
rect 676180 580048 676186 580100
rect 663794 579912 663800 579964
rect 663852 579952 663858 579964
rect 676214 579952 676220 579964
rect 663852 579924 676220 579952
rect 663852 579912 663858 579924
rect 676214 579912 676220 579924
rect 676272 579912 676278 579964
rect 663702 579776 663708 579828
rect 663760 579816 663766 579828
rect 676306 579816 676312 579828
rect 663760 579788 676312 579816
rect 663760 579776 663766 579788
rect 676306 579776 676312 579788
rect 676364 579776 676370 579828
rect 672534 579232 672540 579284
rect 672592 579272 672598 579284
rect 673270 579272 673276 579284
rect 672592 579244 673276 579272
rect 672592 579232 672598 579244
rect 673270 579232 673276 579244
rect 673328 579272 673334 579284
rect 676214 579272 676220 579284
rect 673328 579244 676220 579272
rect 673328 579232 673334 579244
rect 676214 579232 676220 579244
rect 676272 579232 676278 579284
rect 42150 578960 42156 579012
rect 42208 579000 42214 579012
rect 43530 579000 43536 579012
rect 42208 578972 43536 579000
rect 42208 578960 42214 578972
rect 43530 578960 43536 578972
rect 43588 578960 43594 579012
rect 42150 578416 42156 578468
rect 42208 578456 42214 578468
rect 43714 578456 43720 578468
rect 42208 578428 43720 578456
rect 42208 578416 42214 578428
rect 43714 578416 43720 578428
rect 43772 578416 43778 578468
rect 673086 578416 673092 578468
rect 673144 578456 673150 578468
rect 676214 578456 676220 578468
rect 673144 578428 676220 578456
rect 673144 578416 673150 578428
rect 676214 578416 676220 578428
rect 676272 578416 676278 578468
rect 42150 577804 42156 577856
rect 42208 577844 42214 577856
rect 43622 577844 43628 577856
rect 42208 577816 43628 577844
rect 42208 577804 42214 577816
rect 43622 577804 43628 577816
rect 43680 577804 43686 577856
rect 43622 577668 43628 577720
rect 43680 577708 43686 577720
rect 43990 577708 43996 577720
rect 43680 577680 43996 577708
rect 43680 577668 43686 577680
rect 43990 577668 43996 577680
rect 44048 577668 44054 577720
rect 672626 577600 672632 577652
rect 672684 577640 672690 577652
rect 673178 577640 673184 577652
rect 672684 577612 673184 577640
rect 672684 577600 672690 577612
rect 673178 577600 673184 577612
rect 673236 577640 673242 577652
rect 676214 577640 676220 577652
rect 673236 577612 676220 577640
rect 673236 577600 673242 577612
rect 676214 577600 676220 577612
rect 676272 577600 676278 577652
rect 42150 576920 42156 576972
rect 42208 576960 42214 576972
rect 44082 576960 44088 576972
rect 42208 576932 44088 576960
rect 42208 576920 42214 576932
rect 44082 576920 44088 576932
rect 44140 576920 44146 576972
rect 670510 576920 670516 576972
rect 670568 576960 670574 576972
rect 676214 576960 676220 576972
rect 670568 576932 676220 576960
rect 670568 576920 670574 576932
rect 676214 576920 676220 576932
rect 676272 576920 676278 576972
rect 655054 576852 655060 576904
rect 655112 576892 655118 576904
rect 663702 576892 663708 576904
rect 655112 576864 663708 576892
rect 655112 576852 655118 576864
rect 663702 576852 663708 576864
rect 663760 576852 663766 576904
rect 673362 576852 673368 576904
rect 673420 576892 673426 576904
rect 676030 576892 676036 576904
rect 673420 576864 676036 576892
rect 673420 576852 673426 576864
rect 676030 576852 676036 576864
rect 676088 576852 676094 576904
rect 674190 576784 674196 576836
rect 674248 576824 674254 576836
rect 675938 576824 675944 576836
rect 674248 576796 675944 576824
rect 674248 576784 674254 576796
rect 675938 576784 675944 576796
rect 675996 576784 676002 576836
rect 674558 576716 674564 576768
rect 674616 576756 674622 576768
rect 676030 576756 676036 576768
rect 674616 576728 676036 576756
rect 674616 576716 674622 576728
rect 676030 576716 676036 576728
rect 676088 576716 676094 576768
rect 673454 576648 673460 576700
rect 673512 576688 673518 576700
rect 676122 576688 676128 576700
rect 673512 576660 676128 576688
rect 673512 576648 673518 576660
rect 676122 576648 676128 576660
rect 676180 576648 676186 576700
rect 673546 576036 673552 576088
rect 673604 576076 673610 576088
rect 675938 576076 675944 576088
rect 673604 576048 675944 576076
rect 673604 576036 673610 576048
rect 675938 576036 675944 576048
rect 675996 576036 676002 576088
rect 42150 574676 42156 574728
rect 42208 574716 42214 574728
rect 43898 574716 43904 574728
rect 42208 574688 43904 574716
rect 42208 574676 42214 574688
rect 43898 574676 43904 574688
rect 43956 574676 43962 574728
rect 42150 573792 42156 573844
rect 42208 573832 42214 573844
rect 43162 573832 43168 573844
rect 42208 573804 43168 573832
rect 42208 573792 42214 573804
rect 43162 573792 43168 573804
rect 43220 573792 43226 573844
rect 674006 573588 674012 573640
rect 674064 573628 674070 573640
rect 676030 573628 676036 573640
rect 674064 573600 676036 573628
rect 674064 573588 674070 573600
rect 676030 573588 676036 573600
rect 676088 573588 676094 573640
rect 42150 573452 42156 573504
rect 42208 573492 42214 573504
rect 43622 573492 43628 573504
rect 42208 573464 43628 573492
rect 42208 573452 42214 573464
rect 43622 573452 43628 573464
rect 43680 573452 43686 573504
rect 673638 572772 673644 572824
rect 673696 572812 673702 572824
rect 676030 572812 676036 572824
rect 673696 572784 676036 572812
rect 673696 572772 673702 572784
rect 676030 572772 676036 572784
rect 676088 572772 676094 572824
rect 42058 572636 42064 572688
rect 42116 572676 42122 572688
rect 43806 572676 43812 572688
rect 42116 572648 43812 572676
rect 42116 572636 42122 572648
rect 43806 572636 43812 572648
rect 43864 572636 43870 572688
rect 42058 570868 42064 570920
rect 42116 570908 42122 570920
rect 43070 570908 43076 570920
rect 42116 570880 43076 570908
rect 42116 570868 42122 570880
rect 43070 570868 43076 570880
rect 43128 570868 43134 570920
rect 42150 570256 42156 570308
rect 42208 570296 42214 570308
rect 42978 570296 42984 570308
rect 42208 570268 42984 570296
rect 42208 570256 42214 570268
rect 42978 570256 42984 570268
rect 43036 570256 43042 570308
rect 42058 569576 42064 569628
rect 42116 569616 42122 569628
rect 42886 569616 42892 569628
rect 42116 569588 42892 569616
rect 42116 569576 42122 569588
rect 42886 569576 42892 569588
rect 42944 569576 42950 569628
rect 672534 568556 672540 568608
rect 672592 568596 672598 568608
rect 678974 568596 678980 568608
rect 672592 568568 678980 568596
rect 672592 568556 672598 568568
rect 678974 568556 678980 568568
rect 679032 568556 679038 568608
rect 673546 559512 673552 559564
rect 673604 559552 673610 559564
rect 675478 559552 675484 559564
rect 673604 559524 675484 559552
rect 673604 559512 673610 559524
rect 675478 559512 675484 559524
rect 675536 559512 675542 559564
rect 41506 558764 41512 558816
rect 41564 558804 41570 558816
rect 48958 558804 48964 558816
rect 41564 558776 48964 558804
rect 41564 558764 41570 558776
rect 48958 558764 48964 558776
rect 49016 558764 49022 558816
rect 41414 558492 41420 558544
rect 41472 558532 41478 558544
rect 53742 558532 53748 558544
rect 41472 558504 53748 558532
rect 41472 558492 41478 558504
rect 53742 558492 53748 558504
rect 53800 558492 53806 558544
rect 41506 558424 41512 558476
rect 41564 558464 41570 558476
rect 58434 558464 58440 558476
rect 41564 558436 58440 558464
rect 41564 558424 41570 558436
rect 58434 558424 58440 558436
rect 58492 558424 58498 558476
rect 49050 557540 49056 557592
rect 49108 557580 49114 557592
rect 58342 557580 58348 557592
rect 49108 557552 58348 557580
rect 49108 557540 49114 557552
rect 58342 557540 58348 557552
rect 58400 557540 58406 557592
rect 654318 556112 654324 556164
rect 654376 556152 654382 556164
rect 675294 556152 675300 556164
rect 654376 556124 675300 556152
rect 654376 556112 654382 556124
rect 675294 556112 675300 556124
rect 675352 556112 675358 556164
rect 673914 555228 673920 555280
rect 673972 555268 673978 555280
rect 675386 555268 675392 555280
rect 673972 555240 675392 555268
rect 673972 555228 673978 555240
rect 675386 555228 675392 555240
rect 675444 555228 675450 555280
rect 673454 554548 673460 554600
rect 673512 554588 673518 554600
rect 675386 554588 675392 554600
rect 673512 554560 675392 554588
rect 673512 554548 673518 554560
rect 675386 554548 675392 554560
rect 675444 554548 675450 554600
rect 674006 553732 674012 553784
rect 674064 553772 674070 553784
rect 675386 553772 675392 553784
rect 674064 553744 675392 553772
rect 674064 553732 674070 553744
rect 675386 553732 675392 553744
rect 675444 553732 675450 553784
rect 673638 553188 673644 553240
rect 673696 553228 673702 553240
rect 675386 553228 675392 553240
rect 673696 553200 675392 553228
rect 673696 553188 673702 553200
rect 675386 553188 675392 553200
rect 675444 553188 675450 553240
rect 674190 551896 674196 551948
rect 674248 551936 674254 551948
rect 675386 551936 675392 551948
rect 674248 551908 675392 551936
rect 674248 551896 674254 551908
rect 675386 551896 675392 551908
rect 675444 551896 675450 551948
rect 654686 549244 654692 549296
rect 654744 549284 654750 549296
rect 663794 549284 663800 549296
rect 654744 549256 663800 549284
rect 654744 549244 654750 549256
rect 663794 549244 663800 549256
rect 663852 549244 663858 549296
rect 41506 548632 41512 548684
rect 41564 548672 41570 548684
rect 43530 548672 43536 548684
rect 41564 548644 43536 548672
rect 41564 548632 41570 548644
rect 43530 548632 43536 548644
rect 43588 548632 43594 548684
rect 674558 548292 674564 548344
rect 674616 548332 674622 548344
rect 675386 548332 675392 548344
rect 674616 548304 675392 548332
rect 674616 548292 674622 548304
rect 675386 548292 675392 548304
rect 675444 548292 675450 548344
rect 674650 548224 674656 548276
rect 674708 548264 674714 548276
rect 675294 548264 675300 548276
rect 674708 548236 675300 548264
rect 674708 548224 674714 548236
rect 675294 548224 675300 548236
rect 675352 548224 675358 548276
rect 41598 546864 41604 546916
rect 41656 546904 41662 546916
rect 48958 546904 48964 546916
rect 41656 546876 48964 546904
rect 41656 546864 41662 546876
rect 48958 546864 48964 546876
rect 49016 546864 49022 546916
rect 41506 546728 41512 546780
rect 41564 546768 41570 546780
rect 42794 546768 42800 546780
rect 41564 546740 42800 546768
rect 41564 546728 41570 546740
rect 42794 546728 42800 546740
rect 42852 546728 42858 546780
rect 673086 546252 673092 546304
rect 673144 546292 673150 546304
rect 679066 546292 679072 546304
rect 673144 546264 679072 546292
rect 673144 546252 673150 546264
rect 679066 546252 679072 546264
rect 679124 546252 679130 546304
rect 53834 543736 53840 543788
rect 53892 543776 53898 543788
rect 58342 543776 58348 543788
rect 53892 543748 58348 543776
rect 53892 543736 53898 543748
rect 58342 543736 58348 543748
rect 58400 543736 58406 543788
rect 43714 541696 43720 541748
rect 43772 541736 43778 541748
rect 50982 541736 50988 541748
rect 43772 541708 50988 541736
rect 43772 541696 43778 541708
rect 50982 541696 50988 541708
rect 51040 541696 51046 541748
rect 41782 541016 41788 541068
rect 41840 541016 41846 541068
rect 41800 540796 41828 541016
rect 41782 540744 41788 540796
rect 41840 540744 41846 540796
rect 42058 538908 42064 538960
rect 42116 538948 42122 538960
rect 42702 538948 42708 538960
rect 42116 538920 42708 538948
rect 42116 538908 42122 538920
rect 42702 538908 42708 538920
rect 42760 538908 42766 538960
rect 42150 538092 42156 538144
rect 42208 538132 42214 538144
rect 43714 538132 43720 538144
rect 42208 538104 43720 538132
rect 42208 538092 42214 538104
rect 43714 538092 43720 538104
rect 43772 538092 43778 538144
rect 42058 537072 42064 537124
rect 42116 537112 42122 537124
rect 42978 537112 42984 537124
rect 42116 537084 42984 537112
rect 42116 537072 42122 537084
rect 42978 537072 42984 537084
rect 43036 537072 43042 537124
rect 42978 536936 42984 536988
rect 43036 536976 43042 536988
rect 43162 536976 43168 536988
rect 43036 536948 43168 536976
rect 43036 536936 43042 536948
rect 43162 536936 43168 536948
rect 43220 536936 43226 536988
rect 43162 536800 43168 536852
rect 43220 536840 43226 536852
rect 43346 536840 43352 536852
rect 43220 536812 43352 536840
rect 43220 536800 43226 536812
rect 43346 536800 43352 536812
rect 43404 536800 43410 536852
rect 43346 536664 43352 536716
rect 43404 536704 43410 536716
rect 43622 536704 43628 536716
rect 43404 536676 43628 536704
rect 43404 536664 43410 536676
rect 43622 536664 43628 536676
rect 43680 536664 43686 536716
rect 654870 536392 654876 536444
rect 654928 536432 654934 536444
rect 666462 536432 666468 536444
rect 654928 536404 666468 536432
rect 654928 536392 654934 536404
rect 666462 536392 666468 536404
rect 666520 536392 666526 536444
rect 42150 535780 42156 535832
rect 42208 535820 42214 535832
rect 42794 535820 42800 535832
rect 42208 535792 42800 535820
rect 42208 535780 42214 535792
rect 42794 535780 42800 535792
rect 42852 535780 42858 535832
rect 663886 535712 663892 535764
rect 663944 535752 663950 535764
rect 676214 535752 676220 535764
rect 663944 535724 676220 535752
rect 663944 535712 663950 535724
rect 676214 535712 676220 535724
rect 676272 535712 676278 535764
rect 660942 535576 660948 535628
rect 661000 535616 661006 535628
rect 676030 535616 676036 535628
rect 661000 535588 676036 535616
rect 661000 535576 661006 535588
rect 676030 535576 676036 535588
rect 676088 535576 676094 535628
rect 42058 535032 42064 535084
rect 42116 535072 42122 535084
rect 43254 535072 43260 535084
rect 42116 535044 43260 535072
rect 42116 535032 42122 535044
rect 43254 535032 43260 535044
rect 43312 535032 43318 535084
rect 673270 534896 673276 534948
rect 673328 534936 673334 534948
rect 676030 534936 676036 534948
rect 673328 534908 676036 534936
rect 673328 534896 673334 534908
rect 676030 534896 676036 534908
rect 676088 534896 676094 534948
rect 42150 534420 42156 534472
rect 42208 534460 42214 534472
rect 43530 534460 43536 534472
rect 42208 534432 43536 534460
rect 42208 534420 42214 534432
rect 43530 534420 43536 534432
rect 43588 534420 43594 534472
rect 42150 533944 42156 533996
rect 42208 533984 42214 533996
rect 43346 533984 43352 533996
rect 42208 533956 43352 533984
rect 42208 533944 42214 533956
rect 43346 533944 43352 533956
rect 43404 533944 43410 533996
rect 673178 533264 673184 533316
rect 673236 533304 673242 533316
rect 676030 533304 676036 533316
rect 673236 533276 676036 533304
rect 673236 533264 673242 533276
rect 676030 533264 676036 533276
rect 676088 533264 676094 533316
rect 669038 532856 669044 532908
rect 669096 532896 669102 532908
rect 678974 532896 678980 532908
rect 669096 532868 678980 532896
rect 669096 532856 669102 532868
rect 678974 532856 678980 532868
rect 679032 532856 679038 532908
rect 670050 532788 670056 532840
rect 670108 532828 670114 532840
rect 675846 532828 675852 532840
rect 670108 532800 675852 532828
rect 670108 532788 670114 532800
rect 675846 532788 675852 532800
rect 675904 532828 675910 532840
rect 676122 532828 676128 532840
rect 675904 532800 676128 532828
rect 675904 532788 675910 532800
rect 676122 532788 676128 532800
rect 676180 532788 676186 532840
rect 674742 532652 674748 532704
rect 674800 532692 674806 532704
rect 676030 532692 676036 532704
rect 674800 532664 676036 532692
rect 674800 532652 674806 532664
rect 676030 532652 676036 532664
rect 676088 532652 676094 532704
rect 672810 532584 672816 532636
rect 672868 532624 672874 532636
rect 673362 532624 673368 532636
rect 672868 532596 673368 532624
rect 672868 532584 672874 532596
rect 673362 532584 673368 532596
rect 673420 532624 673426 532636
rect 676214 532624 676220 532636
rect 673420 532596 676220 532624
rect 673420 532584 673426 532596
rect 676214 532584 676220 532596
rect 676272 532584 676278 532636
rect 42150 531428 42156 531480
rect 42208 531468 42214 531480
rect 43898 531468 43904 531480
rect 42208 531440 43904 531468
rect 42208 531428 42214 531440
rect 43898 531428 43904 531440
rect 43956 531428 43962 531480
rect 674282 531088 674288 531140
rect 674340 531128 674346 531140
rect 676030 531128 676036 531140
rect 674340 531100 676036 531128
rect 674340 531088 674346 531100
rect 676030 531088 676036 531100
rect 676088 531088 676094 531140
rect 42150 530680 42156 530732
rect 42208 530720 42214 530732
rect 43990 530720 43996 530732
rect 42208 530692 43996 530720
rect 42208 530680 42214 530692
rect 43990 530680 43996 530692
rect 44048 530680 44054 530732
rect 42150 530272 42156 530324
rect 42208 530312 42214 530324
rect 43070 530312 43076 530324
rect 42208 530284 43076 530312
rect 42208 530272 42214 530284
rect 43070 530272 43076 530284
rect 43128 530272 43134 530324
rect 674466 529864 674472 529916
rect 674524 529904 674530 529916
rect 676030 529904 676036 529916
rect 674524 529876 676036 529904
rect 674524 529864 674530 529876
rect 676030 529864 676036 529876
rect 676088 529864 676094 529916
rect 42150 529456 42156 529508
rect 42208 529496 42214 529508
rect 43162 529496 43168 529508
rect 42208 529468 43168 529496
rect 42208 529456 42214 529468
rect 43162 529456 43168 529468
rect 43220 529456 43226 529508
rect 674374 529456 674380 529508
rect 674432 529496 674438 529508
rect 676030 529496 676036 529508
rect 674432 529468 676036 529496
rect 674432 529456 674438 529468
rect 676030 529456 676036 529468
rect 676088 529456 676094 529508
rect 673730 527824 673736 527876
rect 673788 527864 673794 527876
rect 676030 527864 676036 527876
rect 673788 527836 676036 527864
rect 673788 527824 673794 527836
rect 676030 527824 676036 527836
rect 676088 527824 676094 527876
rect 42150 527212 42156 527264
rect 42208 527252 42214 527264
rect 43438 527252 43444 527264
rect 42208 527224 43444 527252
rect 42208 527212 42214 527224
rect 43438 527212 43444 527224
rect 43496 527212 43502 527264
rect 42058 527144 42064 527196
rect 42116 527184 42122 527196
rect 43806 527184 43812 527196
rect 42116 527156 43812 527184
rect 42116 527144 42122 527156
rect 43806 527144 43812 527156
rect 43864 527144 43870 527196
rect 673822 527076 673828 527128
rect 673880 527116 673886 527128
rect 676030 527116 676036 527128
rect 673880 527088 676036 527116
rect 673880 527076 673886 527088
rect 676030 527076 676036 527088
rect 676088 527076 676094 527128
rect 42150 526600 42156 526652
rect 42208 526640 42214 526652
rect 42978 526640 42984 526652
rect 42208 526612 42984 526640
rect 42208 526600 42214 526612
rect 42978 526600 42984 526612
rect 43036 526600 43042 526652
rect 672626 524424 672632 524476
rect 672684 524464 672690 524476
rect 678974 524464 678980 524476
rect 672684 524436 678980 524464
rect 672684 524424 672690 524436
rect 678974 524424 678980 524436
rect 679032 524424 679038 524476
rect 677492 524356 677498 524408
rect 677550 524396 677556 524408
rect 679066 524396 679072 524408
rect 677550 524368 679072 524396
rect 677550 524356 677556 524368
rect 679066 524356 679072 524368
rect 679124 524356 679130 524408
rect 675846 523948 675852 524000
rect 675904 523988 675910 524000
rect 676122 523988 676128 524000
rect 675904 523960 676128 523988
rect 675904 523948 675910 523960
rect 676122 523948 676128 523960
rect 676180 523948 676186 524000
rect 654134 522452 654140 522504
rect 654192 522492 654198 522504
rect 661218 522492 661224 522504
rect 654192 522464 661224 522492
rect 654192 522452 654198 522464
rect 661218 522452 661224 522464
rect 661276 522452 661282 522504
rect 51258 518916 51264 518968
rect 51316 518956 51322 518968
rect 58434 518956 58440 518968
rect 51316 518928 58440 518956
rect 51316 518916 51322 518928
rect 58434 518916 58440 518928
rect 58492 518916 58498 518968
rect 654870 510824 654876 510876
rect 654928 510864 654934 510876
rect 670510 510864 670516 510876
rect 654928 510836 670516 510864
rect 654928 510824 654934 510836
rect 670510 510824 670516 510836
rect 670568 510824 670574 510876
rect 50982 505112 50988 505164
rect 51040 505152 51046 505164
rect 58434 505152 58440 505164
rect 51040 505124 58440 505152
rect 51040 505112 51046 505124
rect 58434 505112 58440 505124
rect 58492 505112 58498 505164
rect 656802 497632 656808 497684
rect 656860 497672 656866 497684
rect 663886 497672 663892 497684
rect 656860 497644 663892 497672
rect 656860 497632 656866 497644
rect 663886 497632 663892 497644
rect 663944 497632 663950 497684
rect 675570 492192 675576 492244
rect 675628 492232 675634 492244
rect 676030 492232 676036 492244
rect 675628 492204 676036 492232
rect 675628 492192 675634 492204
rect 676030 492192 676036 492204
rect 676088 492192 676094 492244
rect 669130 491648 669136 491700
rect 669188 491688 669194 491700
rect 676030 491688 676036 491700
rect 669188 491660 676036 491688
rect 669188 491648 669194 491660
rect 676030 491648 676036 491660
rect 676088 491648 676094 491700
rect 663702 491512 663708 491564
rect 663760 491552 663766 491564
rect 676030 491552 676036 491564
rect 663760 491524 676036 491552
rect 663760 491512 663766 491524
rect 676030 491512 676036 491524
rect 676088 491512 676094 491564
rect 661034 491376 661040 491428
rect 661092 491416 661098 491428
rect 675938 491416 675944 491428
rect 661092 491388 675944 491416
rect 661092 491376 661098 491388
rect 675938 491376 675944 491388
rect 675996 491376 676002 491428
rect 49142 491308 49148 491360
rect 49200 491348 49206 491360
rect 57974 491348 57980 491360
rect 49200 491320 57980 491348
rect 49200 491308 49206 491320
rect 57974 491308 57980 491320
rect 58032 491308 58038 491360
rect 676214 491240 676220 491292
rect 676272 491280 676278 491292
rect 677502 491280 677508 491292
rect 676272 491252 677508 491280
rect 676272 491240 676278 491252
rect 677502 491240 677508 491252
rect 677560 491240 677566 491292
rect 669682 488520 669688 488572
rect 669740 488560 669746 488572
rect 675662 488560 675668 488572
rect 669740 488532 675668 488560
rect 669740 488520 669746 488532
rect 675662 488520 675668 488532
rect 675720 488560 675726 488572
rect 675938 488560 675944 488572
rect 675720 488532 675944 488560
rect 675720 488520 675726 488532
rect 675938 488520 675944 488532
rect 675996 488520 676002 488572
rect 674650 488180 674656 488232
rect 674708 488220 674714 488232
rect 676030 488220 676036 488232
rect 674708 488192 676036 488220
rect 674708 488180 674714 488192
rect 676030 488180 676036 488192
rect 676088 488180 676094 488232
rect 673546 487908 673552 487960
rect 673604 487948 673610 487960
rect 675662 487948 675668 487960
rect 673604 487920 675668 487948
rect 673604 487908 673610 487920
rect 675662 487908 675668 487920
rect 675720 487908 675726 487960
rect 673914 487092 673920 487144
rect 673972 487132 673978 487144
rect 676030 487132 676036 487144
rect 673972 487104 676036 487132
rect 673972 487092 673978 487104
rect 676030 487092 676036 487104
rect 676088 487092 676094 487144
rect 669682 485800 669688 485852
rect 669740 485840 669746 485852
rect 675570 485840 675576 485852
rect 669740 485812 675576 485840
rect 669740 485800 669746 485812
rect 675570 485800 675576 485812
rect 675628 485800 675634 485852
rect 674558 485732 674564 485784
rect 674616 485772 674622 485784
rect 676030 485772 676036 485784
rect 674616 485744 676036 485772
rect 674616 485732 674622 485744
rect 676030 485732 676036 485744
rect 676088 485732 676094 485784
rect 674190 485460 674196 485512
rect 674248 485500 674254 485512
rect 676030 485500 676036 485512
rect 674248 485472 676036 485500
rect 674248 485460 674254 485472
rect 676030 485460 676036 485472
rect 676088 485460 676094 485512
rect 654870 483012 654876 483064
rect 654928 483052 654934 483064
rect 669130 483052 669136 483064
rect 654928 483024 669136 483052
rect 654928 483012 654934 483024
rect 669130 483012 669136 483024
rect 669188 483012 669194 483064
rect 673638 482944 673644 482996
rect 673696 482984 673702 482996
rect 676030 482984 676036 482996
rect 673696 482956 676036 482984
rect 673696 482944 673702 482956
rect 676030 482944 676036 482956
rect 676088 482944 676094 482996
rect 673454 482876 673460 482928
rect 673512 482916 673518 482928
rect 675662 482916 675668 482928
rect 673512 482888 675668 482916
rect 673512 482876 673518 482888
rect 675662 482876 675668 482888
rect 675720 482876 675726 482928
rect 672718 480700 672724 480752
rect 672776 480740 672782 480752
rect 676030 480740 676036 480752
rect 672776 480712 676036 480740
rect 672776 480700 672782 480712
rect 676030 480700 676036 480712
rect 676088 480700 676094 480752
rect 51166 480224 51172 480276
rect 51224 480264 51230 480276
rect 58434 480264 58440 480276
rect 51224 480236 58440 480264
rect 51224 480224 51230 480236
rect 58434 480224 58440 480236
rect 58492 480224 58498 480276
rect 675938 478592 675944 478644
rect 675996 478592 676002 478644
rect 675956 478428 675984 478592
rect 676030 478428 676036 478440
rect 675956 478400 676036 478428
rect 676030 478388 676036 478400
rect 676088 478388 676094 478440
rect 654870 470772 654876 470824
rect 654928 470812 654934 470824
rect 660942 470812 660948 470824
rect 654928 470784 660948 470812
rect 654928 470772 654934 470784
rect 660942 470772 660948 470784
rect 661000 470772 661006 470824
rect 54018 466420 54024 466472
rect 54076 466460 54082 466472
rect 58710 466460 58716 466472
rect 54076 466432 58716 466460
rect 54076 466420 54082 466432
rect 58710 466420 58716 466432
rect 58768 466420 58774 466472
rect 654226 457444 654232 457496
rect 654284 457484 654290 457496
rect 667014 457484 667020 457496
rect 654284 457456 667020 457484
rect 654284 457444 654290 457456
rect 667014 457444 667020 457456
rect 667072 457444 667078 457496
rect 53742 452616 53748 452668
rect 53800 452656 53806 452668
rect 59170 452656 59176 452668
rect 53800 452628 59176 452656
rect 53800 452616 53806 452628
rect 59170 452616 59176 452628
rect 59228 452616 59234 452668
rect 654410 444456 654416 444508
rect 654468 444496 654474 444508
rect 663978 444496 663984 444508
rect 654468 444468 663984 444496
rect 654468 444456 654474 444468
rect 663978 444456 663984 444468
rect 664036 444456 664042 444508
rect 51074 438880 51080 438932
rect 51132 438920 51138 438932
rect 58434 438920 58440 438932
rect 51132 438892 58440 438920
rect 51132 438880 51138 438892
rect 58434 438880 58440 438892
rect 58492 438880 58498 438932
rect 41782 430788 41788 430840
rect 41840 430828 41846 430840
rect 59262 430828 59268 430840
rect 41840 430800 59268 430828
rect 41840 430788 41846 430800
rect 59262 430788 59268 430800
rect 59320 430788 59326 430840
rect 654686 430584 654692 430636
rect 654744 430624 654750 430636
rect 663702 430624 663708 430636
rect 654744 430596 663708 430624
rect 654744 430584 654750 430596
rect 663702 430584 663708 430596
rect 663760 430584 663766 430636
rect 53926 427864 53932 427916
rect 53984 427904 53990 427916
rect 58250 427904 58256 427916
rect 53984 427876 58256 427904
rect 53984 427864 53990 427876
rect 58250 427864 58256 427876
rect 58308 427864 58314 427916
rect 41782 427796 41788 427848
rect 41840 427836 41846 427848
rect 44082 427836 44088 427848
rect 41840 427808 44088 427836
rect 41840 427796 41846 427808
rect 44082 427796 44088 427808
rect 44140 427836 44146 427848
rect 62758 427836 62764 427848
rect 44140 427808 62764 427836
rect 44140 427796 44146 427808
rect 62758 427796 62764 427808
rect 62816 427796 62822 427848
rect 41782 419432 41788 419484
rect 41840 419472 41846 419484
rect 46658 419472 46664 419484
rect 41840 419444 46664 419472
rect 41840 419432 41846 419444
rect 46658 419432 46664 419444
rect 46716 419432 46722 419484
rect 655054 416780 655060 416832
rect 655112 416820 655118 416832
rect 661034 416820 661040 416832
rect 655112 416792 661040 416820
rect 655112 416780 655118 416792
rect 661034 416780 661040 416792
rect 661092 416780 661098 416832
rect 41874 416304 41880 416356
rect 41932 416344 41938 416356
rect 43070 416344 43076 416356
rect 41932 416316 43076 416344
rect 41932 416304 41938 416316
rect 43070 416304 43076 416316
rect 43128 416304 43134 416356
rect 49234 413992 49240 414044
rect 49292 414032 49298 414044
rect 58434 414032 58440 414044
rect 49292 414004 58440 414032
rect 49292 413992 49298 414004
rect 58434 413992 58440 414004
rect 58492 413992 58498 414044
rect 42150 413108 42156 413160
rect 42208 413148 42214 413160
rect 42334 413148 42340 413160
rect 42208 413120 42340 413148
rect 42208 413108 42214 413120
rect 42334 413108 42340 413120
rect 42392 413108 42398 413160
rect 42794 411340 42800 411392
rect 42852 411340 42858 411392
rect 42150 411272 42156 411324
rect 42208 411312 42214 411324
rect 42812 411312 42840 411340
rect 42208 411284 42840 411312
rect 42208 411272 42214 411284
rect 675754 411068 675760 411120
rect 675812 411108 675818 411120
rect 676122 411108 676128 411120
rect 675812 411080 676128 411108
rect 675812 411068 675818 411080
rect 676122 411068 676128 411080
rect 676180 411068 676186 411120
rect 42150 410660 42156 410712
rect 42208 410700 42214 410712
rect 49050 410700 49056 410712
rect 42208 410672 49056 410700
rect 42208 410660 42214 410672
rect 49050 410660 49056 410672
rect 49108 410660 49114 410712
rect 42150 409436 42156 409488
rect 42208 409476 42214 409488
rect 42978 409476 42984 409488
rect 42208 409448 42984 409476
rect 42208 409436 42214 409448
rect 42978 409436 42984 409448
rect 43036 409436 43042 409488
rect 42058 408144 42064 408196
rect 42116 408184 42122 408196
rect 42518 408184 42524 408196
rect 42116 408156 42524 408184
rect 42116 408144 42122 408156
rect 42518 408144 42524 408156
rect 42576 408144 42582 408196
rect 42150 407464 42156 407516
rect 42208 407504 42214 407516
rect 43162 407504 43168 407516
rect 42208 407476 43168 407504
rect 42208 407464 42214 407476
rect 43162 407464 43168 407476
rect 43220 407464 43226 407516
rect 42058 406988 42064 407040
rect 42116 407028 42122 407040
rect 43070 407028 43076 407040
rect 42116 407000 43076 407028
rect 42116 406988 42122 407000
rect 43070 406988 43076 407000
rect 43128 406988 43134 407040
rect 42150 406172 42156 406224
rect 42208 406212 42214 406224
rect 43438 406212 43444 406224
rect 42208 406184 43444 406212
rect 42208 406172 42214 406184
rect 43438 406172 43444 406184
rect 43496 406172 43502 406224
rect 654870 403996 654876 404048
rect 654928 404036 654934 404048
rect 661126 404036 661132 404048
rect 654928 404008 661132 404036
rect 654928 403996 654934 404008
rect 661126 403996 661132 404008
rect 661184 403996 661190 404048
rect 42150 403860 42156 403912
rect 42208 403900 42214 403912
rect 43990 403900 43996 403912
rect 42208 403872 43996 403900
rect 42208 403860 42214 403872
rect 43990 403860 43996 403872
rect 44048 403860 44054 403912
rect 666462 403384 666468 403436
rect 666520 403424 666526 403436
rect 676214 403424 676220 403436
rect 666520 403396 676220 403424
rect 666520 403384 666526 403396
rect 676214 403384 676220 403396
rect 676272 403384 676278 403436
rect 42150 403316 42156 403368
rect 42208 403356 42214 403368
rect 43530 403356 43536 403368
rect 42208 403328 43536 403356
rect 42208 403316 42214 403328
rect 43530 403316 43536 403328
rect 43588 403316 43594 403368
rect 663794 403248 663800 403300
rect 663852 403288 663858 403300
rect 676214 403288 676220 403300
rect 663852 403260 676220 403288
rect 663852 403248 663858 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 661218 403112 661224 403164
rect 661276 403152 661282 403164
rect 675938 403152 675944 403164
rect 661276 403124 675944 403152
rect 661276 403112 661282 403124
rect 675938 403112 675944 403124
rect 675996 403112 676002 403164
rect 42150 402500 42156 402552
rect 42208 402540 42214 402552
rect 43714 402540 43720 402552
rect 42208 402512 43720 402540
rect 42208 402500 42214 402512
rect 43714 402500 43720 402512
rect 43772 402500 43778 402552
rect 43806 402432 43812 402484
rect 43864 402432 43870 402484
rect 43824 402280 43852 402432
rect 43806 402228 43812 402280
rect 43864 402228 43870 402280
rect 42150 402024 42156 402076
rect 42208 402064 42214 402076
rect 43346 402064 43352 402076
rect 42208 402036 43352 402064
rect 42208 402024 42214 402036
rect 43346 402024 43352 402036
rect 43404 402024 43410 402076
rect 675110 400392 675116 400444
rect 675168 400432 675174 400444
rect 676122 400432 676128 400444
rect 675168 400404 676128 400432
rect 675168 400392 675174 400404
rect 676122 400392 676128 400404
rect 676180 400392 676186 400444
rect 49050 400188 49056 400240
rect 49108 400228 49114 400240
rect 58434 400228 58440 400240
rect 49108 400200 58440 400228
rect 49108 400188 49114 400200
rect 58434 400188 58440 400200
rect 58492 400188 58498 400240
rect 42150 399984 42156 400036
rect 42208 400024 42214 400036
rect 42886 400024 42892 400036
rect 42208 399996 42892 400024
rect 42208 399984 42214 399996
rect 42886 399984 42892 399996
rect 42944 399984 42950 400036
rect 42150 399440 42156 399492
rect 42208 399480 42214 399492
rect 43714 399480 43720 399492
rect 42208 399452 43720 399480
rect 42208 399440 42214 399452
rect 43714 399440 43720 399452
rect 43772 399440 43778 399492
rect 674374 399440 674380 399492
rect 674432 399480 674438 399492
rect 676030 399480 676036 399492
rect 674432 399452 676036 399480
rect 674432 399440 674438 399452
rect 676030 399440 676036 399452
rect 676088 399440 676094 399492
rect 42150 398760 42156 398812
rect 42208 398800 42214 398812
rect 43254 398800 43260 398812
rect 42208 398772 43260 398800
rect 42208 398760 42214 398772
rect 43254 398760 43260 398772
rect 43312 398760 43318 398812
rect 674466 398216 674472 398268
rect 674524 398256 674530 398268
rect 676030 398256 676036 398268
rect 674524 398228 676036 398256
rect 674524 398216 674530 398228
rect 676030 398216 676036 398228
rect 676088 398216 676094 398268
rect 673822 397604 673828 397656
rect 673880 397644 673886 397656
rect 675938 397644 675944 397656
rect 673880 397616 675944 397644
rect 673880 397604 673886 397616
rect 675938 397604 675944 397616
rect 675996 397604 676002 397656
rect 674282 397536 674288 397588
rect 674340 397576 674346 397588
rect 676122 397576 676128 397588
rect 674340 397548 676128 397576
rect 674340 397536 674346 397548
rect 676122 397536 676128 397548
rect 676180 397536 676186 397588
rect 674650 397468 674656 397520
rect 674708 397508 674714 397520
rect 676030 397508 676036 397520
rect 674708 397480 676036 397508
rect 674708 397468 674714 397480
rect 676030 397468 676036 397480
rect 676088 397468 676094 397520
rect 673454 396584 673460 396636
rect 673512 396624 673518 396636
rect 676030 396624 676036 396636
rect 673512 396596 676036 396624
rect 673512 396584 673518 396596
rect 676030 396584 676036 396596
rect 676088 396584 676094 396636
rect 673546 395360 673552 395412
rect 673604 395400 673610 395412
rect 675938 395400 675944 395412
rect 673604 395372 675944 395400
rect 673604 395360 673610 395372
rect 675938 395360 675944 395372
rect 675996 395360 676002 395412
rect 675018 394952 675024 395004
rect 675076 394992 675082 395004
rect 676030 394992 676036 395004
rect 675076 394964 676036 394992
rect 675076 394952 675082 394964
rect 676030 394952 676036 394964
rect 676088 394952 676094 395004
rect 673638 394816 673644 394868
rect 673696 394856 673702 394868
rect 675938 394856 675944 394868
rect 673696 394828 675944 394856
rect 673696 394816 673702 394828
rect 675938 394816 675944 394828
rect 675996 394816 676002 394868
rect 674926 394748 674932 394800
rect 674984 394788 674990 394800
rect 676122 394788 676128 394800
rect 674984 394760 676128 394788
rect 674984 394748 674990 394760
rect 676122 394748 676128 394760
rect 676180 394748 676186 394800
rect 675202 394680 675208 394732
rect 675260 394720 675266 394732
rect 676030 394720 676036 394732
rect 675260 394692 676036 394720
rect 675260 394680 675266 394692
rect 676030 394680 676036 394692
rect 676088 394680 676094 394732
rect 672902 392096 672908 392148
rect 672960 392136 672966 392148
rect 679066 392136 679072 392148
rect 672960 392108 679072 392136
rect 672960 392096 672966 392108
rect 679066 392096 679072 392108
rect 679124 392096 679130 392148
rect 673730 392028 673736 392080
rect 673788 392068 673794 392080
rect 676122 392068 676128 392080
rect 673788 392040 676128 392068
rect 673788 392028 673794 392040
rect 676122 392028 676128 392040
rect 676180 392028 676186 392080
rect 674006 391960 674012 392012
rect 674064 392000 674070 392012
rect 676030 392000 676036 392012
rect 674064 391972 676036 392000
rect 674064 391960 674070 391972
rect 676030 391960 676036 391972
rect 676088 391960 676094 392012
rect 674742 390532 674748 390584
rect 674800 390572 674806 390584
rect 675754 390572 675760 390584
rect 674800 390544 675760 390572
rect 674800 390532 674806 390544
rect 675754 390532 675760 390544
rect 675812 390532 675818 390584
rect 674558 390464 674564 390516
rect 674616 390504 674622 390516
rect 675662 390504 675668 390516
rect 674616 390476 675668 390504
rect 674616 390464 674622 390476
rect 675662 390464 675668 390476
rect 675720 390464 675726 390516
rect 654318 389852 654324 389904
rect 654376 389892 654382 389904
rect 666462 389892 666468 389904
rect 654376 389864 666468 389892
rect 654376 389852 654382 389864
rect 666462 389852 666468 389864
rect 666520 389852 666526 389904
rect 53834 389172 53840 389224
rect 53892 389212 53898 389224
rect 57974 389212 57980 389224
rect 53892 389184 57980 389212
rect 53892 389172 53898 389184
rect 57974 389172 57980 389184
rect 58032 389172 58038 389224
rect 41506 387948 41512 388000
rect 41564 387988 41570 388000
rect 51166 387988 51172 388000
rect 41564 387960 51172 387988
rect 41564 387948 41570 387960
rect 51166 387948 51172 387960
rect 51224 387948 51230 388000
rect 41506 387608 41512 387660
rect 41564 387648 41570 387660
rect 54018 387648 54024 387660
rect 41564 387620 54024 387648
rect 41564 387608 41570 387620
rect 54018 387608 54024 387620
rect 54076 387608 54082 387660
rect 41506 387132 41512 387184
rect 41564 387172 41570 387184
rect 49142 387172 49148 387184
rect 41564 387144 49148 387172
rect 41564 387132 41570 387144
rect 49142 387132 49148 387144
rect 49200 387132 49206 387184
rect 42794 386384 42800 386436
rect 42852 386424 42858 386436
rect 63126 386424 63132 386436
rect 42852 386396 63132 386424
rect 42852 386384 42858 386396
rect 63126 386384 63132 386396
rect 63184 386384 63190 386436
rect 675754 386384 675760 386436
rect 675812 386384 675818 386436
rect 675772 386164 675800 386384
rect 675754 386112 675760 386164
rect 675812 386112 675818 386164
rect 674466 384956 674472 385008
rect 674524 384996 674530 385008
rect 675294 384996 675300 385008
rect 674524 384968 675300 384996
rect 674524 384956 674530 384968
rect 675294 384956 675300 384968
rect 675352 384956 675358 385008
rect 675202 384072 675208 384124
rect 675260 384072 675266 384124
rect 675220 383908 675248 384072
rect 675294 383908 675300 383920
rect 675220 383880 675300 383908
rect 675294 383868 675300 383880
rect 675352 383868 675358 383920
rect 674650 383120 674656 383172
rect 674708 383160 674714 383172
rect 675386 383160 675392 383172
rect 674708 383132 675392 383160
rect 674708 383120 674714 383132
rect 675386 383120 675392 383132
rect 675444 383120 675450 383172
rect 674374 382984 674380 383036
rect 674432 383024 674438 383036
rect 674650 383024 674656 383036
rect 674432 382996 674656 383024
rect 674432 382984 674438 382996
rect 674650 382984 674656 382996
rect 674708 382984 674714 383036
rect 675018 382440 675024 382492
rect 675076 382480 675082 382492
rect 675386 382480 675392 382492
rect 675076 382452 675392 382480
rect 675076 382440 675082 382452
rect 675386 382440 675392 382452
rect 675444 382440 675450 382492
rect 674926 381896 674932 381948
rect 674984 381936 674990 381948
rect 675386 381936 675392 381948
rect 674984 381908 675392 381936
rect 674984 381896 674990 381908
rect 675386 381896 675392 381908
rect 675444 381896 675450 381948
rect 673822 379448 673828 379500
rect 673880 379488 673886 379500
rect 675294 379488 675300 379500
rect 673880 379460 675300 379488
rect 673880 379448 673886 379460
rect 675294 379448 675300 379460
rect 675352 379448 675358 379500
rect 656802 378156 656808 378208
rect 656860 378196 656866 378208
rect 670050 378196 670056 378208
rect 656860 378168 670056 378196
rect 656860 378156 656866 378168
rect 670050 378156 670056 378168
rect 670108 378156 670114 378208
rect 674006 378156 674012 378208
rect 674064 378196 674070 378208
rect 675478 378196 675484 378208
rect 674064 378168 675484 378196
rect 674064 378156 674070 378168
rect 675478 378156 675484 378168
rect 675536 378156 675542 378208
rect 673638 378088 673644 378140
rect 673696 378128 673702 378140
rect 675294 378128 675300 378140
rect 673696 378100 675300 378128
rect 673696 378088 673702 378100
rect 675294 378088 675300 378100
rect 675352 378088 675358 378140
rect 673730 376932 673736 376984
rect 673788 376972 673794 376984
rect 675478 376972 675484 376984
rect 673788 376944 675484 376972
rect 673788 376932 673794 376944
rect 675478 376932 675484 376944
rect 675536 376932 675542 376984
rect 673546 376864 673552 376916
rect 673604 376904 673610 376916
rect 675294 376904 675300 376916
rect 673604 376876 675300 376904
rect 673604 376864 673610 376876
rect 675294 376864 675300 376876
rect 675352 376864 675358 376916
rect 41598 376048 41604 376100
rect 41656 376088 41662 376100
rect 46842 376088 46848 376100
rect 41656 376060 46848 376088
rect 41656 376048 41662 376060
rect 46842 376048 46848 376060
rect 46900 376048 46906 376100
rect 49142 375368 49148 375420
rect 49200 375408 49206 375420
rect 58434 375408 58440 375420
rect 49200 375380 58440 375408
rect 49200 375368 49206 375380
rect 58434 375368 58440 375380
rect 58492 375368 58498 375420
rect 675110 374076 675116 374128
rect 675168 374116 675174 374128
rect 675294 374116 675300 374128
rect 675168 374088 675300 374116
rect 675168 374076 675174 374088
rect 675294 374076 675300 374088
rect 675352 374076 675358 374128
rect 674282 373872 674288 373924
rect 674340 373912 674346 373924
rect 675386 373912 675392 373924
rect 674340 373884 675392 373912
rect 674340 373872 674346 373884
rect 675386 373872 675392 373884
rect 675444 373872 675450 373924
rect 675294 372852 675300 372904
rect 675352 372852 675358 372904
rect 675312 372700 675340 372852
rect 675294 372648 675300 372700
rect 675352 372648 675358 372700
rect 673454 372036 673460 372088
rect 673512 372076 673518 372088
rect 675386 372076 675392 372088
rect 673512 372048 675392 372076
rect 673512 372036 673518 372048
rect 675386 372036 675392 372048
rect 675444 372036 675450 372088
rect 41506 371424 41512 371476
rect 41564 371464 41570 371476
rect 42702 371464 42708 371476
rect 41564 371436 42708 371464
rect 41564 371424 41570 371436
rect 42702 371424 42708 371436
rect 42760 371424 42766 371476
rect 674742 370744 674748 370796
rect 674800 370784 674806 370796
rect 675754 370784 675760 370796
rect 674800 370756 675760 370784
rect 674800 370744 674806 370756
rect 675754 370744 675760 370756
rect 675812 370744 675818 370796
rect 674558 370676 674564 370728
rect 674616 370716 674622 370728
rect 675662 370716 675668 370728
rect 674616 370688 675668 370716
rect 674616 370676 674622 370688
rect 675662 370676 675668 370688
rect 675720 370676 675726 370728
rect 42150 369928 42156 369980
rect 42208 369968 42214 369980
rect 42334 369968 42340 369980
rect 42208 369940 42340 369968
rect 42208 369928 42214 369940
rect 42334 369928 42340 369940
rect 42392 369928 42398 369980
rect 42150 368092 42156 368144
rect 42208 368132 42214 368144
rect 42794 368132 42800 368144
rect 42208 368104 42800 368132
rect 42208 368092 42214 368104
rect 42794 368092 42800 368104
rect 42852 368092 42858 368144
rect 42150 366800 42156 366852
rect 42208 366840 42214 366852
rect 50982 366840 50988 366852
rect 42208 366812 50988 366840
rect 42208 366800 42214 366812
rect 50982 366800 50988 366812
rect 51040 366800 51046 366852
rect 42150 366256 42156 366308
rect 42208 366296 42214 366308
rect 42886 366296 42892 366308
rect 42208 366268 42892 366296
rect 42208 366256 42214 366268
rect 42886 366256 42892 366268
rect 42944 366256 42950 366308
rect 42886 366120 42892 366172
rect 42944 366160 42950 366172
rect 43438 366160 43444 366172
rect 42944 366132 43444 366160
rect 42944 366120 42950 366132
rect 43438 366120 43444 366132
rect 43496 366120 43502 366172
rect 42150 364964 42156 365016
rect 42208 365004 42214 365016
rect 42702 365004 42708 365016
rect 42208 364976 42708 365004
rect 42208 364964 42214 364976
rect 42702 364964 42708 364976
rect 42760 364964 42766 365016
rect 42150 364420 42156 364472
rect 42208 364460 42214 364472
rect 43162 364460 43168 364472
rect 42208 364432 43168 364460
rect 42208 364420 42214 364432
rect 43162 364420 43168 364432
rect 43220 364420 43226 364472
rect 656802 364420 656808 364472
rect 656860 364460 656866 364472
rect 669038 364460 669044 364472
rect 656860 364432 669044 364460
rect 656860 364420 656866 364432
rect 669038 364420 669044 364432
rect 669096 364420 669102 364472
rect 42150 363808 42156 363860
rect 42208 363848 42214 363860
rect 43070 363848 43076 363860
rect 42208 363820 43076 363848
rect 42208 363808 42214 363820
rect 43070 363808 43076 363820
rect 43128 363808 43134 363860
rect 43070 363672 43076 363724
rect 43128 363712 43134 363724
rect 43622 363712 43628 363724
rect 43128 363684 43628 363712
rect 43128 363672 43134 363684
rect 43622 363672 43628 363684
rect 43680 363672 43686 363724
rect 42150 363128 42156 363180
rect 42208 363168 42214 363180
rect 43898 363168 43904 363180
rect 42208 363140 43904 363168
rect 42208 363128 42214 363140
rect 43898 363128 43904 363140
rect 43956 363128 43962 363180
rect 51166 361564 51172 361616
rect 51224 361604 51230 361616
rect 58434 361604 58440 361616
rect 51224 361576 58440 361604
rect 51224 361564 51230 361576
rect 58434 361564 58440 361576
rect 58492 361564 58498 361616
rect 42058 360680 42064 360732
rect 42116 360720 42122 360732
rect 43254 360720 43260 360732
rect 42116 360692 43260 360720
rect 42116 360680 42122 360692
rect 43254 360680 43260 360692
rect 43312 360680 43318 360732
rect 42150 359932 42156 359984
rect 42208 359972 42214 359984
rect 43622 359972 43628 359984
rect 42208 359944 43628 359972
rect 42208 359932 42214 359944
rect 43622 359932 43628 359944
rect 43680 359932 43686 359984
rect 42150 359456 42156 359508
rect 42208 359496 42214 359508
rect 43070 359496 43076 359508
rect 42208 359468 43076 359496
rect 42208 359456 42214 359468
rect 43070 359456 43076 359468
rect 43128 359456 43134 359508
rect 42058 358640 42064 358692
rect 42116 358680 42122 358692
rect 42978 358680 42984 358692
rect 42116 358652 42984 358680
rect 42116 358640 42122 358652
rect 42978 358640 42984 358652
rect 43036 358640 43042 358692
rect 673270 357008 673276 357060
rect 673328 357048 673334 357060
rect 675754 357048 675760 357060
rect 673328 357020 675760 357048
rect 673328 357008 673334 357020
rect 675754 357008 675760 357020
rect 675812 357008 675818 357060
rect 42058 356940 42064 356992
rect 42116 356980 42122 356992
rect 43346 356980 43352 356992
rect 42116 356952 43352 356980
rect 42116 356940 42122 356952
rect 43346 356940 43352 356952
rect 43404 356940 43410 356992
rect 670510 356464 670516 356516
rect 670568 356504 670574 356516
rect 675938 356504 675944 356516
rect 670568 356476 675944 356504
rect 670568 356464 670574 356476
rect 675938 356464 675944 356476
rect 675996 356464 676002 356516
rect 42150 356396 42156 356448
rect 42208 356436 42214 356448
rect 42886 356436 42892 356448
rect 42208 356408 42892 356436
rect 42208 356396 42214 356408
rect 42886 356396 42892 356408
rect 42944 356396 42950 356448
rect 669130 356328 669136 356380
rect 669188 356368 669194 356380
rect 676030 356368 676036 356380
rect 669188 356340 676036 356368
rect 669188 356328 669194 356340
rect 676030 356328 676036 356340
rect 676088 356328 676094 356380
rect 663886 356192 663892 356244
rect 663944 356232 663950 356244
rect 675846 356232 675852 356244
rect 663944 356204 675852 356232
rect 663944 356192 663950 356204
rect 675846 356192 675852 356204
rect 675904 356192 675910 356244
rect 673362 356124 673368 356176
rect 673420 356164 673426 356176
rect 676030 356164 676036 356176
rect 673420 356136 676036 356164
rect 673420 356124 673426 356136
rect 676030 356124 676036 356136
rect 676088 356124 676094 356176
rect 669590 356056 669596 356108
rect 669648 356096 669654 356108
rect 672994 356096 673000 356108
rect 669648 356068 673000 356096
rect 669648 356056 669654 356068
rect 672994 356056 673000 356068
rect 673052 356096 673058 356108
rect 673270 356096 673276 356108
rect 673052 356068 673276 356096
rect 673052 356056 673058 356068
rect 673270 356056 673276 356068
rect 673328 356056 673334 356108
rect 673178 355376 673184 355428
rect 673236 355416 673242 355428
rect 676030 355416 676036 355428
rect 673236 355388 676036 355416
rect 673236 355376 673242 355388
rect 676030 355376 676036 355388
rect 676088 355376 676094 355428
rect 673270 354560 673276 354612
rect 673328 354600 673334 354612
rect 676030 354600 676036 354612
rect 673328 354572 676036 354600
rect 673328 354560 673334 354572
rect 676030 354560 676036 354572
rect 676088 354560 676094 354612
rect 669498 353472 669504 353524
rect 669556 353512 669562 353524
rect 673086 353512 673092 353524
rect 669556 353484 673092 353512
rect 669556 353472 669562 353484
rect 673086 353472 673092 353484
rect 673144 353512 673150 353524
rect 673270 353512 673276 353524
rect 673144 353484 673276 353512
rect 673144 353472 673150 353484
rect 673270 353472 673276 353484
rect 673328 353472 673334 353524
rect 673822 353472 673828 353524
rect 673880 353512 673886 353524
rect 676030 353512 676036 353524
rect 673880 353484 676036 353512
rect 673880 353472 673886 353484
rect 676030 353472 676036 353484
rect 676088 353472 676094 353524
rect 669406 353336 669412 353388
rect 669464 353376 669470 353388
rect 673178 353376 673184 353388
rect 669464 353348 673184 353376
rect 669464 353336 669470 353348
rect 673178 353336 673184 353348
rect 673236 353336 673242 353388
rect 674098 353268 674104 353320
rect 674156 353308 674162 353320
rect 676030 353308 676036 353320
rect 674156 353280 676036 353308
rect 674156 353268 674162 353280
rect 676030 353268 676036 353280
rect 676088 353268 676094 353320
rect 672994 351772 673000 351824
rect 673052 351812 673058 351824
rect 673270 351812 673276 351824
rect 673052 351784 673276 351812
rect 673052 351772 673058 351784
rect 673270 351772 673276 351784
rect 673328 351772 673334 351824
rect 674190 351432 674196 351484
rect 674248 351472 674254 351484
rect 676030 351472 676036 351484
rect 674248 351444 676036 351472
rect 674248 351432 674254 351444
rect 676030 351432 676036 351444
rect 676088 351432 676094 351484
rect 673454 351024 673460 351076
rect 673512 351064 673518 351076
rect 675938 351064 675944 351076
rect 673512 351036 675944 351064
rect 673512 351024 673518 351036
rect 675938 351024 675944 351036
rect 675996 351024 676002 351076
rect 673914 350616 673920 350668
rect 673972 350656 673978 350668
rect 675938 350656 675944 350668
rect 673972 350628 675944 350656
rect 673972 350616 673978 350628
rect 675938 350616 675944 350628
rect 675996 350616 676002 350668
rect 654870 350548 654876 350600
rect 654928 350588 654934 350600
rect 669498 350588 669504 350600
rect 654928 350560 669504 350588
rect 654928 350548 654934 350560
rect 669498 350548 669504 350560
rect 669556 350548 669562 350600
rect 674282 350548 674288 350600
rect 674340 350588 674346 350600
rect 676030 350588 676036 350600
rect 674340 350560 676036 350588
rect 674340 350548 674346 350560
rect 676030 350548 676036 350560
rect 676088 350548 676094 350600
rect 673730 349800 673736 349852
rect 673788 349840 673794 349852
rect 676030 349840 676036 349852
rect 673788 349812 676036 349840
rect 673788 349800 673794 349812
rect 676030 349800 676036 349812
rect 676088 349800 676094 349852
rect 673638 348984 673644 349036
rect 673696 349024 673702 349036
rect 675938 349024 675944 349036
rect 673696 348996 675944 349024
rect 673696 348984 673702 348996
rect 675938 348984 675944 348996
rect 675996 348984 676002 349036
rect 673546 347828 673552 347880
rect 673604 347868 673610 347880
rect 675938 347868 675944 347880
rect 673604 347840 675944 347868
rect 673604 347828 673610 347840
rect 675938 347828 675944 347840
rect 675996 347828 676002 347880
rect 50982 347760 50988 347812
rect 51040 347800 51046 347812
rect 58434 347800 58440 347812
rect 51040 347772 58440 347800
rect 51040 347760 51046 347772
rect 58434 347760 58440 347772
rect 58492 347760 58498 347812
rect 674006 347760 674012 347812
rect 674064 347800 674070 347812
rect 676030 347800 676036 347812
rect 674064 347772 676036 347800
rect 674064 347760 674070 347772
rect 676030 347760 676036 347772
rect 676088 347760 676094 347812
rect 672994 347216 673000 347268
rect 673052 347256 673058 347268
rect 676030 347256 676036 347268
rect 673052 347228 676036 347256
rect 673052 347216 673058 347228
rect 676030 347216 676036 347228
rect 676088 347216 676094 347268
rect 44174 344972 44180 345024
rect 44232 345012 44238 345024
rect 48406 345012 48412 345024
rect 44232 344984 48412 345012
rect 44232 344972 44238 344984
rect 48406 344972 48412 344984
rect 48464 344972 48470 345024
rect 41506 344700 41512 344752
rect 41564 344740 41570 344752
rect 43530 344740 43536 344752
rect 41564 344712 43536 344740
rect 41564 344700 41570 344712
rect 43530 344700 43536 344712
rect 43588 344700 43594 344752
rect 41782 344428 41788 344480
rect 41840 344468 41846 344480
rect 53926 344468 53932 344480
rect 41840 344440 53932 344468
rect 41840 344428 41846 344440
rect 53926 344428 53932 344440
rect 53984 344428 53990 344480
rect 41598 344292 41604 344344
rect 41656 344332 41662 344344
rect 49234 344332 49240 344344
rect 41656 344304 49240 344332
rect 41656 344292 41662 344304
rect 49234 344292 49240 344304
rect 49292 344292 49298 344344
rect 41598 343884 41604 343936
rect 41656 343924 41662 343936
rect 51074 343924 51080 343936
rect 41656 343896 51080 343924
rect 41656 343884 41662 343896
rect 51074 343884 51080 343896
rect 51132 343884 51138 343936
rect 41782 343340 41788 343392
rect 41840 343380 41846 343392
rect 44174 343380 44180 343392
rect 41840 343352 44180 343380
rect 41840 343340 41846 343352
rect 44174 343340 44180 343352
rect 44232 343340 44238 343392
rect 674098 340960 674104 341012
rect 674156 341000 674162 341012
rect 675478 341000 675484 341012
rect 674156 340972 675484 341000
rect 674156 340960 674162 340972
rect 675478 340960 675484 340972
rect 675536 340960 675542 341012
rect 673822 339532 673828 339584
rect 673880 339572 673886 339584
rect 675478 339572 675484 339584
rect 673880 339544 675484 339572
rect 673880 339532 673886 339544
rect 675478 339532 675484 339544
rect 675536 339532 675542 339584
rect 674190 337900 674196 337952
rect 674248 337940 674254 337952
rect 675478 337940 675484 337952
rect 674248 337912 675484 337940
rect 674248 337900 674254 337912
rect 675478 337900 675484 337912
rect 675536 337900 675542 337952
rect 674282 337220 674288 337272
rect 674340 337260 674346 337272
rect 675386 337260 675392 337272
rect 674340 337232 675392 337260
rect 674340 337220 674346 337232
rect 675386 337220 675392 337232
rect 675444 337220 675450 337272
rect 48406 336744 48412 336796
rect 48464 336784 48470 336796
rect 58434 336784 58440 336796
rect 48464 336756 58440 336784
rect 48464 336744 48470 336756
rect 58434 336744 58440 336756
rect 58492 336744 58498 336796
rect 655054 336744 655060 336796
rect 655112 336784 655118 336796
rect 666922 336784 666928 336796
rect 655112 336756 666928 336784
rect 655112 336744 655118 336756
rect 666922 336744 666928 336756
rect 666980 336744 666986 336796
rect 673914 336540 673920 336592
rect 673972 336580 673978 336592
rect 675386 336580 675392 336592
rect 673972 336552 675392 336580
rect 673972 336540 673978 336552
rect 675386 336540 675392 336552
rect 675444 336540 675450 336592
rect 674006 335860 674012 335912
rect 674064 335900 674070 335912
rect 675478 335900 675484 335912
rect 674064 335872 675484 335900
rect 674064 335860 674070 335872
rect 675478 335860 675484 335872
rect 675536 335860 675542 335912
rect 673454 333548 673460 333600
rect 673512 333588 673518 333600
rect 675386 333588 675392 333600
rect 673512 333560 675392 333588
rect 673512 333548 673518 333560
rect 675386 333548 675392 333560
rect 675444 333548 675450 333600
rect 673638 332936 673644 332988
rect 673696 332976 673702 332988
rect 675386 332976 675392 332988
rect 673696 332948 675392 332976
rect 673696 332936 673702 332948
rect 675386 332936 675392 332948
rect 675444 332936 675450 332988
rect 41506 332800 41512 332852
rect 41564 332840 41570 332852
rect 46198 332840 46204 332852
rect 41564 332812 46204 332840
rect 41564 332800 41570 332812
rect 46198 332800 46204 332812
rect 46256 332800 46262 332852
rect 673730 332392 673736 332444
rect 673788 332432 673794 332444
rect 675386 332432 675392 332444
rect 673788 332404 675392 332432
rect 673788 332392 673794 332404
rect 675386 332392 675392 332404
rect 675444 332392 675450 332444
rect 673546 331576 673552 331628
rect 673604 331616 673610 331628
rect 675386 331616 675392 331628
rect 673604 331588 675392 331616
rect 673604 331576 673610 331588
rect 675386 331576 675392 331588
rect 675444 331576 675450 331628
rect 33042 330080 33048 330132
rect 33100 330120 33106 330132
rect 41874 330120 41880 330132
rect 33100 330092 41880 330120
rect 33100 330080 33106 330092
rect 41874 330080 41880 330092
rect 41932 330080 41938 330132
rect 32858 329944 32864 329996
rect 32916 329984 32922 329996
rect 42886 329984 42892 329996
rect 32916 329956 42892 329984
rect 32916 329944 32922 329956
rect 42886 329944 42892 329956
rect 42944 329944 42950 329996
rect 32950 329876 32956 329928
rect 33008 329916 33014 329928
rect 43346 329916 43352 329928
rect 33008 329888 43352 329916
rect 33008 329876 33014 329888
rect 43346 329876 43352 329888
rect 43404 329876 43410 329928
rect 32674 329808 32680 329860
rect 32732 329848 32738 329860
rect 42794 329848 42800 329860
rect 32732 329820 42800 329848
rect 32732 329808 32738 329820
rect 42794 329808 42800 329820
rect 42852 329808 42858 329860
rect 41874 326952 41880 327004
rect 41932 326952 41938 327004
rect 41892 326800 41920 326952
rect 41874 326748 41880 326800
rect 41932 326748 41938 326800
rect 42058 324912 42064 324964
rect 42116 324952 42122 324964
rect 42794 324952 42800 324964
rect 42116 324924 42800 324952
rect 42116 324912 42122 324924
rect 42794 324912 42800 324924
rect 42852 324912 42858 324964
rect 42794 324776 42800 324828
rect 42852 324816 42858 324828
rect 43070 324816 43076 324828
rect 42852 324788 43076 324816
rect 42852 324776 42858 324788
rect 43070 324776 43076 324788
rect 43128 324776 43134 324828
rect 43162 324776 43168 324828
rect 43220 324776 43226 324828
rect 43180 324624 43208 324776
rect 43162 324572 43168 324624
rect 43220 324572 43226 324624
rect 654870 323892 654876 323944
rect 654928 323932 654934 323944
rect 669130 323932 669136 323944
rect 654928 323904 669136 323932
rect 654928 323892 654934 323904
rect 669130 323892 669136 323904
rect 669188 323892 669194 323944
rect 53926 323484 53932 323536
rect 53984 323524 53990 323536
rect 58158 323524 58164 323536
rect 53984 323496 58164 323524
rect 53984 323484 53990 323496
rect 58158 323484 58164 323496
rect 58216 323484 58222 323536
rect 42150 323280 42156 323332
rect 42208 323320 42214 323332
rect 42610 323320 42616 323332
rect 42208 323292 42616 323320
rect 42208 323280 42214 323292
rect 42610 323280 42616 323292
rect 42668 323280 42674 323332
rect 42058 323076 42064 323128
rect 42116 323116 42122 323128
rect 42886 323116 42892 323128
rect 42116 323088 42892 323116
rect 42116 323076 42122 323088
rect 42886 323076 42892 323088
rect 42944 323076 42950 323128
rect 42150 321784 42156 321836
rect 42208 321824 42214 321836
rect 43162 321824 43168 321836
rect 42208 321796 43168 321824
rect 42208 321784 42214 321796
rect 43162 321784 43168 321796
rect 43220 321784 43226 321836
rect 42150 321036 42156 321088
rect 42208 321076 42214 321088
rect 43346 321076 43352 321088
rect 42208 321048 43352 321076
rect 42208 321036 42214 321048
rect 43346 321036 43352 321048
rect 43404 321036 43410 321088
rect 42150 320560 42156 320612
rect 42208 320600 42214 320612
rect 42978 320600 42984 320612
rect 42208 320572 42984 320600
rect 42208 320560 42214 320572
rect 42978 320560 42984 320572
rect 43036 320560 43042 320612
rect 42610 320084 42616 320136
rect 42668 320124 42674 320136
rect 53742 320124 53748 320136
rect 42668 320096 53748 320124
rect 42668 320084 42674 320096
rect 53742 320084 53748 320096
rect 53800 320084 53806 320136
rect 42150 317432 42156 317484
rect 42208 317472 42214 317484
rect 42794 317472 42800 317484
rect 42208 317444 42800 317472
rect 42208 317432 42214 317444
rect 42794 317432 42800 317444
rect 42852 317432 42858 317484
rect 658458 314576 658464 314628
rect 658516 314616 658522 314628
rect 671154 314616 671160 314628
rect 658516 314588 671160 314616
rect 658516 314576 658522 314588
rect 671154 314576 671160 314588
rect 671212 314576 671218 314628
rect 667014 313692 667020 313744
rect 667072 313732 667078 313744
rect 676030 313732 676036 313744
rect 667072 313704 676036 313732
rect 667072 313692 667078 313704
rect 676030 313692 676036 313704
rect 676088 313692 676094 313744
rect 663978 312876 663984 312928
rect 664036 312916 664042 312928
rect 676030 312916 676036 312928
rect 664036 312888 676036 312916
rect 664036 312876 664042 312888
rect 676030 312876 676036 312888
rect 676088 312876 676094 312928
rect 673270 312468 673276 312520
rect 673328 312508 673334 312520
rect 676030 312508 676036 312520
rect 673328 312480 676036 312508
rect 673328 312468 673334 312480
rect 676030 312468 676036 312480
rect 676088 312468 676094 312520
rect 671154 312060 671160 312112
rect 671212 312100 671218 312112
rect 672258 312100 672264 312112
rect 671212 312072 672264 312100
rect 671212 312060 671218 312072
rect 672258 312060 672264 312072
rect 672316 312100 672322 312112
rect 676030 312100 676036 312112
rect 672316 312072 676036 312100
rect 672316 312060 672322 312072
rect 676030 312060 676036 312072
rect 676088 312060 676094 312112
rect 660942 311992 660948 312044
rect 661000 312032 661006 312044
rect 676214 312032 676220 312044
rect 661000 312004 676220 312032
rect 661000 311992 661006 312004
rect 676214 311992 676220 312004
rect 676272 311992 676278 312044
rect 658366 311788 658372 311840
rect 658424 311828 658430 311840
rect 671154 311828 671160 311840
rect 658424 311800 671160 311828
rect 658424 311788 658430 311800
rect 671154 311788 671160 311800
rect 671212 311788 671218 311840
rect 673362 311652 673368 311704
rect 673420 311692 673426 311704
rect 676030 311692 676036 311704
rect 673420 311664 676036 311692
rect 673420 311652 673426 311664
rect 676030 311652 676036 311664
rect 676088 311652 676094 311704
rect 654134 311244 654140 311296
rect 654192 311284 654198 311296
rect 669406 311284 669412 311296
rect 654192 311256 669412 311284
rect 654192 311244 654198 311256
rect 669406 311244 669412 311256
rect 669464 311244 669470 311296
rect 674742 310972 674748 311024
rect 674800 311012 674806 311024
rect 676030 311012 676036 311024
rect 674800 310984 676036 311012
rect 674800 310972 674806 310984
rect 676030 310972 676036 310984
rect 676088 310972 676094 311024
rect 673178 310836 673184 310888
rect 673236 310876 673242 310888
rect 676030 310876 676036 310888
rect 673236 310848 676036 310876
rect 673236 310836 673242 310848
rect 676030 310836 676036 310848
rect 676088 310836 676094 310888
rect 655422 310428 655428 310480
rect 655480 310468 655486 310480
rect 673270 310468 673276 310480
rect 655480 310440 673276 310468
rect 655480 310428 655486 310440
rect 673270 310428 673276 310440
rect 673328 310468 673334 310480
rect 676030 310468 676036 310480
rect 673328 310440 676036 310468
rect 673328 310428 673334 310440
rect 676030 310428 676036 310440
rect 676088 310428 676094 310480
rect 673086 310020 673092 310072
rect 673144 310060 673150 310072
rect 676030 310060 676036 310072
rect 673144 310032 676036 310060
rect 673144 310020 673150 310032
rect 676030 310020 676036 310032
rect 676088 310020 676094 310072
rect 671154 309612 671160 309664
rect 671212 309652 671218 309664
rect 671890 309652 671896 309664
rect 671212 309624 671896 309652
rect 671212 309612 671218 309624
rect 671890 309612 671896 309624
rect 671948 309652 671954 309664
rect 676030 309652 676036 309664
rect 671948 309624 676036 309652
rect 671948 309612 671954 309624
rect 676030 309612 676036 309624
rect 676088 309612 676094 309664
rect 674190 309136 674196 309188
rect 674248 309176 674254 309188
rect 676030 309176 676036 309188
rect 674248 309148 676036 309176
rect 674248 309136 674254 309148
rect 676030 309136 676036 309148
rect 676088 309136 676094 309188
rect 673546 308048 673552 308100
rect 673604 308088 673610 308100
rect 676030 308088 676036 308100
rect 673604 308060 676036 308088
rect 673604 308048 673610 308060
rect 676030 308048 676036 308060
rect 676088 308048 676094 308100
rect 673454 306484 673460 306536
rect 673512 306524 673518 306536
rect 675938 306524 675944 306536
rect 673512 306496 675944 306524
rect 673512 306484 673518 306496
rect 675938 306484 675944 306496
rect 675996 306484 676002 306536
rect 674466 306416 674472 306468
rect 674524 306456 674530 306468
rect 676030 306456 676036 306468
rect 674524 306428 676036 306456
rect 674524 306416 674530 306428
rect 676030 306416 676036 306428
rect 676088 306416 676094 306468
rect 673914 306348 673920 306400
rect 673972 306388 673978 306400
rect 676122 306388 676128 306400
rect 673972 306360 676128 306388
rect 673972 306348 673978 306360
rect 676122 306348 676128 306360
rect 676180 306348 676186 306400
rect 674650 306008 674656 306060
rect 674708 306048 674714 306060
rect 676030 306048 676036 306060
rect 674708 306020 676036 306048
rect 674708 306008 674714 306020
rect 676030 306008 676036 306020
rect 676088 306008 676094 306060
rect 673638 305056 673644 305108
rect 673696 305096 673702 305108
rect 676122 305096 676128 305108
rect 673696 305068 676128 305096
rect 673696 305056 673702 305068
rect 676122 305056 676128 305068
rect 676180 305056 676186 305108
rect 673730 304648 673736 304700
rect 673788 304688 673794 304700
rect 676122 304688 676128 304700
rect 673788 304660 676128 304688
rect 673788 304648 673794 304660
rect 676122 304648 676128 304660
rect 676180 304648 676186 304700
rect 673822 303832 673828 303884
rect 673880 303872 673886 303884
rect 675846 303872 675852 303884
rect 673880 303844 675852 303872
rect 673880 303832 673886 303844
rect 675846 303832 675852 303844
rect 675904 303832 675910 303884
rect 674006 303764 674012 303816
rect 674064 303804 674070 303816
rect 675938 303804 675944 303816
rect 674064 303776 675944 303804
rect 674064 303764 674070 303776
rect 675938 303764 675944 303776
rect 675996 303764 676002 303816
rect 674558 303696 674564 303748
rect 674616 303736 674622 303748
rect 676122 303736 676128 303748
rect 674616 303708 676128 303736
rect 674616 303696 674622 303708
rect 676122 303696 676128 303708
rect 676180 303696 676186 303748
rect 41506 301588 41512 301640
rect 41564 301628 41570 301640
rect 49142 301628 49148 301640
rect 41564 301600 49148 301628
rect 41564 301588 41570 301600
rect 49142 301588 49148 301600
rect 49200 301588 49206 301640
rect 675202 300976 675208 301028
rect 675260 301016 675266 301028
rect 675478 301016 675484 301028
rect 675260 300988 675484 301016
rect 675260 300976 675266 300988
rect 675478 300976 675484 300988
rect 675536 300976 675542 301028
rect 41782 300908 41788 300960
rect 41840 300948 41846 300960
rect 51166 300948 51172 300960
rect 41840 300920 51172 300948
rect 41840 300908 41846 300920
rect 51166 300908 51172 300920
rect 51224 300908 51230 300960
rect 673086 300840 673092 300892
rect 673144 300880 673150 300892
rect 678974 300880 678980 300892
rect 673144 300852 678980 300880
rect 673144 300840 673150 300852
rect 678974 300840 678980 300852
rect 679032 300840 679038 300892
rect 655606 298256 655612 298308
rect 655664 298296 655670 298308
rect 669590 298296 669596 298308
rect 655664 298268 669596 298296
rect 655664 298256 655670 298268
rect 669590 298256 669596 298268
rect 669648 298256 669654 298308
rect 675754 296148 675760 296200
rect 675812 296148 675818 296200
rect 675772 295996 675800 296148
rect 675754 295944 675760 295996
rect 675812 295944 675818 295996
rect 675202 295060 675208 295112
rect 675260 295100 675266 295112
rect 675386 295100 675392 295112
rect 675260 295072 675392 295100
rect 675260 295060 675266 295072
rect 675386 295060 675392 295072
rect 675444 295060 675450 295112
rect 674190 294516 674196 294568
rect 674248 294556 674254 294568
rect 675386 294556 675392 294568
rect 674248 294528 675392 294556
rect 674248 294516 674254 294528
rect 675386 294516 675392 294528
rect 675444 294516 675450 294568
rect 674466 292884 674472 292936
rect 674524 292924 674530 292936
rect 675386 292924 675392 292936
rect 674524 292896 675392 292924
rect 674524 292884 674530 292896
rect 675386 292884 675392 292896
rect 675444 292884 675450 292936
rect 674650 292272 674656 292324
rect 674708 292312 674714 292324
rect 675386 292312 675392 292324
rect 674708 292284 675392 292312
rect 674708 292272 674714 292284
rect 675386 292272 675392 292284
rect 675444 292272 675450 292324
rect 41782 292000 41788 292052
rect 41840 292040 41846 292052
rect 43346 292040 43352 292052
rect 41840 292012 43352 292040
rect 41840 292000 41846 292012
rect 43346 292000 43352 292012
rect 43404 292000 43410 292052
rect 41782 291592 41788 291644
rect 41840 291632 41846 291644
rect 43530 291632 43536 291644
rect 41840 291604 43536 291632
rect 41840 291592 41846 291604
rect 43530 291592 43536 291604
rect 43588 291592 43594 291644
rect 41874 291116 41880 291168
rect 41932 291156 41938 291168
rect 42702 291156 42708 291168
rect 41932 291128 42708 291156
rect 41932 291116 41938 291128
rect 42702 291116 42708 291128
rect 42760 291116 42766 291168
rect 674558 291048 674564 291100
rect 674616 291088 674622 291100
rect 675386 291088 675392 291100
rect 674616 291060 675392 291088
rect 674616 291048 674622 291060
rect 675386 291048 675392 291060
rect 675444 291048 675450 291100
rect 41782 289824 41788 289876
rect 41840 289864 41846 289876
rect 43162 289864 43168 289876
rect 41840 289836 43168 289864
rect 41840 289824 41846 289836
rect 43162 289824 43168 289836
rect 43220 289824 43226 289876
rect 673914 288532 673920 288584
rect 673972 288572 673978 288584
rect 675386 288572 675392 288584
rect 673972 288544 675392 288572
rect 673972 288532 673978 288544
rect 675386 288532 675392 288544
rect 675444 288532 675450 288584
rect 674006 287920 674012 287972
rect 674064 287960 674070 287972
rect 675386 287960 675392 287972
rect 674064 287932 675392 287960
rect 674064 287920 674070 287932
rect 675386 287920 675392 287932
rect 675444 287920 675450 287972
rect 673730 287172 673736 287224
rect 673788 287212 673794 287224
rect 675478 287212 675484 287224
rect 673788 287184 675484 287212
rect 673788 287172 673794 287184
rect 675478 287172 675484 287184
rect 675536 287172 675542 287224
rect 673822 286560 673828 286612
rect 673880 286600 673886 286612
rect 675386 286600 675392 286612
rect 673880 286572 675392 286600
rect 673880 286560 673886 286572
rect 675386 286560 675392 286572
rect 675444 286560 675450 286612
rect 32674 285744 32680 285796
rect 32732 285784 32738 285796
rect 42794 285784 42800 285796
rect 32732 285756 42800 285784
rect 32732 285744 32738 285756
rect 42794 285744 42800 285756
rect 42852 285744 42858 285796
rect 32858 285676 32864 285728
rect 32916 285716 32922 285728
rect 42978 285716 42984 285728
rect 32916 285688 42984 285716
rect 32916 285676 32922 285688
rect 42978 285676 42984 285688
rect 43036 285676 43042 285728
rect 32766 285608 32772 285660
rect 32824 285648 32830 285660
rect 42886 285648 42892 285660
rect 32824 285620 42892 285648
rect 32824 285608 32830 285620
rect 42886 285608 42892 285620
rect 42944 285608 42950 285660
rect 673638 285540 673644 285592
rect 673696 285580 673702 285592
rect 675478 285580 675484 285592
rect 673696 285552 675484 285580
rect 673696 285540 673702 285552
rect 675478 285540 675484 285552
rect 675536 285540 675542 285592
rect 655330 284724 655336 284776
rect 655388 284764 655394 284776
rect 670510 284764 670516 284776
rect 655388 284736 670516 284764
rect 655388 284724 655394 284736
rect 670510 284724 670516 284736
rect 670568 284724 670574 284776
rect 673546 283704 673552 283756
rect 673604 283744 673610 283756
rect 675478 283744 675484 283756
rect 673604 283716 675484 283744
rect 673604 283704 673610 283716
rect 675478 283704 675484 283716
rect 675536 283704 675542 283756
rect 42150 283568 42156 283620
rect 42208 283608 42214 283620
rect 42702 283608 42708 283620
rect 42208 283580 42708 283608
rect 42208 283568 42214 283580
rect 42702 283568 42708 283580
rect 42760 283568 42766 283620
rect 42426 283296 42432 283348
rect 42484 283336 42490 283348
rect 42702 283336 42708 283348
rect 42484 283308 42708 283336
rect 42484 283296 42490 283308
rect 42702 283296 42708 283308
rect 42760 283296 42766 283348
rect 673454 281868 673460 281920
rect 673512 281908 673518 281920
rect 675386 281908 675392 281920
rect 673512 281880 675392 281908
rect 673512 281868 673518 281880
rect 675386 281868 675392 281880
rect 675444 281868 675450 281920
rect 42150 281732 42156 281784
rect 42208 281772 42214 281784
rect 42794 281772 42800 281784
rect 42208 281744 42800 281772
rect 42208 281732 42214 281744
rect 42794 281732 42800 281744
rect 42852 281732 42858 281784
rect 42150 281052 42156 281104
rect 42208 281092 42214 281104
rect 49050 281092 49056 281104
rect 42208 281064 49056 281092
rect 42208 281052 42214 281064
rect 49050 281052 49056 281064
rect 49108 281052 49114 281104
rect 42150 279828 42156 279880
rect 42208 279868 42214 279880
rect 43070 279868 43076 279880
rect 42208 279840 43076 279868
rect 42208 279828 42214 279840
rect 43070 279828 43076 279840
rect 43128 279828 43134 279880
rect 42058 278604 42064 278656
rect 42116 278644 42122 278656
rect 43162 278644 43168 278656
rect 42116 278616 43168 278644
rect 42116 278604 42122 278616
rect 43162 278604 43168 278616
rect 43220 278604 43226 278656
rect 46474 278536 46480 278588
rect 46532 278576 46538 278588
rect 672810 278576 672816 278588
rect 46532 278548 672816 278576
rect 46532 278536 46538 278548
rect 672810 278536 672816 278548
rect 672868 278536 672874 278588
rect 46566 278468 46572 278520
rect 46624 278508 46630 278520
rect 670234 278508 670240 278520
rect 46624 278480 670240 278508
rect 46624 278468 46630 278480
rect 670234 278468 670240 278480
rect 670292 278468 670298 278520
rect 46750 278400 46756 278452
rect 46808 278440 46814 278452
rect 670418 278440 670424 278452
rect 46808 278412 670424 278440
rect 46808 278400 46814 278412
rect 670418 278400 670424 278412
rect 670476 278400 670482 278452
rect 62574 278332 62580 278384
rect 62632 278372 62638 278384
rect 670142 278372 670148 278384
rect 62632 278344 670148 278372
rect 62632 278332 62638 278344
rect 670142 278332 670148 278344
rect 670200 278332 670206 278384
rect 62758 278264 62764 278316
rect 62816 278304 62822 278316
rect 668762 278304 668768 278316
rect 62816 278276 668768 278304
rect 62816 278264 62822 278276
rect 668762 278264 668768 278276
rect 668820 278264 668826 278316
rect 62942 278196 62948 278248
rect 63000 278236 63006 278248
rect 670326 278236 670332 278248
rect 63000 278208 670332 278236
rect 63000 278196 63006 278208
rect 670326 278196 670332 278208
rect 670384 278196 670390 278248
rect 62390 278128 62396 278180
rect 62448 278168 62454 278180
rect 669682 278168 669688 278180
rect 62448 278140 669688 278168
rect 62448 278128 62454 278140
rect 669682 278128 669688 278140
rect 669740 278128 669746 278180
rect 63126 278060 63132 278112
rect 63184 278100 63190 278112
rect 669774 278100 669780 278112
rect 63184 278072 669780 278100
rect 63184 278060 63190 278072
rect 669774 278060 669780 278072
rect 669832 278060 669838 278112
rect 63218 277992 63224 278044
rect 63276 278032 63282 278044
rect 669866 278032 669872 278044
rect 63276 278004 669872 278032
rect 63276 277992 63282 278004
rect 669866 277992 669872 278004
rect 669924 277992 669930 278044
rect 63310 277924 63316 277976
rect 63368 277964 63374 277976
rect 669958 277964 669964 277976
rect 63368 277936 669964 277964
rect 63368 277924 63374 277936
rect 669958 277924 669964 277936
rect 670016 277924 670022 277976
rect 42150 277856 42156 277908
rect 42208 277896 42214 277908
rect 43254 277896 43260 277908
rect 42208 277868 43260 277896
rect 42208 277856 42214 277868
rect 43254 277856 43260 277868
rect 43312 277856 43318 277908
rect 42150 277380 42156 277432
rect 42208 277420 42214 277432
rect 43530 277420 43536 277432
rect 42208 277392 43536 277420
rect 42208 277380 42214 277392
rect 43530 277380 43536 277392
rect 43588 277380 43594 277432
rect 42058 276700 42064 276752
rect 42116 276740 42122 276752
rect 42978 276740 42984 276752
rect 42116 276712 42984 276740
rect 42116 276700 42122 276712
rect 42978 276700 42984 276712
rect 43036 276700 43042 276752
rect 345106 275952 345112 276004
rect 345164 275992 345170 276004
rect 471330 275992 471336 276004
rect 345164 275964 471336 275992
rect 345164 275952 345170 275964
rect 471330 275952 471336 275964
rect 471388 275952 471394 276004
rect 343726 275884 343732 275936
rect 343784 275924 343790 275936
rect 467834 275924 467840 275936
rect 343784 275896 467840 275924
rect 343784 275884 343790 275896
rect 467834 275884 467840 275896
rect 467892 275884 467898 275936
rect 349062 275816 349068 275868
rect 349120 275856 349126 275868
rect 482002 275856 482008 275868
rect 349120 275828 482008 275856
rect 349120 275816 349126 275828
rect 482002 275816 482008 275828
rect 482060 275816 482066 275868
rect 350350 275748 350356 275800
rect 350408 275788 350414 275800
rect 485498 275788 485504 275800
rect 350408 275760 485504 275788
rect 350408 275748 350414 275760
rect 485498 275748 485504 275760
rect 485556 275748 485562 275800
rect 354398 275680 354404 275732
rect 354456 275720 354462 275732
rect 496170 275720 496176 275732
rect 354456 275692 496176 275720
rect 354456 275680 354462 275692
rect 496170 275680 496176 275692
rect 496228 275680 496234 275732
rect 355778 275612 355784 275664
rect 355836 275652 355842 275664
rect 499758 275652 499764 275664
rect 355836 275624 499764 275652
rect 355836 275612 355842 275624
rect 499758 275612 499764 275624
rect 499816 275612 499822 275664
rect 358446 275544 358452 275596
rect 358504 275584 358510 275596
rect 506842 275584 506848 275596
rect 358504 275556 506848 275584
rect 358504 275544 358510 275556
rect 506842 275544 506848 275556
rect 506900 275544 506906 275596
rect 361114 275476 361120 275528
rect 361172 275516 361178 275528
rect 513926 275516 513932 275528
rect 361172 275488 513932 275516
rect 361172 275476 361178 275488
rect 513926 275476 513932 275488
rect 513984 275476 513990 275528
rect 364058 275408 364064 275460
rect 364116 275448 364122 275460
rect 521010 275448 521016 275460
rect 364116 275420 521016 275448
rect 364116 275408 364122 275420
rect 521010 275408 521016 275420
rect 521068 275408 521074 275460
rect 366450 275340 366456 275392
rect 366508 275380 366514 275392
rect 528094 275380 528100 275392
rect 366508 275352 528100 275380
rect 366508 275340 366514 275352
rect 528094 275340 528100 275352
rect 528152 275340 528158 275392
rect 369118 275272 369124 275324
rect 369176 275312 369182 275324
rect 535178 275312 535184 275324
rect 369176 275284 535184 275312
rect 369176 275272 369182 275284
rect 535178 275272 535184 275284
rect 535236 275272 535242 275324
rect 371786 275204 371792 275256
rect 371844 275244 371850 275256
rect 542262 275244 542268 275256
rect 371844 275216 542268 275244
rect 371844 275204 371850 275216
rect 542262 275204 542268 275216
rect 542320 275204 542326 275256
rect 374914 275136 374920 275188
rect 374972 275176 374978 275188
rect 550542 275176 550548 275188
rect 374972 275148 550548 275176
rect 374972 275136 374978 275148
rect 550542 275136 550548 275148
rect 550600 275136 550606 275188
rect 377582 275068 377588 275120
rect 377640 275108 377646 275120
rect 557626 275108 557632 275120
rect 377640 275080 557632 275108
rect 377640 275068 377646 275080
rect 557626 275068 557632 275080
rect 557684 275068 557690 275120
rect 380250 275000 380256 275052
rect 380308 275040 380314 275052
rect 564710 275040 564716 275052
rect 380308 275012 564716 275040
rect 380308 275000 380314 275012
rect 564710 275000 564716 275012
rect 564768 275000 564774 275052
rect 382918 274932 382924 274984
rect 382976 274972 382982 274984
rect 571794 274972 571800 274984
rect 382976 274944 571800 274972
rect 382976 274932 382982 274944
rect 571794 274932 571800 274944
rect 571852 274932 571858 274984
rect 385586 274864 385592 274916
rect 385644 274904 385650 274916
rect 578878 274904 578884 274916
rect 385644 274876 578884 274904
rect 385644 274864 385650 274876
rect 578878 274864 578884 274876
rect 578936 274864 578942 274916
rect 318886 274796 318892 274848
rect 318944 274836 318950 274848
rect 401594 274836 401600 274848
rect 318944 274808 401600 274836
rect 318944 274796 318950 274808
rect 401594 274796 401600 274808
rect 401652 274796 401658 274848
rect 403894 274796 403900 274848
rect 403952 274836 403958 274848
rect 403952 274808 411392 274836
rect 403952 274796 403958 274808
rect 320174 274728 320180 274780
rect 320232 274768 320238 274780
rect 405182 274768 405188 274780
rect 320232 274740 405188 274768
rect 320232 274728 320238 274740
rect 405182 274728 405188 274740
rect 405240 274728 405246 274780
rect 406562 274728 406568 274780
rect 406620 274768 406626 274780
rect 411364 274768 411392 274808
rect 411438 274796 411444 274848
rect 411496 274836 411502 274848
rect 620278 274836 620284 274848
rect 411496 274808 620284 274836
rect 411496 274796 411502 274808
rect 620278 274796 620284 274808
rect 620336 274796 620342 274848
rect 627362 274768 627368 274780
rect 406620 274740 411300 274768
rect 411364 274740 627368 274768
rect 406620 274728 406626 274740
rect 321002 274660 321008 274712
rect 321060 274700 321066 274712
rect 407482 274700 407488 274712
rect 321060 274672 407488 274700
rect 321060 274660 321066 274672
rect 407482 274660 407488 274672
rect 407540 274660 407546 274712
rect 409230 274660 409236 274712
rect 409288 274700 409294 274712
rect 411272 274700 411300 274740
rect 627362 274728 627368 274740
rect 627420 274728 627426 274780
rect 634446 274700 634452 274712
rect 409288 274672 411208 274700
rect 411272 274672 634452 274700
rect 409288 274660 409294 274672
rect 322842 274592 322848 274644
rect 322900 274632 322906 274644
rect 411070 274632 411076 274644
rect 322900 274604 411076 274632
rect 322900 274592 322906 274604
rect 411070 274592 411076 274604
rect 411128 274592 411134 274644
rect 411180 274632 411208 274672
rect 634446 274660 634452 274672
rect 634504 274660 634510 274712
rect 641622 274632 641628 274644
rect 411180 274604 641628 274632
rect 641622 274592 641628 274604
rect 641680 274592 641686 274644
rect 342530 274524 342536 274576
rect 342588 274564 342594 274576
rect 464246 274564 464252 274576
rect 342588 274536 464252 274564
rect 342588 274524 342594 274536
rect 464246 274524 464252 274536
rect 464304 274524 464310 274576
rect 341058 274456 341064 274508
rect 341116 274496 341122 274508
rect 460658 274496 460664 274508
rect 341116 274468 460664 274496
rect 341116 274456 341122 274468
rect 460658 274456 460664 274468
rect 460716 274456 460722 274508
rect 337102 274388 337108 274440
rect 337160 274428 337166 274440
rect 450078 274428 450084 274440
rect 337160 274400 450084 274428
rect 337160 274388 337166 274400
rect 450078 274388 450084 274400
rect 450136 274388 450142 274440
rect 335722 274320 335728 274372
rect 335780 274360 335786 274372
rect 446490 274360 446496 274372
rect 335780 274332 446496 274360
rect 335780 274320 335786 274332
rect 446490 274320 446496 274332
rect 446548 274320 446554 274372
rect 42150 274252 42156 274304
rect 42208 274292 42214 274304
rect 42886 274292 42892 274304
rect 42208 274264 42892 274292
rect 42208 274252 42214 274264
rect 42886 274252 42892 274264
rect 42944 274252 42950 274304
rect 334342 274252 334348 274304
rect 334400 274292 334406 274304
rect 427078 274292 427084 274304
rect 334400 274264 427084 274292
rect 334400 274252 334406 274264
rect 427078 274252 427084 274264
rect 427136 274252 427142 274304
rect 333422 274184 333428 274236
rect 333480 274224 333486 274236
rect 439406 274224 439412 274236
rect 333480 274196 439412 274224
rect 333480 274184 333486 274196
rect 439406 274184 439412 274196
rect 439464 274184 439470 274236
rect 332134 274116 332140 274168
rect 332192 274156 332198 274168
rect 437014 274156 437020 274168
rect 332192 274128 437020 274156
rect 332192 274116 332198 274128
rect 437014 274116 437020 274128
rect 437072 274116 437078 274168
rect 351822 274048 351828 274100
rect 351880 274088 351886 274100
rect 432322 274088 432328 274100
rect 351880 274060 432328 274088
rect 351880 274048 351886 274060
rect 432322 274048 432328 274060
rect 432380 274048 432386 274100
rect 331674 273980 331680 274032
rect 331732 274020 331738 274032
rect 435910 274020 435916 274032
rect 331732 273992 435916 274020
rect 331732 273980 331738 273992
rect 435910 273980 435916 273992
rect 435968 273980 435974 274032
rect 327718 273912 327724 273964
rect 327776 273952 327782 273964
rect 425238 273952 425244 273964
rect 327776 273924 425244 273952
rect 327776 273912 327782 273924
rect 425238 273912 425244 273924
rect 425296 273912 425302 273964
rect 329098 273844 329104 273896
rect 329156 273884 329162 273896
rect 428826 273884 428832 273896
rect 329156 273856 428832 273884
rect 329156 273844 329162 273856
rect 428826 273844 428832 273856
rect 428884 273844 428890 273896
rect 326798 273776 326804 273828
rect 326856 273816 326862 273828
rect 326856 273788 419534 273816
rect 326856 273776 326862 273788
rect 42058 273708 42064 273760
rect 42116 273748 42122 273760
rect 42702 273748 42708 273760
rect 42116 273720 42708 273748
rect 42116 273708 42122 273720
rect 42702 273708 42708 273720
rect 42760 273708 42766 273760
rect 325418 273708 325424 273760
rect 325476 273748 325482 273760
rect 418154 273748 418160 273760
rect 325476 273720 418160 273748
rect 325476 273708 325482 273720
rect 418154 273708 418160 273720
rect 418212 273708 418218 273760
rect 326338 273640 326344 273692
rect 326396 273680 326402 273692
rect 419506 273680 419534 273788
rect 427078 273776 427084 273828
rect 427136 273816 427142 273828
rect 442994 273816 443000 273828
rect 427136 273788 443000 273816
rect 427136 273776 427142 273788
rect 442994 273776 443000 273788
rect 443052 273776 443058 273828
rect 422846 273680 422852 273692
rect 326396 273652 409828 273680
rect 419506 273652 422852 273680
rect 326396 273640 326402 273652
rect 323670 273572 323676 273624
rect 323728 273612 323734 273624
rect 409800 273612 409828 273652
rect 422846 273640 422852 273652
rect 422904 273640 422910 273692
rect 323728 273584 400214 273612
rect 409800 273584 419534 273612
rect 323728 273572 323734 273584
rect 330386 273504 330392 273556
rect 330444 273544 330450 273556
rect 351822 273544 351828 273556
rect 330444 273516 351828 273544
rect 330444 273504 330450 273516
rect 351822 273504 351828 273516
rect 351880 273504 351886 273556
rect 400186 273544 400214 273584
rect 414566 273544 414572 273556
rect 400186 273516 414572 273544
rect 414566 273504 414572 273516
rect 414624 273504 414630 273556
rect 419506 273544 419534 273584
rect 421650 273544 421656 273556
rect 419506 273516 421656 273544
rect 421650 273504 421656 273516
rect 421708 273504 421714 273556
rect 401134 273436 401140 273488
rect 401192 273476 401198 273488
rect 411438 273476 411444 273488
rect 401192 273448 411444 273476
rect 401192 273436 401198 273448
rect 411438 273436 411444 273448
rect 411496 273436 411502 273488
rect 225874 273204 225880 273216
rect 168346 273176 225880 273204
rect 155678 273096 155684 273148
rect 155736 273136 155742 273148
rect 168346 273136 168374 273176
rect 225874 273164 225880 273176
rect 225932 273164 225938 273216
rect 263226 273164 263232 273216
rect 263284 273204 263290 273216
rect 266722 273204 266728 273216
rect 263284 273176 266728 273204
rect 263284 273164 263290 273176
rect 266722 273164 266728 273176
rect 266780 273164 266786 273216
rect 292114 273164 292120 273216
rect 292172 273204 292178 273216
rect 330662 273204 330668 273216
rect 292172 273176 330668 273204
rect 292172 273164 292178 273176
rect 330662 273164 330668 273176
rect 330720 273164 330726 273216
rect 339494 273164 339500 273216
rect 339552 273204 339558 273216
rect 344830 273204 344836 273216
rect 339552 273176 344836 273204
rect 339552 273164 339558 273176
rect 344830 273164 344836 273176
rect 344888 273164 344894 273216
rect 362770 273164 362776 273216
rect 362828 273204 362834 273216
rect 491478 273204 491484 273216
rect 362828 273176 491484 273204
rect 362828 273164 362834 273176
rect 491478 273164 491484 273176
rect 491536 273164 491542 273216
rect 155736 273108 168374 273136
rect 155736 273096 155742 273108
rect 177850 273096 177856 273148
rect 177908 273136 177914 273148
rect 177908 273108 226334 273136
rect 177908 273096 177914 273108
rect 149790 273028 149796 273080
rect 149848 273068 149854 273080
rect 224402 273068 224408 273080
rect 149848 273040 224408 273068
rect 149848 273028 149854 273040
rect 224402 273028 224408 273040
rect 224460 273028 224466 273080
rect 150986 272960 150992 273012
rect 151044 273000 151050 273012
rect 223942 273000 223948 273012
rect 151044 272972 223948 273000
rect 151044 272960 151050 272972
rect 223942 272960 223948 272972
rect 224000 272960 224006 273012
rect 42150 272892 42156 272944
rect 42208 272932 42214 272944
rect 43346 272932 43352 272944
rect 42208 272904 43352 272932
rect 42208 272892 42214 272904
rect 43346 272892 43352 272904
rect 43404 272892 43410 272944
rect 143902 272892 143908 272944
rect 143960 272932 143966 272944
rect 221274 272932 221280 272944
rect 143960 272904 221280 272932
rect 143960 272892 143966 272904
rect 221274 272892 221280 272904
rect 221332 272892 221338 272944
rect 148594 272824 148600 272876
rect 148652 272864 148658 272876
rect 223206 272864 223212 272876
rect 148652 272836 223212 272864
rect 148652 272824 148658 272836
rect 223206 272824 223212 272836
rect 223264 272824 223270 272876
rect 146202 272756 146208 272808
rect 146260 272796 146266 272808
rect 223022 272796 223028 272808
rect 146260 272768 223028 272796
rect 146260 272756 146266 272768
rect 223022 272756 223028 272768
rect 223080 272756 223086 272808
rect 145006 272688 145012 272740
rect 145064 272728 145070 272740
rect 222194 272728 222200 272740
rect 145064 272700 222200 272728
rect 145064 272688 145070 272700
rect 222194 272688 222200 272700
rect 222252 272688 222258 272740
rect 139118 272620 139124 272672
rect 139176 272660 139182 272672
rect 220354 272660 220360 272672
rect 139176 272632 220360 272660
rect 139176 272620 139182 272632
rect 220354 272620 220360 272632
rect 220412 272620 220418 272672
rect 136818 272552 136824 272604
rect 136876 272592 136882 272604
rect 218606 272592 218612 272604
rect 136876 272564 218612 272592
rect 136876 272552 136882 272564
rect 218606 272552 218612 272564
rect 218664 272552 218670 272604
rect 137922 272484 137928 272536
rect 137980 272524 137986 272536
rect 219434 272524 219440 272536
rect 137980 272496 219440 272524
rect 137980 272484 137986 272496
rect 219434 272484 219440 272496
rect 219492 272484 219498 272536
rect 132034 272416 132040 272468
rect 132092 272456 132098 272468
rect 217686 272456 217692 272468
rect 132092 272428 217692 272456
rect 132092 272416 132098 272428
rect 217686 272416 217692 272428
rect 217744 272416 217750 272468
rect 129642 272348 129648 272400
rect 129700 272388 129706 272400
rect 215662 272388 215668 272400
rect 129700 272360 215668 272388
rect 129700 272348 129706 272360
rect 215662 272348 215668 272360
rect 215720 272348 215726 272400
rect 124950 272280 124956 272332
rect 125008 272320 125014 272332
rect 215018 272320 215024 272332
rect 125008 272292 215024 272320
rect 125008 272280 125014 272292
rect 215018 272280 215024 272292
rect 215076 272280 215082 272332
rect 117866 272212 117872 272264
rect 117924 272252 117930 272264
rect 205542 272252 205548 272264
rect 117924 272224 205548 272252
rect 117924 272212 117930 272224
rect 205542 272212 205548 272224
rect 205600 272212 205606 272264
rect 226306 272252 226334 273108
rect 264422 273096 264428 273148
rect 264480 273136 264486 273148
rect 267182 273136 267188 273148
rect 264480 273108 267188 273136
rect 264480 273096 264486 273108
rect 267182 273096 267188 273108
rect 267240 273096 267246 273148
rect 292574 273096 292580 273148
rect 292632 273136 292638 273148
rect 331858 273136 331864 273148
rect 292632 273108 331864 273136
rect 292632 273096 292638 273108
rect 331858 273096 331864 273108
rect 331916 273096 331922 273148
rect 331950 273096 331956 273148
rect 332008 273136 332014 273148
rect 337746 273136 337752 273148
rect 332008 273108 337752 273136
rect 332008 273096 332014 273108
rect 337746 273096 337752 273108
rect 337804 273096 337810 273148
rect 355318 273096 355324 273148
rect 355376 273136 355382 273148
rect 498562 273136 498568 273148
rect 355376 273108 362816 273136
rect 355376 273096 355382 273108
rect 243170 273028 243176 273080
rect 243228 273068 243234 273080
rect 259178 273068 259184 273080
rect 243228 273040 259184 273068
rect 243228 273028 243234 273040
rect 259178 273028 259184 273040
rect 259236 273028 259242 273080
rect 260926 273028 260932 273080
rect 260984 273068 260990 273080
rect 265802 273068 265808 273080
rect 260984 273040 265808 273068
rect 260984 273028 260990 273040
rect 265802 273028 265808 273040
rect 265860 273028 265866 273080
rect 293402 273028 293408 273080
rect 293460 273068 293466 273080
rect 334158 273068 334164 273080
rect 293460 273040 334164 273068
rect 293460 273028 293466 273040
rect 334158 273028 334164 273040
rect 334216 273028 334222 273080
rect 358814 273028 358820 273080
rect 358872 273068 358878 273080
rect 362788 273068 362816 273108
rect 363064 273108 498568 273136
rect 363064 273068 363092 273108
rect 498562 273096 498568 273108
rect 498620 273096 498626 273148
rect 358872 273040 362724 273068
rect 362788 273040 363092 273068
rect 358872 273028 358878 273040
rect 293862 272960 293868 273012
rect 293920 273000 293926 273012
rect 335354 273000 335360 273012
rect 293920 272972 335360 273000
rect 293920 272960 293926 272972
rect 335354 272960 335360 272972
rect 335412 272960 335418 273012
rect 344002 272960 344008 273012
rect 344060 273000 344066 273012
rect 362586 273000 362592 273012
rect 344060 272972 362592 273000
rect 344060 272960 344066 272972
rect 362586 272960 362592 272972
rect 362644 272960 362650 273012
rect 362696 273000 362724 273040
rect 363138 273028 363144 273080
rect 363196 273068 363202 273080
rect 497366 273068 497372 273080
rect 363196 273040 497372 273068
rect 363196 273028 363202 273040
rect 497366 273028 497372 273040
rect 497424 273028 497430 273080
rect 498838 273028 498844 273080
rect 498896 273068 498902 273080
rect 617978 273068 617984 273080
rect 498896 273040 617984 273068
rect 498896 273028 498902 273040
rect 617978 273028 617984 273040
rect 618036 273028 618042 273080
rect 504450 273000 504456 273012
rect 362696 272972 504456 273000
rect 504450 272960 504456 272972
rect 504508 272960 504514 273012
rect 239582 272892 239588 272944
rect 239640 272932 239646 272944
rect 257798 272932 257804 272944
rect 239640 272904 257804 272932
rect 239640 272892 239646 272904
rect 257798 272892 257804 272904
rect 257856 272892 257862 272944
rect 304902 272892 304908 272944
rect 304960 272932 304966 272944
rect 332502 272932 332508 272944
rect 304960 272904 332508 272932
rect 304960 272892 304966 272904
rect 332502 272892 332508 272904
rect 332560 272892 332566 272944
rect 357986 272892 357992 272944
rect 358044 272932 358050 272944
rect 505646 272932 505652 272944
rect 358044 272904 505652 272932
rect 358044 272892 358050 272904
rect 505646 272892 505652 272904
rect 505704 272892 505710 272944
rect 236086 272824 236092 272876
rect 236144 272864 236150 272876
rect 256418 272864 256424 272876
rect 236144 272836 256424 272864
rect 236144 272824 236150 272836
rect 256418 272824 256424 272836
rect 256476 272824 256482 272876
rect 307846 272824 307852 272876
rect 307904 272864 307910 272876
rect 348418 272864 348424 272876
rect 307904 272836 348424 272864
rect 307904 272824 307910 272836
rect 348418 272824 348424 272836
rect 348476 272824 348482 272876
rect 354858 272824 354864 272876
rect 354916 272864 354922 272876
rect 362862 272864 362868 272876
rect 354916 272836 362868 272864
rect 354916 272824 354922 272836
rect 362862 272824 362868 272836
rect 362920 272824 362926 272876
rect 512730 272864 512736 272876
rect 362972 272836 512736 272864
rect 234890 272756 234896 272808
rect 234948 272796 234954 272808
rect 256050 272796 256056 272808
rect 234948 272768 256056 272796
rect 234948 272756 234954 272768
rect 256050 272756 256056 272768
rect 256108 272756 256114 272808
rect 300762 272756 300768 272808
rect 300820 272796 300826 272808
rect 353110 272796 353116 272808
rect 300820 272768 353116 272796
rect 300820 272756 300826 272768
rect 353110 272756 353116 272768
rect 353168 272756 353174 272808
rect 360654 272756 360660 272808
rect 360712 272796 360718 272808
rect 362972 272796 363000 272836
rect 512730 272824 512736 272836
rect 512788 272824 512794 272876
rect 360712 272768 363000 272796
rect 360712 272756 360718 272768
rect 363230 272756 363236 272808
rect 363288 272796 363294 272808
rect 511534 272796 511540 272808
rect 363288 272768 511540 272796
rect 363288 272756 363294 272768
rect 511534 272756 511540 272768
rect 511592 272756 511598 272808
rect 511626 272756 511632 272808
rect 511684 272796 511690 272808
rect 610802 272796 610808 272808
rect 511684 272768 610808 272796
rect 511684 272756 511690 272768
rect 610802 272756 610808 272768
rect 610860 272756 610866 272808
rect 237282 272688 237288 272740
rect 237340 272728 237346 272740
rect 257154 272728 257160 272740
rect 237340 272700 257160 272728
rect 237340 272688 237346 272700
rect 257154 272688 257160 272700
rect 257212 272688 257218 272740
rect 296070 272688 296076 272740
rect 296128 272728 296134 272740
rect 341334 272728 341340 272740
rect 296128 272700 341340 272728
rect 296128 272688 296134 272700
rect 341334 272688 341340 272700
rect 341392 272688 341398 272740
rect 344922 272688 344928 272740
rect 344980 272728 344986 272740
rect 470134 272728 470140 272740
rect 344980 272700 362908 272728
rect 344980 272688 344986 272700
rect 300670 272620 300676 272672
rect 300728 272660 300734 272672
rect 351914 272660 351920 272672
rect 300728 272632 351920 272660
rect 300728 272620 300734 272632
rect 351914 272620 351920 272632
rect 351972 272620 351978 272672
rect 353018 272620 353024 272672
rect 353076 272660 353082 272672
rect 362770 272660 362776 272672
rect 353076 272632 362776 272660
rect 353076 272620 353082 272632
rect 362770 272620 362776 272632
rect 362828 272620 362834 272672
rect 362880 272660 362908 272700
rect 363064 272700 470140 272728
rect 363064 272660 363092 272700
rect 470134 272688 470140 272700
rect 470192 272688 470198 272740
rect 471974 272688 471980 272740
rect 472032 272728 472038 272740
rect 625062 272728 625068 272740
rect 472032 272700 625068 272728
rect 472032 272688 472038 272700
rect 625062 272688 625068 272700
rect 625120 272688 625126 272740
rect 362880 272632 363092 272660
rect 363138 272620 363144 272672
rect 363196 272660 363202 272672
rect 518618 272660 518624 272672
rect 363196 272632 518624 272660
rect 363196 272620 363202 272632
rect 518618 272620 518624 272632
rect 518676 272620 518682 272672
rect 232498 272552 232504 272604
rect 232556 272592 232562 272604
rect 255130 272592 255136 272604
rect 232556 272564 255136 272592
rect 232556 272552 232562 272564
rect 255130 272552 255136 272564
rect 255188 272552 255194 272604
rect 301406 272552 301412 272604
rect 301464 272592 301470 272604
rect 355502 272592 355508 272604
rect 301464 272564 355508 272592
rect 301464 272552 301470 272564
rect 355502 272552 355508 272564
rect 355560 272552 355566 272604
rect 368198 272552 368204 272604
rect 368256 272592 368262 272604
rect 532786 272592 532792 272604
rect 368256 272564 532792 272592
rect 368256 272552 368262 272564
rect 532786 272552 532792 272564
rect 532844 272552 532850 272604
rect 295242 272484 295248 272536
rect 295300 272524 295306 272536
rect 338942 272524 338948 272536
rect 295300 272496 338948 272524
rect 295300 272484 295306 272496
rect 338942 272484 338948 272496
rect 339000 272484 339006 272536
rect 342806 272484 342812 272536
rect 342864 272524 342870 272536
rect 465442 272524 465448 272536
rect 342864 272496 465448 272524
rect 342864 272484 342870 272496
rect 465442 272484 465448 272496
rect 465500 272484 465506 272536
rect 466270 272484 466276 272536
rect 466328 272524 466334 272536
rect 632146 272524 632152 272536
rect 466328 272496 632152 272524
rect 466328 272484 466334 272496
rect 632146 272484 632152 272496
rect 632204 272484 632210 272536
rect 230198 272416 230204 272468
rect 230256 272456 230262 272468
rect 254210 272456 254216 272468
rect 230256 272428 254216 272456
rect 230256 272416 230262 272428
rect 254210 272416 254216 272428
rect 254268 272416 254274 272468
rect 301866 272416 301872 272468
rect 301924 272456 301930 272468
rect 356698 272456 356704 272468
rect 301924 272428 356704 272456
rect 301924 272416 301930 272428
rect 356698 272416 356704 272428
rect 356756 272416 356762 272468
rect 360562 272416 360568 272468
rect 360620 272456 360626 272468
rect 363230 272456 363236 272468
rect 360620 272428 363236 272456
rect 360620 272416 360626 272428
rect 363230 272416 363236 272428
rect 363288 272416 363294 272468
rect 373166 272416 373172 272468
rect 373224 272456 373230 272468
rect 545850 272456 545856 272468
rect 373224 272428 545856 272456
rect 373224 272416 373230 272428
rect 545850 272416 545856 272428
rect 545908 272416 545914 272468
rect 303522 272348 303528 272400
rect 303580 272388 303586 272400
rect 360194 272388 360200 272400
rect 303580 272360 360200 272388
rect 303580 272348 303586 272360
rect 360194 272348 360200 272360
rect 360252 272348 360258 272400
rect 376662 272348 376668 272400
rect 376720 272388 376726 272400
rect 555234 272388 555240 272400
rect 376720 272360 555240 272388
rect 376720 272348 376726 272360
rect 555234 272348 555240 272360
rect 555292 272348 555298 272400
rect 295058 272280 295064 272332
rect 295116 272320 295122 272332
rect 331950 272320 331956 272332
rect 295116 272292 331956 272320
rect 295116 272280 295122 272292
rect 331950 272280 331956 272292
rect 332008 272280 332014 272332
rect 332502 272280 332508 272332
rect 332560 272320 332566 272332
rect 346026 272320 346032 272332
rect 332560 272292 346032 272320
rect 332560 272280 332566 272292
rect 346026 272280 346032 272292
rect 346084 272280 346090 272332
rect 351822 272280 351828 272332
rect 351880 272320 351886 272332
rect 458358 272320 458364 272332
rect 351880 272292 458364 272320
rect 351880 272280 351886 272292
rect 458358 272280 458364 272292
rect 458416 272280 458422 272332
rect 459462 272280 459468 272332
rect 459520 272320 459526 272332
rect 639230 272320 639236 272332
rect 459520 272292 639236 272320
rect 459520 272280 459526 272292
rect 639230 272280 639236 272292
rect 639288 272280 639294 272332
rect 227070 272252 227076 272264
rect 226306 272224 227076 272252
rect 227070 272212 227076 272224
rect 227128 272212 227134 272264
rect 303338 272212 303344 272264
rect 303396 272252 303402 272264
rect 358998 272252 359004 272264
rect 303396 272224 359004 272252
rect 303396 272212 303402 272224
rect 358998 272212 359004 272224
rect 359056 272212 359062 272264
rect 381998 272212 382004 272264
rect 382056 272252 382062 272264
rect 569494 272252 569500 272264
rect 382056 272224 569500 272252
rect 382056 272212 382062 272224
rect 569494 272212 569500 272224
rect 569552 272212 569558 272264
rect 93026 272144 93032 272196
rect 93084 272184 93090 272196
rect 184934 272184 184940 272196
rect 93084 272156 184940 272184
rect 93084 272144 93090 272156
rect 184934 272144 184940 272156
rect 184992 272144 184998 272196
rect 188798 272144 188804 272196
rect 188856 272184 188862 272196
rect 234798 272184 234804 272196
rect 188856 272156 234804 272184
rect 188856 272144 188862 272156
rect 234798 272144 234804 272156
rect 234856 272144 234862 272196
rect 238478 272144 238484 272196
rect 238536 272184 238542 272196
rect 257246 272184 257252 272196
rect 238536 272156 257252 272184
rect 238536 272144 238542 272156
rect 257246 272144 257252 272156
rect 257304 272144 257310 272196
rect 306282 272144 306288 272196
rect 306340 272184 306346 272196
rect 367278 272184 367284 272196
rect 306340 272156 367284 272184
rect 306340 272144 306346 272156
rect 367278 272144 367284 272156
rect 367336 272144 367342 272196
rect 384666 272144 384672 272196
rect 384724 272184 384730 272196
rect 576578 272184 576584 272196
rect 384724 272156 576584 272184
rect 384724 272144 384730 272156
rect 576578 272144 576584 272156
rect 576636 272144 576642 272196
rect 104894 272076 104900 272128
rect 104952 272116 104958 272128
rect 202690 272116 202696 272128
rect 104952 272088 202696 272116
rect 104952 272076 104958 272088
rect 202690 272076 202696 272088
rect 202748 272076 202754 272128
rect 205358 272076 205364 272128
rect 205416 272116 205422 272128
rect 240134 272116 240140 272128
rect 205416 272088 240140 272116
rect 205416 272076 205422 272088
rect 240134 272076 240140 272088
rect 240192 272076 240198 272128
rect 308950 272076 308956 272128
rect 309008 272116 309014 272128
rect 374362 272116 374368 272128
rect 309008 272088 374368 272116
rect 309008 272076 309014 272088
rect 374362 272076 374368 272088
rect 374420 272076 374426 272128
rect 387334 272076 387340 272128
rect 387392 272116 387398 272128
rect 583662 272116 583668 272128
rect 387392 272088 583668 272116
rect 387392 272076 387398 272088
rect 583662 272076 583668 272088
rect 583720 272076 583726 272128
rect 89530 272008 89536 272060
rect 89588 272048 89594 272060
rect 178034 272048 178040 272060
rect 89588 272020 178040 272048
rect 89588 272008 89594 272020
rect 178034 272008 178040 272020
rect 178092 272008 178098 272060
rect 178126 272008 178132 272060
rect 178184 272048 178190 272060
rect 197262 272048 197268 272060
rect 178184 272020 197268 272048
rect 178184 272008 178190 272020
rect 197262 272008 197268 272020
rect 197320 272008 197326 272060
rect 199470 272008 199476 272060
rect 199528 272048 199534 272060
rect 242618 272048 242624 272060
rect 199528 272020 242624 272048
rect 199528 272008 199534 272020
rect 242618 272008 242624 272020
rect 242676 272008 242682 272060
rect 284202 272008 284208 272060
rect 284260 272048 284266 272060
rect 309410 272048 309416 272060
rect 284260 272020 309416 272048
rect 284260 272008 284266 272020
rect 309410 272008 309416 272020
rect 309468 272008 309474 272060
rect 311618 272008 311624 272060
rect 311676 272048 311682 272060
rect 381538 272048 381544 272060
rect 311676 272020 381544 272048
rect 311676 272008 311682 272020
rect 381538 272008 381544 272020
rect 381596 272008 381602 272060
rect 394602 272008 394608 272060
rect 394660 272048 394666 272060
rect 590746 272048 590752 272060
rect 394660 272020 590752 272048
rect 394660 272008 394666 272020
rect 590746 272008 590752 272020
rect 590804 272008 590810 272060
rect 75270 271940 75276 271992
rect 75328 271980 75334 271992
rect 195422 271980 195428 271992
rect 75328 271952 195428 271980
rect 75328 271940 75334 271952
rect 195422 271940 195428 271952
rect 195480 271940 195486 271992
rect 201770 271940 201776 271992
rect 201828 271980 201834 271992
rect 243538 271980 243544 271992
rect 201828 271952 243544 271980
rect 201828 271940 201834 271952
rect 243538 271940 243544 271952
rect 243596 271940 243602 271992
rect 259546 271980 259552 271992
rect 245626 271952 259552 271980
rect 66990 271872 66996 271924
rect 67048 271912 67054 271924
rect 192478 271912 192484 271924
rect 67048 271884 192484 271912
rect 67048 271872 67054 271884
rect 192478 271872 192484 271884
rect 192536 271872 192542 271924
rect 242250 271912 242256 271924
rect 198706 271884 242256 271912
rect 65886 271804 65892 271856
rect 65944 271844 65950 271856
rect 192110 271844 192116 271856
rect 65944 271816 192116 271844
rect 65944 271804 65950 271816
rect 192110 271804 192116 271816
rect 192168 271804 192174 271856
rect 197170 271844 197176 271856
rect 194612 271816 197176 271844
rect 120258 271736 120264 271788
rect 120316 271776 120322 271788
rect 156782 271776 156788 271788
rect 120316 271748 156788 271776
rect 120316 271736 120322 271748
rect 156782 271736 156788 271748
rect 156840 271736 156846 271788
rect 156874 271736 156880 271788
rect 156932 271776 156938 271788
rect 177850 271776 177856 271788
rect 156932 271748 177856 271776
rect 156932 271736 156938 271748
rect 177850 271736 177856 271748
rect 177908 271736 177914 271788
rect 177942 271736 177948 271788
rect 178000 271776 178006 271788
rect 194502 271776 194508 271788
rect 178000 271748 194508 271776
rect 178000 271736 178006 271748
rect 194502 271736 194508 271748
rect 194560 271736 194566 271788
rect 130838 271668 130844 271720
rect 130896 271708 130902 271720
rect 194612 271708 194640 271816
rect 197170 271804 197176 271816
rect 197228 271804 197234 271856
rect 198274 271804 198280 271856
rect 198332 271844 198338 271856
rect 198706 271844 198734 271884
rect 242250 271872 242256 271884
rect 242308 271872 242314 271924
rect 240870 271844 240876 271856
rect 198332 271816 198734 271844
rect 208412 271816 240876 271844
rect 198332 271804 198338 271816
rect 130896 271680 194640 271708
rect 130896 271668 130902 271680
rect 194686 271668 194692 271720
rect 194744 271708 194750 271720
rect 208412 271708 208440 271816
rect 240870 271804 240876 271816
rect 240928 271804 240934 271856
rect 244366 271804 244372 271856
rect 244424 271844 244430 271856
rect 245626 271844 245654 271952
rect 259546 271940 259552 271952
rect 259604 271940 259610 271992
rect 285398 271940 285404 271992
rect 285456 271980 285462 271992
rect 312906 271980 312912 271992
rect 285456 271952 312912 271980
rect 285456 271940 285462 271952
rect 312906 271940 312912 271952
rect 312964 271940 312970 271992
rect 314286 271940 314292 271992
rect 314344 271980 314350 271992
rect 388622 271980 388628 271992
rect 314344 271952 388628 271980
rect 314344 271940 314350 271952
rect 388622 271940 388628 271952
rect 388680 271940 388686 271992
rect 395430 271940 395436 271992
rect 395488 271980 395494 271992
rect 604914 271980 604920 271992
rect 395488 271952 604920 271980
rect 395488 271940 395494 271952
rect 604914 271940 604920 271952
rect 604972 271940 604978 271992
rect 258718 271912 258724 271924
rect 244424 271816 245654 271844
rect 246500 271884 258724 271912
rect 244424 271804 244430 271816
rect 226518 271776 226524 271788
rect 226306 271748 226524 271776
rect 194744 271680 208440 271708
rect 194744 271668 194750 271680
rect 208486 271668 208492 271720
rect 208544 271708 208550 271720
rect 226306 271708 226334 271748
rect 226518 271736 226524 271748
rect 226576 271736 226582 271788
rect 241974 271736 241980 271788
rect 242032 271776 242038 271788
rect 246500 271776 246528 271884
rect 258718 271872 258724 271884
rect 258776 271872 258782 271924
rect 290274 271872 290280 271924
rect 290332 271912 290338 271924
rect 325970 271912 325976 271924
rect 290332 271884 325976 271912
rect 290332 271872 290338 271884
rect 325970 271872 325976 271884
rect 326028 271872 326034 271924
rect 326706 271872 326712 271924
rect 326764 271912 326770 271924
rect 402790 271912 402796 271924
rect 326764 271884 402796 271912
rect 326764 271872 326770 271884
rect 402790 271872 402796 271884
rect 402848 271872 402854 271924
rect 402882 271872 402888 271924
rect 402940 271912 402946 271924
rect 619082 271912 619088 271924
rect 402940 271884 619088 271912
rect 402940 271872 402946 271884
rect 619082 271872 619088 271884
rect 619140 271872 619146 271924
rect 258258 271844 258264 271856
rect 242032 271748 246528 271776
rect 246592 271816 258264 271844
rect 242032 271736 242038 271748
rect 208544 271680 226334 271708
rect 208544 271668 208550 271680
rect 240778 271668 240784 271720
rect 240836 271708 240842 271720
rect 246592 271708 246620 271816
rect 258258 271804 258264 271816
rect 258316 271804 258322 271856
rect 289538 271804 289544 271856
rect 289596 271844 289602 271856
rect 323578 271844 323584 271856
rect 289596 271816 323584 271844
rect 289596 271804 289602 271816
rect 323578 271804 323584 271816
rect 323636 271804 323642 271856
rect 325602 271804 325608 271856
rect 325660 271844 325666 271856
rect 409874 271844 409880 271856
rect 325660 271816 409880 271844
rect 325660 271804 325666 271816
rect 409874 271804 409880 271816
rect 409932 271804 409938 271856
rect 412818 271804 412824 271856
rect 412876 271844 412882 271856
rect 633342 271844 633348 271856
rect 412876 271816 633348 271844
rect 412876 271804 412882 271816
rect 633342 271804 633348 271816
rect 633400 271804 633406 271856
rect 255590 271776 255596 271788
rect 240836 271680 246620 271708
rect 246684 271748 255596 271776
rect 240836 271668 240842 271680
rect 163958 271600 163964 271652
rect 164016 271640 164022 271652
rect 229738 271640 229744 271652
rect 164016 271612 229744 271640
rect 164016 271600 164022 271612
rect 229738 271600 229744 271612
rect 229796 271600 229802 271652
rect 233694 271600 233700 271652
rect 233752 271640 233758 271652
rect 246684 271640 246712 271748
rect 255590 271736 255596 271748
rect 255648 271736 255654 271788
rect 262122 271736 262128 271788
rect 262180 271776 262186 271788
rect 266262 271776 266268 271788
rect 262180 271748 266268 271776
rect 262180 271736 262186 271748
rect 266262 271736 266268 271748
rect 266320 271736 266326 271788
rect 291746 271736 291752 271788
rect 291804 271776 291810 271788
rect 329466 271776 329472 271788
rect 291804 271748 329472 271776
rect 291804 271736 291810 271748
rect 329466 271736 329472 271748
rect 329524 271736 329530 271788
rect 340230 271736 340236 271788
rect 340288 271776 340294 271788
rect 351822 271776 351828 271788
rect 340288 271748 351828 271776
rect 340288 271736 340294 271748
rect 351822 271736 351828 271748
rect 351880 271736 351886 271788
rect 484302 271776 484308 271788
rect 351932 271748 484308 271776
rect 246758 271668 246764 271720
rect 246816 271708 246822 271720
rect 260466 271708 260472 271720
rect 246816 271680 260472 271708
rect 246816 271668 246822 271680
rect 260466 271668 260472 271680
rect 260524 271668 260530 271720
rect 290734 271668 290740 271720
rect 290792 271708 290798 271720
rect 327074 271708 327080 271720
rect 290792 271680 327080 271708
rect 290792 271668 290798 271680
rect 327074 271668 327080 271680
rect 327132 271668 327138 271720
rect 336734 271668 336740 271720
rect 336792 271708 336798 271720
rect 343634 271708 343640 271720
rect 336792 271680 343640 271708
rect 336792 271668 336798 271680
rect 343634 271668 343640 271680
rect 343692 271668 343698 271720
rect 233752 271612 246712 271640
rect 233752 271600 233758 271612
rect 247862 271600 247868 271652
rect 247920 271640 247926 271652
rect 260926 271640 260932 271652
rect 247920 271612 260932 271640
rect 247920 271600 247926 271612
rect 260926 271600 260932 271612
rect 260984 271600 260990 271652
rect 289814 271600 289820 271652
rect 289872 271640 289878 271652
rect 324774 271640 324780 271652
rect 289872 271612 324780 271640
rect 289872 271600 289878 271612
rect 324774 271600 324780 271612
rect 324832 271600 324838 271652
rect 350258 271600 350264 271652
rect 350316 271640 350322 271652
rect 351932 271640 351960 271748
rect 484302 271736 484308 271748
rect 484360 271736 484366 271788
rect 352374 271668 352380 271720
rect 352432 271708 352438 271720
rect 486694 271708 486700 271720
rect 352432 271680 486700 271708
rect 352432 271668 352438 271680
rect 486694 271668 486700 271680
rect 486752 271668 486758 271720
rect 479610 271640 479616 271652
rect 350316 271612 351960 271640
rect 352024 271612 479616 271640
rect 350316 271600 350322 271612
rect 165154 271532 165160 271584
rect 165212 271572 165218 271584
rect 229462 271572 229468 271584
rect 165212 271544 229468 271572
rect 165212 271532 165218 271544
rect 229462 271532 229468 271544
rect 229520 271532 229526 271584
rect 245562 271532 245568 271584
rect 245620 271572 245626 271584
rect 250162 271572 250168 271584
rect 245620 271544 250168 271572
rect 245620 271532 245626 271544
rect 250162 271532 250168 271544
rect 250220 271532 250226 271584
rect 250254 271532 250260 271584
rect 250312 271572 250318 271584
rect 261846 271572 261852 271584
rect 250312 271544 261852 271572
rect 250312 271532 250318 271544
rect 261846 271532 261852 271544
rect 261904 271532 261910 271584
rect 291194 271532 291200 271584
rect 291252 271572 291258 271584
rect 328270 271572 328276 271584
rect 291252 271544 328276 271572
rect 291252 271532 291258 271544
rect 328270 271532 328276 271544
rect 328328 271532 328334 271584
rect 348234 271532 348240 271584
rect 348292 271572 348298 271584
rect 352024 271572 352052 271612
rect 479610 271600 479616 271612
rect 479668 271600 479674 271652
rect 348292 271544 352052 271572
rect 348292 271532 348298 271544
rect 352098 271532 352104 271584
rect 352156 271572 352162 271584
rect 477218 271572 477224 271584
rect 352156 271544 477224 271572
rect 352156 271532 352162 271544
rect 477218 271532 477224 271544
rect 477276 271532 477282 271584
rect 158070 271464 158076 271516
rect 158128 271504 158134 271516
rect 177942 271504 177948 271516
rect 158128 271476 177948 271504
rect 158128 271464 158134 271476
rect 177942 271464 177948 271476
rect 178000 271464 178006 271516
rect 178126 271464 178132 271516
rect 178184 271504 178190 271516
rect 228818 271504 228824 271516
rect 178184 271476 228824 271504
rect 178184 271464 178190 271476
rect 228818 271464 228824 271476
rect 228876 271464 228882 271516
rect 231394 271464 231400 271516
rect 231452 271504 231458 271516
rect 254670 271504 254676 271516
rect 231452 271476 254676 271504
rect 231452 271464 231458 271476
rect 254670 271464 254676 271476
rect 254728 271464 254734 271516
rect 255038 271464 255044 271516
rect 255096 271504 255102 271516
rect 263594 271504 263600 271516
rect 255096 271476 263600 271504
rect 255096 271464 255102 271476
rect 263594 271464 263600 271476
rect 263652 271464 263658 271516
rect 289354 271464 289360 271516
rect 289412 271504 289418 271516
rect 322382 271504 322388 271516
rect 289412 271476 322388 271504
rect 289412 271464 289418 271476
rect 322382 271464 322388 271476
rect 322440 271464 322446 271516
rect 342162 271464 342168 271516
rect 342220 271504 342226 271516
rect 463050 271504 463056 271516
rect 342220 271476 352052 271504
rect 342220 271464 342226 271476
rect 171042 271396 171048 271448
rect 171100 271436 171106 271448
rect 232406 271436 232412 271448
rect 171100 271408 232412 271436
rect 171100 271396 171106 271408
rect 232406 271396 232412 271408
rect 232464 271396 232470 271448
rect 258534 271396 258540 271448
rect 258592 271436 258598 271448
rect 264882 271436 264888 271448
rect 258592 271408 264888 271436
rect 258592 271396 258598 271408
rect 264882 271396 264888 271408
rect 264940 271396 264946 271448
rect 288526 271396 288532 271448
rect 288584 271436 288590 271448
rect 321186 271436 321192 271448
rect 288584 271408 321192 271436
rect 288584 271396 288590 271408
rect 321186 271396 321192 271408
rect 321244 271396 321250 271448
rect 347590 271396 347596 271448
rect 347648 271436 347654 271448
rect 351914 271436 351920 271448
rect 347648 271408 351920 271436
rect 347648 271396 347654 271408
rect 351914 271396 351920 271408
rect 351972 271396 351978 271448
rect 352024 271436 352052 271476
rect 352300 271476 463056 271504
rect 352300 271436 352328 271476
rect 463050 271464 463056 271476
rect 463108 271464 463114 271516
rect 352024 271408 352328 271436
rect 355962 271396 355968 271448
rect 356020 271436 356026 271448
rect 472526 271436 472532 271448
rect 356020 271408 472532 271436
rect 356020 271396 356026 271408
rect 472526 271396 472532 271408
rect 472584 271396 472590 271448
rect 172238 271328 172244 271380
rect 172296 271368 172302 271380
rect 172296 271340 180012 271368
rect 172296 271328 172302 271340
rect 162762 271260 162768 271312
rect 162820 271300 162826 271312
rect 178126 271300 178132 271312
rect 162820 271272 178132 271300
rect 162820 271260 162826 271272
rect 178126 271260 178132 271272
rect 178184 271260 178190 271312
rect 179984 271300 180012 271340
rect 180058 271328 180064 271380
rect 180116 271368 180122 271380
rect 231486 271368 231492 271380
rect 180116 271340 231492 271368
rect 180116 271328 180122 271340
rect 231486 271328 231492 271340
rect 231544 271328 231550 271380
rect 257338 271328 257344 271380
rect 257396 271368 257402 271380
rect 264514 271368 264520 271380
rect 257396 271340 264520 271368
rect 257396 271328 257402 271340
rect 264514 271328 264520 271340
rect 264572 271328 264578 271380
rect 287606 271328 287612 271380
rect 287664 271368 287670 271380
rect 318794 271368 318800 271380
rect 287664 271340 318800 271368
rect 287664 271328 287670 271340
rect 318794 271328 318800 271340
rect 318852 271328 318858 271380
rect 339402 271328 339408 271380
rect 339460 271368 339466 271380
rect 455966 271368 455972 271380
rect 339460 271340 455972 271368
rect 339460 271328 339466 271340
rect 455966 271328 455972 271340
rect 456024 271328 456030 271380
rect 231762 271300 231768 271312
rect 179984 271272 231768 271300
rect 231762 271260 231768 271272
rect 231820 271260 231826 271312
rect 256142 271260 256148 271312
rect 256200 271300 256206 271312
rect 264054 271300 264060 271312
rect 256200 271272 264060 271300
rect 256200 271260 256206 271272
rect 264054 271260 264060 271272
rect 264112 271260 264118 271312
rect 286778 271260 286784 271312
rect 286836 271300 286842 271312
rect 316494 271300 316500 271312
rect 286836 271272 316500 271300
rect 286836 271260 286842 271272
rect 316494 271260 316500 271272
rect 316552 271260 316558 271312
rect 336458 271260 336464 271312
rect 336516 271300 336522 271312
rect 448882 271300 448888 271312
rect 336516 271272 448888 271300
rect 336516 271260 336522 271272
rect 448882 271260 448888 271272
rect 448940 271260 448946 271312
rect 178034 271192 178040 271244
rect 178092 271232 178098 271244
rect 188614 271232 188620 271244
rect 178092 271204 188620 271232
rect 178092 271192 178098 271204
rect 188614 271192 188620 271204
rect 188672 271192 188678 271244
rect 197262 271192 197268 271244
rect 197320 271232 197326 271244
rect 231946 271232 231952 271244
rect 197320 271204 231952 271232
rect 197320 271192 197326 271204
rect 231946 271192 231952 271204
rect 232004 271192 232010 271244
rect 251450 271192 251456 271244
rect 251508 271232 251514 271244
rect 262214 271232 262220 271244
rect 251508 271204 262220 271232
rect 251508 271192 251514 271204
rect 262214 271192 262220 271204
rect 262272 271192 262278 271244
rect 288158 271192 288164 271244
rect 288216 271232 288222 271244
rect 319990 271232 319996 271244
rect 288216 271204 319996 271232
rect 288216 271192 288222 271204
rect 319990 271192 319996 271204
rect 320048 271192 320054 271244
rect 337470 271192 337476 271244
rect 337528 271232 337534 271244
rect 451274 271232 451280 271244
rect 337528 271204 451280 271232
rect 337528 271192 337534 271204
rect 451274 271192 451280 271204
rect 451332 271192 451338 271244
rect 179322 271124 179328 271176
rect 179380 271164 179386 271176
rect 234522 271164 234528 271176
rect 179380 271136 234528 271164
rect 179380 271124 179386 271136
rect 234522 271124 234528 271136
rect 234580 271124 234586 271176
rect 249058 271124 249064 271176
rect 249116 271164 249122 271176
rect 261386 271164 261392 271176
rect 249116 271136 261392 271164
rect 249116 271124 249122 271136
rect 261386 271124 261392 271136
rect 261444 271124 261450 271176
rect 287146 271124 287152 271176
rect 287204 271164 287210 271176
rect 317690 271164 317696 271176
rect 287204 271136 317696 271164
rect 287204 271124 287210 271136
rect 317690 271124 317696 271136
rect 317748 271124 317754 271176
rect 333974 271124 333980 271176
rect 334032 271164 334038 271176
rect 441798 271164 441804 271176
rect 334032 271136 441804 271164
rect 334032 271124 334038 271136
rect 441798 271124 441804 271136
rect 441856 271124 441862 271176
rect 169846 271056 169852 271108
rect 169904 271096 169910 271108
rect 180058 271096 180064 271108
rect 169904 271068 180064 271096
rect 169904 271056 169910 271068
rect 180058 271056 180064 271068
rect 180116 271056 180122 271108
rect 182910 271056 182916 271108
rect 182968 271096 182974 271108
rect 232038 271096 232044 271108
rect 182968 271068 232044 271096
rect 182968 271056 182974 271068
rect 232038 271056 232044 271068
rect 232096 271056 232102 271108
rect 253842 271056 253848 271108
rect 253900 271096 253906 271108
rect 263134 271096 263140 271108
rect 253900 271068 263140 271096
rect 253900 271056 253906 271068
rect 263134 271056 263140 271068
rect 263192 271056 263198 271108
rect 266814 271056 266820 271108
rect 266872 271096 266878 271108
rect 268010 271096 268016 271108
rect 266872 271068 268016 271096
rect 266872 271056 266878 271068
rect 268010 271056 268016 271068
rect 268068 271056 268074 271108
rect 286686 271056 286692 271108
rect 286744 271096 286750 271108
rect 315298 271096 315304 271108
rect 286744 271068 315304 271096
rect 286744 271056 286750 271068
rect 315298 271056 315304 271068
rect 315356 271056 315362 271108
rect 334802 271056 334808 271108
rect 334860 271096 334866 271108
rect 444190 271096 444196 271108
rect 334860 271068 444196 271096
rect 334860 271056 334866 271068
rect 444190 271056 444196 271068
rect 444248 271056 444254 271108
rect 176930 270988 176936 271040
rect 176988 271028 176994 271040
rect 226426 271028 226432 271040
rect 176988 271000 226432 271028
rect 176988 270988 176994 271000
rect 226426 270988 226432 271000
rect 226484 270988 226490 271040
rect 226610 270988 226616 271040
rect 226668 271028 226674 271040
rect 252922 271028 252928 271040
rect 226668 271000 252928 271028
rect 226668 270988 226674 271000
rect 252922 270988 252928 271000
rect 252980 270988 252986 271040
rect 331306 270988 331312 271040
rect 331364 271028 331370 271040
rect 434714 271028 434720 271040
rect 331364 271000 434720 271028
rect 331364 270988 331370 271000
rect 434714 270988 434720 271000
rect 434772 270988 434778 271040
rect 175826 270920 175832 270972
rect 175884 270960 175890 270972
rect 179322 270960 179328 270972
rect 175884 270932 179328 270960
rect 175884 270920 175890 270932
rect 179322 270920 179328 270932
rect 179380 270920 179386 270972
rect 185210 270920 185216 270972
rect 185268 270960 185274 270972
rect 234706 270960 234712 270972
rect 185268 270932 234712 270960
rect 185268 270920 185274 270932
rect 234706 270920 234712 270932
rect 234764 270920 234770 270972
rect 250162 270920 250168 270972
rect 250220 270960 250226 270972
rect 260006 270960 260012 270972
rect 250220 270932 260012 270960
rect 250220 270920 250226 270932
rect 260006 270920 260012 270932
rect 260064 270920 260070 270972
rect 285858 270920 285864 270972
rect 285916 270960 285922 270972
rect 314102 270960 314108 270972
rect 285916 270932 314108 270960
rect 285916 270920 285922 270932
rect 314102 270920 314108 270932
rect 314160 270920 314166 270972
rect 329926 270920 329932 270972
rect 329984 270960 329990 270972
rect 431126 270960 431132 270972
rect 329984 270932 431132 270960
rect 329984 270920 329990 270932
rect 431126 270920 431132 270932
rect 431184 270920 431190 270972
rect 186406 270852 186412 270904
rect 186464 270892 186470 270904
rect 232130 270892 232136 270904
rect 186464 270864 232136 270892
rect 186464 270852 186470 270864
rect 232130 270852 232136 270864
rect 232188 270852 232194 270904
rect 327258 270852 327264 270904
rect 327316 270892 327322 270904
rect 424042 270892 424048 270904
rect 327316 270864 424048 270892
rect 327316 270852 327322 270864
rect 424042 270852 424048 270864
rect 424100 270852 424106 270904
rect 189994 270784 190000 270836
rect 190052 270824 190058 270836
rect 232498 270824 232504 270836
rect 190052 270796 232504 270824
rect 190052 270784 190058 270796
rect 232498 270784 232504 270796
rect 232556 270784 232562 270836
rect 259730 270784 259736 270836
rect 259788 270824 259794 270836
rect 265342 270824 265348 270836
rect 259788 270796 265348 270824
rect 259788 270784 259794 270796
rect 265342 270784 265348 270796
rect 265400 270784 265406 270836
rect 329006 270784 329012 270836
rect 329064 270824 329070 270836
rect 340138 270824 340144 270836
rect 329064 270796 340144 270824
rect 329064 270784 329070 270796
rect 340138 270784 340144 270796
rect 340196 270784 340202 270836
rect 340322 270784 340328 270836
rect 340380 270824 340386 270836
rect 416958 270824 416964 270836
rect 340380 270796 416964 270824
rect 340380 270784 340386 270796
rect 416958 270784 416964 270796
rect 417016 270784 417022 270836
rect 187602 270716 187608 270768
rect 187660 270756 187666 270768
rect 202782 270756 202788 270768
rect 187660 270728 202788 270756
rect 187660 270716 187666 270728
rect 202782 270716 202788 270728
rect 202840 270716 202846 270768
rect 206738 270716 206744 270768
rect 206796 270756 206802 270768
rect 229370 270756 229376 270768
rect 206796 270728 229376 270756
rect 206796 270716 206802 270728
rect 229370 270716 229376 270728
rect 229428 270716 229434 270768
rect 326430 270716 326436 270768
rect 326488 270756 326494 270768
rect 395706 270756 395712 270768
rect 326488 270728 395712 270756
rect 326488 270716 326494 270728
rect 395706 270716 395712 270728
rect 395764 270716 395770 270768
rect 191190 270648 191196 270700
rect 191248 270688 191254 270700
rect 230198 270688 230204 270700
rect 191248 270660 193214 270688
rect 191248 270648 191254 270660
rect 193186 270620 193214 270660
rect 212506 270660 230204 270688
rect 206738 270620 206744 270632
rect 193186 270592 206744 270620
rect 206738 270580 206744 270592
rect 206796 270580 206802 270632
rect 192294 270512 192300 270564
rect 192352 270552 192358 270564
rect 198642 270552 198648 270564
rect 192352 270524 198648 270552
rect 192352 270512 192358 270524
rect 198642 270512 198648 270524
rect 198700 270512 198706 270564
rect 202782 270512 202788 270564
rect 202840 270552 202846 270564
rect 212506 270552 212534 270660
rect 230198 270648 230204 270660
rect 230256 270648 230262 270700
rect 252646 270648 252652 270700
rect 252704 270688 252710 270700
rect 262858 270688 262864 270700
rect 252704 270660 262864 270688
rect 252704 270648 252710 270660
rect 262858 270648 262864 270660
rect 262916 270648 262922 270700
rect 331122 270648 331128 270700
rect 331180 270688 331186 270700
rect 377950 270688 377956 270700
rect 331180 270660 377956 270688
rect 331180 270648 331186 270660
rect 377950 270648 377956 270660
rect 378008 270648 378014 270700
rect 229002 270580 229008 270632
rect 229060 270620 229066 270632
rect 253750 270620 253756 270632
rect 229060 270592 253756 270620
rect 229060 270580 229066 270592
rect 253750 270580 253756 270592
rect 253808 270580 253814 270632
rect 324590 270580 324596 270632
rect 324648 270620 324654 270632
rect 340322 270620 340328 270632
rect 324648 270592 340328 270620
rect 324648 270580 324654 270592
rect 340322 270580 340328 270592
rect 340380 270580 340386 270632
rect 352006 270580 352012 270632
rect 352064 270620 352070 270632
rect 394510 270620 394516 270632
rect 352064 270592 394516 270620
rect 352064 270580 352070 270592
rect 394510 270580 394516 270592
rect 394568 270580 394574 270632
rect 202840 270524 212534 270552
rect 202840 270512 202846 270524
rect 227806 270512 227812 270564
rect 227864 270552 227870 270564
rect 253382 270552 253388 270564
rect 227864 270524 253388 270552
rect 227864 270512 227870 270524
rect 253382 270512 253388 270524
rect 253440 270512 253446 270564
rect 357434 270512 357440 270564
rect 357492 270552 357498 270564
rect 385034 270552 385040 270564
rect 357492 270524 385040 270552
rect 357492 270512 357498 270524
rect 385034 270512 385040 270524
rect 385092 270512 385098 270564
rect 411806 270512 411812 270564
rect 411864 270552 411870 270564
rect 413094 270552 413100 270564
rect 411864 270524 413100 270552
rect 411864 270512 411870 270524
rect 413094 270512 413100 270524
rect 413152 270512 413158 270564
rect 154482 270444 154488 270496
rect 154540 270484 154546 270496
rect 206462 270484 206468 270496
rect 154540 270456 206468 270484
rect 154540 270444 154546 270456
rect 206462 270444 206468 270456
rect 206520 270444 206526 270496
rect 222654 270484 222660 270496
rect 206572 270456 222660 270484
rect 147398 270376 147404 270428
rect 147456 270416 147462 270428
rect 206572 270416 206600 270456
rect 222654 270444 222660 270456
rect 222712 270444 222718 270496
rect 225414 270444 225420 270496
rect 225472 270484 225478 270496
rect 252462 270484 252468 270496
rect 225472 270456 252468 270484
rect 225472 270444 225478 270456
rect 252462 270444 252468 270456
rect 252520 270444 252526 270496
rect 265618 270444 265624 270496
rect 265676 270484 265682 270496
rect 267550 270484 267556 270496
rect 265676 270456 267556 270484
rect 265676 270444 265682 270456
rect 267550 270444 267556 270456
rect 267608 270444 267614 270496
rect 269850 270444 269856 270496
rect 269908 270484 269914 270496
rect 271506 270484 271512 270496
rect 269908 270456 271512 270484
rect 269908 270444 269914 270456
rect 271506 270444 271512 270456
rect 271564 270444 271570 270496
rect 272058 270444 272064 270496
rect 272116 270484 272122 270496
rect 277486 270484 277492 270496
rect 272116 270456 277492 270484
rect 272116 270444 272122 270456
rect 277486 270444 277492 270456
rect 277544 270444 277550 270496
rect 304074 270444 304080 270496
rect 304132 270484 304138 270496
rect 344002 270484 344008 270496
rect 304132 270456 344008 270484
rect 304132 270444 304138 270456
rect 344002 270444 344008 270456
rect 344060 270444 344066 270496
rect 346854 270444 346860 270496
rect 346912 270484 346918 270496
rect 476114 270484 476120 270496
rect 346912 270456 476120 270484
rect 346912 270444 346918 270456
rect 476114 270444 476120 270456
rect 476172 270444 476178 270496
rect 220814 270416 220820 270428
rect 147456 270388 206600 270416
rect 208228 270388 220820 270416
rect 147456 270376 147462 270388
rect 140314 270308 140320 270360
rect 140372 270348 140378 270360
rect 208026 270348 208032 270360
rect 140372 270320 208032 270348
rect 140372 270308 140378 270320
rect 208026 270308 208032 270320
rect 208084 270308 208090 270360
rect 141510 270240 141516 270292
rect 141568 270280 141574 270292
rect 208228 270280 208256 270388
rect 220814 270376 220820 270388
rect 220872 270376 220878 270428
rect 224218 270376 224224 270428
rect 224276 270416 224282 270428
rect 252002 270416 252008 270428
rect 224276 270388 252008 270416
rect 224276 270376 224282 270388
rect 252002 270376 252008 270388
rect 252060 270376 252066 270428
rect 270310 270376 270316 270428
rect 270368 270416 270374 270428
rect 272702 270416 272708 270428
rect 270368 270388 272708 270416
rect 270368 270376 270374 270388
rect 272702 270376 272708 270388
rect 272760 270376 272766 270428
rect 272978 270376 272984 270428
rect 273036 270416 273042 270428
rect 279786 270416 279792 270428
rect 273036 270388 279792 270416
rect 273036 270376 273042 270388
rect 279786 270376 279792 270388
rect 279844 270376 279850 270428
rect 294322 270376 294328 270428
rect 294380 270416 294386 270428
rect 336550 270416 336556 270428
rect 294380 270388 336556 270416
rect 294380 270376 294386 270388
rect 336550 270376 336556 270388
rect 336608 270376 336614 270428
rect 348602 270376 348608 270428
rect 348660 270416 348666 270428
rect 480806 270416 480812 270428
rect 348660 270388 480812 270416
rect 348660 270376 348666 270388
rect 480806 270376 480812 270388
rect 480864 270376 480870 270428
rect 208302 270308 208308 270360
rect 208360 270348 208366 270360
rect 219986 270348 219992 270360
rect 208360 270320 219992 270348
rect 208360 270308 208366 270320
rect 219986 270308 219992 270320
rect 220044 270308 220050 270360
rect 220722 270308 220728 270360
rect 220780 270348 220786 270360
rect 250714 270348 250720 270360
rect 220780 270320 250720 270348
rect 220780 270308 220786 270320
rect 250714 270308 250720 270320
rect 250772 270308 250778 270360
rect 270678 270308 270684 270360
rect 270736 270348 270742 270360
rect 273898 270348 273904 270360
rect 270736 270320 273904 270348
rect 270736 270308 270742 270320
rect 273898 270308 273904 270320
rect 273956 270308 273962 270360
rect 274266 270308 274272 270360
rect 274324 270348 274330 270360
rect 283374 270348 283380 270360
rect 274324 270320 283380 270348
rect 274324 270308 274330 270320
rect 283374 270308 283380 270320
rect 283432 270308 283438 270360
rect 296990 270308 296996 270360
rect 297048 270348 297054 270360
rect 336734 270348 336740 270360
rect 297048 270320 336740 270348
rect 297048 270308 297054 270320
rect 336734 270308 336740 270320
rect 336792 270308 336798 270360
rect 349522 270308 349528 270360
rect 349580 270348 349586 270360
rect 483198 270348 483204 270360
rect 349580 270320 483204 270348
rect 349580 270308 349586 270320
rect 483198 270308 483204 270320
rect 483256 270308 483262 270360
rect 219066 270280 219072 270292
rect 141568 270252 208256 270280
rect 208320 270252 219072 270280
rect 141568 270240 141574 270252
rect 135622 270172 135628 270224
rect 135680 270212 135686 270224
rect 208320 270212 208348 270252
rect 219066 270240 219072 270252
rect 219124 270240 219130 270292
rect 221918 270240 221924 270292
rect 221976 270280 221982 270292
rect 251082 270280 251088 270292
rect 221976 270252 251088 270280
rect 221976 270240 221982 270252
rect 251082 270240 251088 270252
rect 251140 270240 251146 270292
rect 271138 270240 271144 270292
rect 271196 270280 271202 270292
rect 275094 270280 275100 270292
rect 271196 270252 275100 270280
rect 271196 270240 271202 270252
rect 275094 270240 275100 270252
rect 275152 270240 275158 270292
rect 277394 270240 277400 270292
rect 277452 270280 277458 270292
rect 291654 270280 291660 270292
rect 277452 270252 291660 270280
rect 277452 270240 277458 270252
rect 291654 270240 291660 270252
rect 291712 270240 291718 270292
rect 297450 270240 297456 270292
rect 297508 270280 297514 270292
rect 339494 270280 339500 270292
rect 297508 270252 339500 270280
rect 297508 270240 297514 270252
rect 339494 270240 339500 270252
rect 339552 270240 339558 270292
rect 351270 270240 351276 270292
rect 351328 270280 351334 270292
rect 487890 270280 487896 270292
rect 351328 270252 487896 270280
rect 351328 270240 351334 270252
rect 487890 270240 487896 270252
rect 487948 270240 487954 270292
rect 135680 270184 208348 270212
rect 135680 270172 135686 270184
rect 208394 270172 208400 270224
rect 208452 270212 208458 270224
rect 218146 270212 218152 270224
rect 208452 270184 218152 270212
rect 208452 270172 208458 270184
rect 218146 270172 218152 270184
rect 218204 270172 218210 270224
rect 218330 270172 218336 270224
rect 218388 270212 218394 270224
rect 249794 270212 249800 270224
rect 218388 270184 249800 270212
rect 218388 270172 218394 270184
rect 249794 270172 249800 270184
rect 249852 270172 249858 270224
rect 272518 270172 272524 270224
rect 272576 270212 272582 270224
rect 278682 270212 278688 270224
rect 272576 270184 278688 270212
rect 272576 270172 272582 270184
rect 278682 270172 278688 270184
rect 278740 270172 278746 270224
rect 278774 270172 278780 270224
rect 278832 270212 278838 270224
rect 290458 270212 290464 270224
rect 278832 270184 290464 270212
rect 278832 270172 278838 270184
rect 290458 270172 290464 270184
rect 290516 270172 290522 270224
rect 296530 270172 296536 270224
rect 296588 270212 296594 270224
rect 342438 270212 342444 270224
rect 296588 270184 342444 270212
rect 296588 270172 296594 270184
rect 342438 270172 342444 270184
rect 342496 270172 342502 270224
rect 352190 270172 352196 270224
rect 352248 270212 352254 270224
rect 490282 270212 490288 270224
rect 352248 270184 490288 270212
rect 352248 270172 352254 270184
rect 490282 270172 490288 270184
rect 490340 270172 490346 270224
rect 133230 270104 133236 270156
rect 133288 270144 133294 270156
rect 133288 270116 215892 270144
rect 133288 270104 133294 270116
rect 134426 270036 134432 270088
rect 134484 270076 134490 270088
rect 208210 270076 208216 270088
rect 134484 270048 208216 270076
rect 134484 270036 134490 270048
rect 208210 270036 208216 270048
rect 208268 270036 208274 270088
rect 215864 270076 215892 270116
rect 215938 270104 215944 270156
rect 215996 270144 216002 270156
rect 248874 270144 248880 270156
rect 215996 270116 248880 270144
rect 215996 270104 216002 270116
rect 248874 270104 248880 270116
rect 248932 270104 248938 270156
rect 273714 270104 273720 270156
rect 273772 270144 273778 270156
rect 280982 270144 280988 270156
rect 273772 270116 280988 270144
rect 273772 270104 273778 270116
rect 280982 270104 280988 270116
rect 281040 270104 281046 270156
rect 295150 270144 295156 270156
rect 281276 270116 295156 270144
rect 217318 270076 217324 270088
rect 215864 270048 217324 270076
rect 217318 270036 217324 270048
rect 217376 270036 217382 270088
rect 223114 270036 223120 270088
rect 223172 270076 223178 270088
rect 251542 270076 251548 270088
rect 223172 270048 251548 270076
rect 223172 270036 223178 270048
rect 251542 270036 251548 270048
rect 251600 270036 251606 270088
rect 271598 270036 271604 270088
rect 271656 270076 271662 270088
rect 276290 270076 276296 270088
rect 271656 270048 276296 270076
rect 271656 270036 271662 270048
rect 276290 270036 276296 270048
rect 276348 270036 276354 270088
rect 278682 270036 278688 270088
rect 278740 270076 278746 270088
rect 281276 270076 281304 270116
rect 295150 270104 295156 270116
rect 295208 270104 295214 270156
rect 298278 270104 298284 270156
rect 298336 270144 298342 270156
rect 347222 270144 347228 270156
rect 298336 270116 347228 270144
rect 298336 270104 298342 270116
rect 347222 270104 347228 270116
rect 347280 270104 347286 270156
rect 350902 270104 350908 270156
rect 350960 270144 350966 270156
rect 352374 270144 352380 270156
rect 350960 270116 352380 270144
rect 350960 270104 350966 270116
rect 352374 270104 352380 270116
rect 352432 270104 352438 270156
rect 353570 270104 353576 270156
rect 353628 270144 353634 270156
rect 493778 270144 493784 270156
rect 353628 270116 493784 270144
rect 353628 270104 353634 270116
rect 493778 270104 493784 270116
rect 493836 270104 493842 270156
rect 294046 270076 294052 270088
rect 278740 270048 281304 270076
rect 281368 270048 294052 270076
rect 278740 270036 278746 270048
rect 126146 269968 126152 270020
rect 126204 270008 126210 270020
rect 126204 269980 213592 270008
rect 126204 269968 126210 269980
rect 119062 269900 119068 269952
rect 119120 269940 119126 269952
rect 211890 269940 211896 269952
rect 119120 269912 211896 269940
rect 119120 269900 119126 269912
rect 211890 269900 211896 269912
rect 211948 269900 211954 269952
rect 213564 269940 213592 269980
rect 213638 269968 213644 270020
rect 213696 270008 213702 270020
rect 248046 270008 248052 270020
rect 213696 269980 248052 270008
rect 213696 269968 213702 269980
rect 248046 269968 248052 269980
rect 248104 269968 248110 270020
rect 278314 269968 278320 270020
rect 278372 270008 278378 270020
rect 281368 270008 281396 270048
rect 294046 270036 294052 270048
rect 294104 270036 294110 270088
rect 299198 270036 299204 270088
rect 299256 270076 299262 270088
rect 349614 270076 349620 270088
rect 299256 270048 349620 270076
rect 299256 270036 299262 270048
rect 349614 270036 349620 270048
rect 349672 270036 349678 270088
rect 355962 270076 355968 270088
rect 349724 270048 355968 270076
rect 278372 269980 281396 270008
rect 278372 269968 278378 269980
rect 281534 269968 281540 270020
rect 281592 270008 281598 270020
rect 292850 270008 292856 270020
rect 281592 269980 292856 270008
rect 281592 269968 281598 269980
rect 292850 269968 292856 269980
rect 292908 269968 292914 270020
rect 345474 269968 345480 270020
rect 345532 270008 345538 270020
rect 349724 270008 349752 270048
rect 355962 270036 355968 270048
rect 356020 270036 356026 270088
rect 356238 270036 356244 270088
rect 356296 270076 356302 270088
rect 500862 270076 500868 270088
rect 356296 270048 500868 270076
rect 356296 270036 356302 270048
rect 500862 270036 500868 270048
rect 500920 270036 500926 270088
rect 345532 269980 349752 270008
rect 345532 269968 345538 269980
rect 351730 269968 351736 270020
rect 351788 270008 351794 270020
rect 363782 270008 363788 270020
rect 351788 269980 363788 270008
rect 351788 269968 351794 269980
rect 363782 269968 363788 269980
rect 363840 269968 363846 270020
rect 364702 269968 364708 270020
rect 364760 270008 364766 270020
rect 364760 269980 382412 270008
rect 364760 269968 364766 269980
rect 214650 269940 214656 269952
rect 213564 269912 214656 269940
rect 214650 269900 214656 269912
rect 214708 269900 214714 269952
rect 217134 269900 217140 269952
rect 217192 269940 217198 269952
rect 249334 269940 249340 269952
rect 217192 269912 249340 269940
rect 217192 269900 217198 269912
rect 249334 269900 249340 269912
rect 249392 269900 249398 269952
rect 276934 269900 276940 269952
rect 276992 269940 276998 269952
rect 278774 269940 278780 269952
rect 276992 269912 278780 269940
rect 276992 269900 276998 269912
rect 278774 269900 278780 269912
rect 278832 269900 278838 269952
rect 279602 269900 279608 269952
rect 279660 269940 279666 269952
rect 297542 269940 297548 269952
rect 279660 269912 297548 269940
rect 279660 269900 279666 269912
rect 297542 269900 297548 269912
rect 297600 269900 297606 269952
rect 305454 269900 305460 269952
rect 305512 269940 305518 269952
rect 366082 269940 366088 269952
rect 305512 269912 366088 269940
rect 305512 269900 305518 269912
rect 366082 269900 366088 269912
rect 366140 269900 366146 269952
rect 367370 269900 367376 269952
rect 367428 269940 367434 269952
rect 382384 269940 382412 269980
rect 382458 269968 382464 270020
rect 382516 270008 382522 270020
rect 515122 270008 515128 270020
rect 382516 269980 515128 270008
rect 382516 269968 382522 269980
rect 515122 269968 515128 269980
rect 515180 269968 515186 270020
rect 523402 269940 523408 269952
rect 367428 269912 382136 269940
rect 382384 269912 523408 269940
rect 367428 269900 367434 269912
rect 110782 269832 110788 269884
rect 110840 269872 110846 269884
rect 209682 269872 209688 269884
rect 110840 269844 209688 269872
rect 110840 269832 110846 269844
rect 209682 269832 209688 269844
rect 209740 269832 209746 269884
rect 210050 269832 210056 269884
rect 210108 269872 210114 269884
rect 246666 269872 246672 269884
rect 210108 269844 246672 269872
rect 210108 269832 210114 269844
rect 246666 269832 246672 269844
rect 246724 269832 246730 269884
rect 279142 269832 279148 269884
rect 279200 269872 279206 269884
rect 296346 269872 296352 269884
rect 279200 269844 296352 269872
rect 279200 269832 279206 269844
rect 296346 269832 296352 269844
rect 296404 269832 296410 269884
rect 306742 269832 306748 269884
rect 306800 269872 306806 269884
rect 369670 269872 369676 269884
rect 306800 269844 369676 269872
rect 306800 269832 306806 269844
rect 369670 269832 369676 269844
rect 369728 269832 369734 269884
rect 370038 269832 370044 269884
rect 370096 269872 370102 269884
rect 382108 269872 382136 269912
rect 523402 269900 523408 269912
rect 523460 269900 523466 269952
rect 530486 269872 530492 269884
rect 370096 269844 382044 269872
rect 382108 269844 530492 269872
rect 370096 269832 370102 269844
rect 114278 269764 114284 269816
rect 114336 269804 114342 269816
rect 211062 269804 211068 269816
rect 114336 269776 211068 269804
rect 114336 269764 114342 269776
rect 211062 269764 211068 269776
rect 211120 269764 211126 269816
rect 214834 269764 214840 269816
rect 214892 269804 214898 269816
rect 248414 269804 248420 269816
rect 214892 269776 248420 269804
rect 214892 269764 214898 269776
rect 248414 269764 248420 269776
rect 248472 269764 248478 269816
rect 280522 269764 280528 269816
rect 280580 269804 280586 269816
rect 299934 269804 299940 269816
rect 280580 269776 299940 269804
rect 280580 269764 280586 269776
rect 299934 269764 299940 269776
rect 299992 269764 299998 269816
rect 307202 269764 307208 269816
rect 307260 269804 307266 269816
rect 370866 269804 370872 269816
rect 307260 269776 370872 269804
rect 307260 269764 307266 269776
rect 370866 269764 370872 269776
rect 370924 269764 370930 269816
rect 373258 269804 373264 269816
rect 372586 269776 373264 269804
rect 109586 269696 109592 269748
rect 109644 269736 109650 269748
rect 208854 269736 208860 269748
rect 109644 269708 208860 269736
rect 109644 269696 109650 269708
rect 208854 269696 208860 269708
rect 208912 269696 208918 269748
rect 212442 269696 212448 269748
rect 212500 269736 212506 269748
rect 247586 269736 247592 269748
rect 212500 269708 247592 269736
rect 212500 269696 212506 269708
rect 247586 269696 247592 269708
rect 247644 269696 247650 269748
rect 280062 269696 280068 269748
rect 280120 269736 280126 269748
rect 298738 269736 298744 269748
rect 280120 269708 298744 269736
rect 280120 269696 280126 269708
rect 298738 269696 298744 269708
rect 298796 269696 298802 269748
rect 308122 269696 308128 269748
rect 308180 269736 308186 269748
rect 372586 269736 372614 269776
rect 373258 269764 373264 269776
rect 373316 269764 373322 269816
rect 382016 269804 382044 269844
rect 530486 269832 530492 269844
rect 530544 269832 530550 269884
rect 537570 269804 537576 269816
rect 382016 269776 537576 269804
rect 537570 269764 537576 269776
rect 537628 269764 537634 269816
rect 308180 269708 372614 269736
rect 308180 269696 308186 269708
rect 375374 269696 375380 269748
rect 375432 269736 375438 269748
rect 375432 269708 382412 269736
rect 375432 269696 375438 269708
rect 102502 269628 102508 269680
rect 102560 269668 102566 269680
rect 206186 269668 206192 269680
rect 102560 269640 206192 269668
rect 102560 269628 102566 269640
rect 206186 269628 206192 269640
rect 206244 269628 206250 269680
rect 209130 269628 209136 269680
rect 209188 269668 209194 269680
rect 246206 269668 246212 269680
rect 209188 269640 246212 269668
rect 209188 269628 209194 269640
rect 246206 269628 246212 269640
rect 246264 269628 246270 269680
rect 277854 269628 277860 269680
rect 277912 269668 277918 269680
rect 281534 269668 281540 269680
rect 277912 269640 281540 269668
rect 277912 269628 277918 269640
rect 281534 269628 281540 269640
rect 281592 269628 281598 269680
rect 281810 269628 281816 269680
rect 281868 269668 281874 269680
rect 303430 269668 303436 269680
rect 281868 269640 303436 269668
rect 281868 269628 281874 269640
rect 303430 269628 303436 269640
rect 303488 269628 303494 269680
rect 343266 269628 343272 269680
rect 343324 269668 343330 269680
rect 352282 269668 352288 269680
rect 343324 269640 352288 269668
rect 343324 269628 343330 269640
rect 352282 269628 352288 269640
rect 352340 269628 352346 269680
rect 361574 269628 361580 269680
rect 361632 269668 361638 269680
rect 382274 269668 382280 269680
rect 361632 269640 382280 269668
rect 361632 269628 361638 269640
rect 382274 269628 382280 269640
rect 382332 269628 382338 269680
rect 382384 269668 382412 269708
rect 382458 269696 382464 269748
rect 382516 269736 382522 269748
rect 544654 269736 544660 269748
rect 382516 269708 544660 269736
rect 382516 269696 382522 269708
rect 544654 269696 544660 269708
rect 544712 269696 544718 269748
rect 551738 269668 551744 269680
rect 382384 269640 551744 269668
rect 551738 269628 551744 269640
rect 551796 269628 551802 269680
rect 188614 269560 188620 269612
rect 188672 269600 188678 269612
rect 200758 269600 200764 269612
rect 188672 269572 200764 269600
rect 188672 269560 188678 269572
rect 200758 269560 200764 269572
rect 200816 269560 200822 269612
rect 207750 269560 207756 269612
rect 207808 269600 207814 269612
rect 245746 269600 245752 269612
rect 207808 269572 245752 269600
rect 207808 269560 207814 269572
rect 245746 269560 245752 269572
rect 245804 269560 245810 269612
rect 281442 269560 281448 269612
rect 281500 269600 281506 269612
rect 302326 269600 302332 269612
rect 281500 269572 302332 269600
rect 281500 269560 281506 269572
rect 302326 269560 302332 269572
rect 302384 269560 302390 269612
rect 310790 269560 310796 269612
rect 310848 269600 310854 269612
rect 380342 269600 380348 269612
rect 310848 269572 380348 269600
rect 310848 269560 310854 269572
rect 380342 269560 380348 269572
rect 380400 269560 380406 269612
rect 380710 269560 380716 269612
rect 380768 269600 380774 269612
rect 565906 269600 565912 269612
rect 380768 269572 565912 269600
rect 380768 269560 380774 269572
rect 565906 269560 565912 269572
rect 565964 269560 565970 269612
rect 94222 269492 94228 269544
rect 94280 269532 94286 269544
rect 202598 269532 202604 269544
rect 94280 269504 202604 269532
rect 94280 269492 94286 269504
rect 202598 269492 202604 269504
rect 202656 269492 202662 269544
rect 202966 269492 202972 269544
rect 203024 269532 203030 269544
rect 226334 269532 226340 269544
rect 203024 269504 226340 269532
rect 203024 269492 203030 269504
rect 226334 269492 226340 269504
rect 226392 269492 226398 269544
rect 226426 269492 226432 269544
rect 226484 269532 226490 269544
rect 234154 269532 234160 269544
rect 226484 269504 234160 269532
rect 226484 269492 226490 269504
rect 234154 269492 234160 269504
rect 234212 269492 234218 269544
rect 280982 269492 280988 269544
rect 281040 269532 281046 269544
rect 301130 269532 301136 269544
rect 281040 269504 301136 269532
rect 281040 269492 281046 269504
rect 301130 269492 301136 269504
rect 301188 269492 301194 269544
rect 312078 269492 312084 269544
rect 312136 269532 312142 269544
rect 383838 269532 383844 269544
rect 312136 269504 383844 269532
rect 312136 269492 312142 269504
rect 383838 269492 383844 269504
rect 383896 269492 383902 269544
rect 386046 269492 386052 269544
rect 386104 269532 386110 269544
rect 580074 269532 580080 269544
rect 386104 269504 580080 269532
rect 386104 269492 386110 269504
rect 580074 269492 580080 269504
rect 580132 269492 580138 269544
rect 198642 269424 198648 269476
rect 198700 269464 198706 269476
rect 239950 269464 239956 269476
rect 198700 269436 239956 269464
rect 198700 269424 198706 269436
rect 239950 269424 239956 269436
rect 240008 269424 240014 269476
rect 282730 269424 282736 269476
rect 282788 269464 282794 269476
rect 305822 269464 305828 269476
rect 282788 269436 305828 269464
rect 282788 269424 282794 269436
rect 305822 269424 305828 269436
rect 305880 269424 305886 269476
rect 313458 269424 313464 269476
rect 313516 269464 313522 269476
rect 387426 269464 387432 269476
rect 313516 269436 387432 269464
rect 313516 269424 313522 269436
rect 387426 269424 387432 269436
rect 387484 269424 387490 269476
rect 388714 269424 388720 269476
rect 388772 269464 388778 269476
rect 587158 269464 587164 269476
rect 388772 269436 587164 269464
rect 388772 269424 388778 269436
rect 587158 269424 587164 269436
rect 587216 269424 587222 269476
rect 74074 269356 74080 269408
rect 74132 269396 74138 269408
rect 195882 269396 195888 269408
rect 74132 269368 195888 269396
rect 74132 269356 74138 269368
rect 195882 269356 195888 269368
rect 195940 269356 195946 269408
rect 204162 269356 204168 269408
rect 204220 269396 204226 269408
rect 244458 269396 244464 269408
rect 204220 269368 244464 269396
rect 204220 269356 204226 269368
rect 244458 269356 244464 269368
rect 244516 269356 244522 269408
rect 282270 269356 282276 269408
rect 282328 269396 282334 269408
rect 304626 269396 304632 269408
rect 282328 269368 304632 269396
rect 282328 269356 282334 269368
rect 304626 269356 304632 269368
rect 304684 269356 304690 269408
rect 314838 269356 314844 269408
rect 314896 269396 314902 269408
rect 390922 269396 390928 269408
rect 314896 269368 390928 269396
rect 314896 269356 314902 269368
rect 390922 269356 390928 269368
rect 390980 269356 390986 269408
rect 394050 269356 394056 269408
rect 394108 269396 394114 269408
rect 601418 269396 601424 269408
rect 394108 269368 601424 269396
rect 394108 269356 394114 269368
rect 601418 269356 601424 269368
rect 601476 269356 601482 269408
rect 80054 269288 80060 269340
rect 80112 269328 80118 269340
rect 197262 269328 197268 269340
rect 80112 269300 197268 269328
rect 80112 269288 80118 269300
rect 197262 269288 197268 269300
rect 197320 269288 197326 269340
rect 197354 269288 197360 269340
rect 197412 269328 197418 269340
rect 241790 269328 241796 269340
rect 197412 269300 241796 269328
rect 197412 269288 197418 269300
rect 241790 269288 241796 269300
rect 241848 269288 241854 269340
rect 283650 269288 283656 269340
rect 283708 269328 283714 269340
rect 308214 269328 308220 269340
rect 283708 269300 308220 269328
rect 283708 269288 283714 269300
rect 308214 269288 308220 269300
rect 308272 269288 308278 269340
rect 315206 269288 315212 269340
rect 315264 269328 315270 269340
rect 392118 269328 392124 269340
rect 315264 269300 392124 269328
rect 315264 269288 315270 269300
rect 392118 269288 392124 269300
rect 392176 269288 392182 269340
rect 396718 269288 396724 269340
rect 396776 269328 396782 269340
rect 608502 269328 608508 269340
rect 396776 269300 608508 269328
rect 396776 269288 396782 269300
rect 608502 269288 608508 269300
rect 608560 269288 608566 269340
rect 81250 269220 81256 269272
rect 81308 269260 81314 269272
rect 198090 269260 198096 269272
rect 81308 269232 198096 269260
rect 81308 269220 81314 269232
rect 198090 269220 198096 269232
rect 198148 269220 198154 269272
rect 200574 269220 200580 269272
rect 200632 269260 200638 269272
rect 243078 269260 243084 269272
rect 200632 269232 243084 269260
rect 200632 269220 200638 269232
rect 243078 269220 243084 269232
rect 243136 269220 243142 269272
rect 283190 269220 283196 269272
rect 283248 269260 283254 269272
rect 307018 269260 307024 269272
rect 283248 269232 307024 269260
rect 283248 269220 283254 269232
rect 307018 269220 307024 269232
rect 307076 269220 307082 269272
rect 317874 269220 317880 269272
rect 317932 269260 317938 269272
rect 399202 269260 399208 269272
rect 317932 269232 399208 269260
rect 317932 269220 317938 269232
rect 399202 269220 399208 269232
rect 399260 269220 399266 269272
rect 399386 269220 399392 269272
rect 399444 269260 399450 269272
rect 615586 269260 615592 269272
rect 399444 269232 615592 269260
rect 399444 269220 399450 269232
rect 615586 269220 615592 269232
rect 615644 269220 615650 269272
rect 71774 269152 71780 269204
rect 71832 269192 71838 269204
rect 194594 269192 194600 269204
rect 71832 269164 194600 269192
rect 71832 269152 71838 269164
rect 194594 269152 194600 269164
rect 194652 269152 194658 269204
rect 195790 269152 195796 269204
rect 195848 269192 195854 269204
rect 241330 269192 241336 269204
rect 195848 269164 241336 269192
rect 195848 269152 195854 269164
rect 241330 269152 241336 269164
rect 241388 269152 241394 269204
rect 284938 269152 284944 269204
rect 284996 269192 285002 269204
rect 311710 269192 311716 269204
rect 284996 269164 311716 269192
rect 284996 269152 285002 269164
rect 311710 269152 311716 269164
rect 311768 269152 311774 269204
rect 320542 269152 320548 269204
rect 320600 269192 320606 269204
rect 406286 269192 406292 269204
rect 320600 269164 406292 269192
rect 320600 269152 320606 269164
rect 406286 269152 406292 269164
rect 406344 269152 406350 269204
rect 411438 269152 411444 269204
rect 411496 269192 411502 269204
rect 647510 269192 647516 269204
rect 411496 269164 647516 269192
rect 411496 269152 411502 269164
rect 647510 269152 647516 269164
rect 647568 269152 647574 269204
rect 193490 269084 193496 269136
rect 193548 269124 193554 269136
rect 240410 269124 240416 269136
rect 193548 269096 240416 269124
rect 193548 269084 193554 269096
rect 240410 269084 240416 269096
rect 240468 269084 240474 269136
rect 284478 269084 284484 269136
rect 284536 269124 284542 269136
rect 310514 269124 310520 269136
rect 284536 269096 310520 269124
rect 284536 269084 284542 269096
rect 310514 269084 310520 269096
rect 310572 269084 310578 269136
rect 323210 269084 323216 269136
rect 323268 269124 323274 269136
rect 411806 269124 411812 269136
rect 323268 269096 411812 269124
rect 323268 269084 323274 269096
rect 411806 269084 411812 269096
rect 411864 269084 411870 269136
rect 411898 269084 411904 269136
rect 411956 269124 411962 269136
rect 648706 269124 648712 269136
rect 411956 269096 648712 269124
rect 411956 269084 411962 269096
rect 648706 269084 648712 269096
rect 648764 269084 648770 269136
rect 152182 269016 152188 269068
rect 152240 269056 152246 269068
rect 224862 269056 224868 269068
rect 152240 269028 224868 269056
rect 152240 269016 152246 269028
rect 224862 269016 224868 269028
rect 224920 269016 224926 269068
rect 226334 269016 226340 269068
rect 226392 269056 226398 269068
rect 243998 269056 244004 269068
rect 226392 269028 244004 269056
rect 226392 269016 226398 269028
rect 243998 269016 244004 269028
rect 244056 269016 244062 269068
rect 292942 269016 292948 269068
rect 293000 269056 293006 269068
rect 333054 269056 333060 269068
rect 293000 269028 333060 269056
rect 293000 269016 293006 269028
rect 333054 269016 333060 269028
rect 333112 269016 333118 269068
rect 351822 269056 351828 269068
rect 342226 269028 351828 269056
rect 159266 268948 159272 269000
rect 159324 268988 159330 269000
rect 227530 268988 227536 269000
rect 159324 268960 227536 268988
rect 159324 268948 159330 268960
rect 227530 268948 227536 268960
rect 227588 268948 227594 269000
rect 232130 268948 232136 269000
rect 232188 268988 232194 269000
rect 237282 268988 237288 269000
rect 232188 268960 237288 268988
rect 232188 268948 232194 268960
rect 237282 268948 237288 268960
rect 237340 268948 237346 269000
rect 269390 268948 269396 269000
rect 269448 268988 269454 269000
rect 270402 268988 270408 269000
rect 269448 268960 270408 268988
rect 269448 268948 269454 268960
rect 270402 268948 270408 268960
rect 270460 268948 270466 269000
rect 295610 268948 295616 269000
rect 295668 268988 295674 269000
rect 329006 268988 329012 269000
rect 295668 268960 329012 268988
rect 295668 268948 295674 268960
rect 329006 268948 329012 268960
rect 329064 268948 329070 269000
rect 330846 268948 330852 269000
rect 330904 268988 330910 269000
rect 342226 268988 342254 269028
rect 351822 269016 351828 269028
rect 351880 269016 351886 269068
rect 473722 269056 473728 269068
rect 351932 269028 473728 269056
rect 330904 268960 342254 268988
rect 330904 268948 330910 268960
rect 345934 268948 345940 269000
rect 345992 268988 345998 269000
rect 351932 268988 351960 269028
rect 473722 269016 473728 269028
rect 473780 269016 473786 269068
rect 345992 268960 351960 268988
rect 345992 268948 345998 268960
rect 352282 268948 352288 269000
rect 352340 268988 352346 269000
rect 466638 268988 466644 269000
rect 352340 268960 466644 268988
rect 352340 268948 352346 268960
rect 466638 268948 466644 268960
rect 466696 268948 466702 269000
rect 160462 268880 160468 268932
rect 160520 268920 160526 268932
rect 228450 268920 228456 268932
rect 160520 268892 228456 268920
rect 160520 268880 160526 268892
rect 228450 268880 228456 268892
rect 228508 268880 228514 268932
rect 230198 268880 230204 268932
rect 230256 268920 230262 268932
rect 238202 268920 238208 268932
rect 230256 268892 238208 268920
rect 230256 268880 230262 268892
rect 238202 268880 238208 268892
rect 238260 268880 238266 268932
rect 309870 268880 309876 268932
rect 309928 268920 309934 268932
rect 331122 268920 331128 268932
rect 309928 268892 331128 268920
rect 309928 268880 309934 268892
rect 331122 268880 331128 268892
rect 331180 268880 331186 268932
rect 351914 268920 351920 268932
rect 331232 268892 351920 268920
rect 161566 268812 161572 268864
rect 161624 268852 161630 268864
rect 227990 268852 227996 268864
rect 161624 268824 227996 268852
rect 161624 268812 161630 268824
rect 227990 268812 227996 268824
rect 228048 268812 228054 268864
rect 229370 268812 229376 268864
rect 229428 268852 229434 268864
rect 239582 268852 239588 268864
rect 229428 268824 239588 268852
rect 229428 268812 229434 268824
rect 239582 268812 239588 268824
rect 239640 268812 239646 268864
rect 328638 268812 328644 268864
rect 328696 268852 328702 268864
rect 331232 268852 331260 268892
rect 351914 268880 351920 268892
rect 351972 268880 351978 268932
rect 352098 268880 352104 268932
rect 352156 268920 352162 268932
rect 468938 268920 468944 268932
rect 352156 268892 468944 268920
rect 352156 268880 352162 268892
rect 468938 268880 468944 268892
rect 468996 268880 469002 268932
rect 328696 268824 331260 268852
rect 328696 268812 328702 268824
rect 341518 268812 341524 268864
rect 341576 268852 341582 268864
rect 461854 268852 461860 268864
rect 341576 268824 461860 268852
rect 341576 268812 341582 268824
rect 461854 268812 461860 268824
rect 461912 268812 461918 268864
rect 166350 268744 166356 268796
rect 166408 268784 166414 268796
rect 230198 268784 230204 268796
rect 166408 268756 230204 268784
rect 166408 268744 166414 268756
rect 230198 268744 230204 268756
rect 230256 268744 230262 268796
rect 340598 268744 340604 268796
rect 340656 268784 340662 268796
rect 459554 268784 459560 268796
rect 340656 268756 459560 268784
rect 340656 268744 340662 268756
rect 459554 268744 459560 268756
rect 459612 268744 459618 268796
rect 167546 268676 167552 268728
rect 167604 268716 167610 268728
rect 231118 268716 231124 268728
rect 167604 268688 231124 268716
rect 167604 268676 167610 268688
rect 231118 268676 231124 268688
rect 231176 268676 231182 268728
rect 273806 268676 273812 268728
rect 273864 268716 273870 268728
rect 282178 268716 282184 268728
rect 273864 268688 282184 268716
rect 273864 268676 273870 268688
rect 282178 268676 282184 268688
rect 282236 268676 282242 268728
rect 338850 268676 338856 268728
rect 338908 268716 338914 268728
rect 454770 268716 454776 268728
rect 338908 268688 454776 268716
rect 338908 268676 338914 268688
rect 454770 268676 454776 268688
rect 454828 268676 454834 268728
rect 173434 268608 173440 268660
rect 173492 268648 173498 268660
rect 232866 268648 232872 268660
rect 173492 268620 232872 268648
rect 173492 268608 173498 268620
rect 232866 268608 232872 268620
rect 232924 268608 232930 268660
rect 250254 268648 250260 268660
rect 235920 268620 250260 268648
rect 168650 268540 168656 268592
rect 168708 268580 168714 268592
rect 230658 268580 230664 268592
rect 168708 268552 230664 268580
rect 168708 268540 168714 268552
rect 230658 268540 230664 268552
rect 230716 268540 230722 268592
rect 156782 268472 156788 268524
rect 156840 268512 156846 268524
rect 212810 268512 212816 268524
rect 156840 268484 212816 268512
rect 156840 268472 156846 268484
rect 212810 268472 212816 268484
rect 212868 268472 212874 268524
rect 219526 268472 219532 268524
rect 219584 268512 219590 268524
rect 235920 268512 235948 268620
rect 250254 268608 250260 268620
rect 250312 268608 250318 268660
rect 337930 268608 337936 268660
rect 337988 268648 337994 268660
rect 452470 268648 452476 268660
rect 337988 268620 452476 268648
rect 337988 268608 337994 268620
rect 452470 268608 452476 268620
rect 452528 268608 452534 268660
rect 240134 268540 240140 268592
rect 240192 268580 240198 268592
rect 244918 268580 244924 268592
rect 240192 268552 244924 268580
rect 240192 268540 240198 268552
rect 244918 268540 244924 268552
rect 244976 268540 244982 268592
rect 336182 268540 336188 268592
rect 336240 268580 336246 268592
rect 447686 268580 447692 268592
rect 336240 268552 447692 268580
rect 336240 268540 336246 268552
rect 447686 268540 447692 268552
rect 447744 268540 447750 268592
rect 219584 268484 235948 268512
rect 219584 268472 219590 268484
rect 335262 268472 335268 268524
rect 335320 268512 335326 268524
rect 445294 268512 445300 268524
rect 335320 268484 445300 268512
rect 335320 268472 335326 268484
rect 445294 268472 445300 268484
rect 445352 268472 445358 268524
rect 174630 268404 174636 268456
rect 174688 268444 174694 268456
rect 233786 268444 233792 268456
rect 174688 268416 233792 268444
rect 174688 268404 174694 268416
rect 233786 268404 233792 268416
rect 233844 268404 233850 268456
rect 234798 268404 234804 268456
rect 234856 268444 234862 268456
rect 239122 268444 239128 268456
rect 234856 268416 239128 268444
rect 234856 268404 234862 268416
rect 239122 268404 239128 268416
rect 239180 268404 239186 268456
rect 276474 268404 276480 268456
rect 276532 268444 276538 268456
rect 289262 268444 289268 268456
rect 276532 268416 289268 268444
rect 276532 268404 276538 268416
rect 289262 268404 289268 268416
rect 289320 268404 289326 268456
rect 325970 268404 325976 268456
rect 326028 268444 326034 268456
rect 332778 268444 332784 268456
rect 326028 268416 332784 268444
rect 326028 268404 326034 268416
rect 332778 268404 332784 268416
rect 332836 268404 332842 268456
rect 333514 268404 333520 268456
rect 333572 268444 333578 268456
rect 440602 268444 440608 268456
rect 333572 268416 440608 268444
rect 333572 268404 333578 268416
rect 440602 268404 440608 268416
rect 440660 268404 440666 268456
rect 179322 268336 179328 268388
rect 179380 268376 179386 268388
rect 233326 268376 233332 268388
rect 179380 268348 233332 268376
rect 179380 268336 179386 268348
rect 233326 268336 233332 268348
rect 233384 268336 233390 268388
rect 275186 268336 275192 268388
rect 275244 268376 275250 268388
rect 285766 268376 285772 268388
rect 275244 268348 285772 268376
rect 275244 268336 275250 268348
rect 285766 268336 285772 268348
rect 285824 268336 285830 268388
rect 309410 268336 309416 268388
rect 309468 268376 309474 268388
rect 332502 268376 332508 268388
rect 309468 268348 332508 268376
rect 309468 268336 309474 268348
rect 332502 268336 332508 268348
rect 332560 268336 332566 268388
rect 332594 268336 332600 268388
rect 332652 268376 332658 268388
rect 438210 268376 438216 268388
rect 332652 268348 438216 268376
rect 332652 268336 332658 268348
rect 438210 268336 438216 268348
rect 438268 268336 438274 268388
rect 180518 268268 180524 268320
rect 180576 268308 180582 268320
rect 235534 268308 235540 268320
rect 180576 268280 235540 268308
rect 180576 268268 180582 268280
rect 235534 268268 235540 268280
rect 235592 268268 235598 268320
rect 274726 268268 274732 268320
rect 274784 268308 274790 268320
rect 284570 268308 284576 268320
rect 274784 268280 284576 268308
rect 274784 268268 274790 268280
rect 284570 268268 284576 268280
rect 284628 268268 284634 268320
rect 312538 268268 312544 268320
rect 312596 268308 312602 268320
rect 312596 268280 332640 268308
rect 312596 268268 312602 268280
rect 181714 268200 181720 268252
rect 181772 268240 181778 268252
rect 236454 268240 236460 268252
rect 181772 268212 236460 268240
rect 181772 268200 181778 268212
rect 236454 268200 236460 268212
rect 236512 268200 236518 268252
rect 275646 268200 275652 268252
rect 275704 268240 275710 268252
rect 286870 268240 286876 268252
rect 275704 268212 286876 268240
rect 275704 268200 275710 268212
rect 286870 268200 286876 268212
rect 286928 268200 286934 268252
rect 316126 268200 316132 268252
rect 316184 268240 316190 268252
rect 316184 268212 332364 268240
rect 316184 268200 316190 268212
rect 206554 268132 206560 268184
rect 206612 268172 206618 268184
rect 245286 268172 245292 268184
rect 206612 268144 245292 268172
rect 206612 268132 206618 268144
rect 245286 268132 245292 268144
rect 245344 268132 245350 268184
rect 316586 268132 316592 268184
rect 316644 268172 316650 268184
rect 326430 268172 326436 268184
rect 316644 268144 326436 268172
rect 316644 268132 316650 268144
rect 326430 268132 326436 268144
rect 326488 268132 326494 268184
rect 184106 268064 184112 268116
rect 184164 268104 184170 268116
rect 236914 268104 236920 268116
rect 184164 268076 236920 268104
rect 184164 268064 184170 268076
rect 236914 268064 236920 268076
rect 236972 268064 236978 268116
rect 82354 267996 82360 268048
rect 82412 268036 82418 268048
rect 198550 268036 198556 268048
rect 82412 268008 198556 268036
rect 82412 267996 82418 268008
rect 198550 267996 198556 268008
rect 198608 267996 198614 268048
rect 201310 267996 201316 268048
rect 201368 268036 201374 268048
rect 203886 268036 203892 268048
rect 201368 268008 203892 268036
rect 201368 267996 201374 268008
rect 203886 267996 203892 268008
rect 203944 267996 203950 268048
rect 206462 267996 206468 268048
rect 206520 268036 206526 268048
rect 225322 268036 225328 268048
rect 206520 268008 225328 268036
rect 206520 267996 206526 268008
rect 225322 267996 225328 268008
rect 225380 267996 225386 268048
rect 231946 267996 231952 268048
rect 232004 268036 232010 268048
rect 235074 268036 235080 268048
rect 232004 268008 235080 268036
rect 232004 267996 232010 268008
rect 235074 267996 235080 268008
rect 235132 267996 235138 268048
rect 319254 267996 319260 268048
rect 319312 268036 319318 268048
rect 326706 268036 326712 268048
rect 319312 268008 326712 268036
rect 319312 267996 319318 268008
rect 326706 267996 326712 268008
rect 326764 267996 326770 268048
rect 197170 267928 197176 267980
rect 197228 267968 197234 267980
rect 216858 267968 216864 267980
rect 197228 267940 216864 267968
rect 197228 267928 197234 267940
rect 216858 267928 216864 267940
rect 216916 267928 216922 267980
rect 232038 267928 232044 267980
rect 232096 267968 232102 267980
rect 235718 267968 235724 267980
rect 232096 267940 235724 267968
rect 232096 267928 232102 267940
rect 235718 267928 235724 267940
rect 235776 267928 235782 267980
rect 298738 267928 298744 267980
rect 298796 267968 298802 267980
rect 307846 267968 307852 267980
rect 298796 267940 307852 267968
rect 298796 267928 298802 267940
rect 307846 267928 307852 267940
rect 307904 267928 307910 267980
rect 321922 267928 321928 267980
rect 321980 267968 321986 267980
rect 325602 267968 325608 267980
rect 321980 267940 325608 267968
rect 321980 267928 321986 267940
rect 325602 267928 325608 267940
rect 325660 267928 325666 267980
rect 332336 267968 332364 268212
rect 332612 268036 332640 268280
rect 351822 268268 351828 268320
rect 351880 268308 351886 268320
rect 433518 268308 433524 268320
rect 351880 268280 433524 268308
rect 351880 268268 351886 268280
rect 433518 268268 433524 268280
rect 433576 268268 433582 268320
rect 332686 268200 332692 268252
rect 332744 268240 332750 268252
rect 426434 268240 426440 268252
rect 332744 268212 426440 268240
rect 332744 268200 332750 268212
rect 426434 268200 426440 268212
rect 426492 268200 426498 268252
rect 351914 268132 351920 268184
rect 351972 268172 351978 268184
rect 427630 268172 427636 268184
rect 351972 268144 427636 268172
rect 351972 268132 351978 268144
rect 427630 268132 427636 268144
rect 427688 268132 427694 268184
rect 332778 268064 332784 268116
rect 332836 268104 332842 268116
rect 420546 268104 420552 268116
rect 332836 268076 420552 268104
rect 332836 268064 332842 268076
rect 420546 268064 420552 268076
rect 420604 268064 420610 268116
rect 663702 268064 663708 268116
rect 663760 268104 663766 268116
rect 676214 268104 676220 268116
rect 663760 268076 676220 268104
rect 663760 268064 663766 268076
rect 676214 268064 676220 268076
rect 676272 268064 676278 268116
rect 357434 268036 357440 268048
rect 332612 268008 357440 268036
rect 357434 267996 357440 268008
rect 357492 267996 357498 268048
rect 357526 267996 357532 268048
rect 357584 268036 357590 268048
rect 358722 268036 358728 268048
rect 357584 268008 358728 268036
rect 357584 267996 357590 268008
rect 358722 267996 358728 268008
rect 358780 267996 358786 268048
rect 372706 267996 372712 268048
rect 372764 268036 372770 268048
rect 382458 268036 382464 268048
rect 372764 268008 382464 268036
rect 372764 267996 372770 268008
rect 382458 267996 382464 268008
rect 382516 267996 382522 268048
rect 390002 267996 390008 268048
rect 390060 268036 390066 268048
rect 394602 268036 394608 268048
rect 390060 268008 394608 268036
rect 390060 267996 390066 268008
rect 394602 267996 394608 268008
rect 394660 267996 394666 268048
rect 400766 267996 400772 268048
rect 400824 268036 400830 268048
rect 402882 268036 402888 268048
rect 400824 268008 402888 268036
rect 400824 267996 400830 268008
rect 402882 267996 402888 268008
rect 402940 267996 402946 268048
rect 406102 267996 406108 268048
rect 406160 268036 406166 268048
rect 412818 268036 412824 268048
rect 406160 268008 412824 268036
rect 406160 267996 406166 268008
rect 412818 267996 412824 268008
rect 412876 267996 412882 268048
rect 352006 267968 352012 267980
rect 332336 267940 352012 267968
rect 352006 267928 352012 267940
rect 352064 267928 352070 267980
rect 661126 267928 661132 267980
rect 661184 267968 661190 267980
rect 676030 267968 676036 267980
rect 661184 267940 676036 267968
rect 661184 267928 661190 267940
rect 676030 267928 676036 267940
rect 676088 267928 676094 267980
rect 88334 267860 88340 267912
rect 88392 267900 88398 267912
rect 201218 267900 201224 267912
rect 88392 267872 201224 267900
rect 88392 267860 88398 267872
rect 201218 267860 201224 267872
rect 201276 267860 201282 267912
rect 211246 267860 211252 267912
rect 211304 267900 211310 267912
rect 247126 267900 247132 267912
rect 211304 267872 247132 267900
rect 211304 267860 211310 267872
rect 247126 267860 247132 267872
rect 247184 267860 247190 267912
rect 276290 267860 276296 267912
rect 276348 267900 276354 267912
rect 288066 267900 288072 267912
rect 276348 267872 288072 267900
rect 276348 267860 276354 267872
rect 288066 267860 288072 267872
rect 288124 267860 288130 267912
rect 297910 267860 297916 267912
rect 297968 267900 297974 267912
rect 304902 267900 304908 267912
rect 297968 267872 304908 267900
rect 297968 267860 297974 267872
rect 304902 267860 304908 267872
rect 304960 267860 304966 267912
rect 327994 267860 328000 267912
rect 328052 267900 328058 267912
rect 332686 267900 332692 267912
rect 328052 267872 332692 267900
rect 328052 267860 328058 267872
rect 332686 267860 332692 267872
rect 332744 267860 332750 267912
rect 344186 267860 344192 267912
rect 344244 267900 344250 267912
rect 352098 267900 352104 267912
rect 344244 267872 352104 267900
rect 344244 267860 344250 267872
rect 352098 267860 352104 267872
rect 352156 267860 352162 267912
rect 95418 267792 95424 267844
rect 95476 267832 95482 267844
rect 203518 267832 203524 267844
rect 95476 267804 203524 267832
rect 95476 267792 95482 267804
rect 203518 267792 203524 267804
rect 203576 267792 203582 267844
rect 205542 267792 205548 267844
rect 205600 267832 205606 267844
rect 212350 267832 212356 267844
rect 205600 267804 212356 267832
rect 205600 267792 205606 267804
rect 212350 267792 212356 267804
rect 212408 267792 212414 267844
rect 234706 267792 234712 267844
rect 234764 267832 234770 267844
rect 237742 267832 237748 267844
rect 234764 267804 237748 267832
rect 234764 267792 234770 267804
rect 237742 267792 237748 267804
rect 237800 267792 237806 267844
rect 304534 267792 304540 267844
rect 304592 267832 304598 267844
rect 351730 267832 351736 267844
rect 304592 267804 351736 267832
rect 304592 267792 304598 267804
rect 351730 267792 351736 267804
rect 351788 267792 351794 267844
rect 202690 267724 202696 267776
rect 202748 267764 202754 267776
rect 206554 267764 206560 267776
rect 202748 267736 206560 267764
rect 202748 267724 202754 267736
rect 206554 267724 206560 267736
rect 206612 267724 206618 267776
rect 232498 267724 232504 267776
rect 232556 267764 232562 267776
rect 238662 267764 238668 267776
rect 232556 267736 238668 267764
rect 232556 267724 232562 267736
rect 238662 267724 238668 267736
rect 238720 267724 238726 267776
rect 332502 267724 332508 267776
rect 332560 267764 332566 267776
rect 376754 267764 376760 267776
rect 332560 267736 376760 267764
rect 332560 267724 332566 267736
rect 376754 267724 376760 267736
rect 376812 267724 376818 267776
rect 661034 267724 661040 267776
rect 661092 267764 661098 267776
rect 676122 267764 676128 267776
rect 661092 267736 676128 267764
rect 661092 267724 661098 267736
rect 676122 267724 676128 267736
rect 676180 267724 676186 267776
rect 359734 267656 359740 267708
rect 359792 267696 359798 267708
rect 510338 267696 510344 267708
rect 359792 267668 510344 267696
rect 359792 267656 359798 267668
rect 510338 267656 510344 267668
rect 510396 267656 510402 267708
rect 674742 267656 674748 267708
rect 674800 267696 674806 267708
rect 676030 267696 676036 267708
rect 674800 267668 676036 267696
rect 674800 267656 674806 267668
rect 676030 267656 676036 267668
rect 676088 267656 676094 267708
rect 362402 267588 362408 267640
rect 362460 267628 362466 267640
rect 517422 267628 517428 267640
rect 362460 267600 517428 267628
rect 362460 267588 362466 267600
rect 517422 267588 517428 267600
rect 517480 267588 517486 267640
rect 365070 267520 365076 267572
rect 365128 267560 365134 267572
rect 524506 267560 524512 267572
rect 365128 267532 524512 267560
rect 365128 267520 365134 267532
rect 524506 267520 524512 267532
rect 524564 267520 524570 267572
rect 367738 267452 367744 267504
rect 367796 267492 367802 267504
rect 531590 267492 531596 267504
rect 367796 267464 531596 267492
rect 367796 267452 367802 267464
rect 531590 267452 531596 267464
rect 531648 267452 531654 267504
rect 672258 267452 672264 267504
rect 672316 267492 672322 267504
rect 675938 267492 675944 267504
rect 672316 267464 675944 267492
rect 672316 267452 672322 267464
rect 675938 267452 675944 267464
rect 675996 267452 676002 267504
rect 370498 267384 370504 267436
rect 370556 267424 370562 267436
rect 538766 267424 538772 267436
rect 370556 267396 538772 267424
rect 370556 267384 370562 267396
rect 538766 267384 538772 267396
rect 538824 267384 538830 267436
rect 373534 267316 373540 267368
rect 373592 267356 373598 267368
rect 547046 267356 547052 267368
rect 373592 267328 547052 267356
rect 373592 267316 373598 267328
rect 547046 267316 547052 267328
rect 547104 267316 547110 267368
rect 374454 267248 374460 267300
rect 374512 267288 374518 267300
rect 549346 267288 549352 267300
rect 374512 267260 549352 267288
rect 374512 267248 374518 267260
rect 549346 267248 549352 267260
rect 549404 267248 549410 267300
rect 376202 267180 376208 267232
rect 376260 267220 376266 267232
rect 554130 267220 554136 267232
rect 376260 267192 554136 267220
rect 376260 267180 376266 267192
rect 554130 267180 554136 267192
rect 554188 267180 554194 267232
rect 299658 267112 299664 267164
rect 299716 267152 299722 267164
rect 350718 267152 350724 267164
rect 299716 267124 350724 267152
rect 299716 267112 299722 267124
rect 350718 267112 350724 267124
rect 350776 267112 350782 267164
rect 375834 267112 375840 267164
rect 375892 267152 375898 267164
rect 552934 267152 552940 267164
rect 375892 267124 552940 267152
rect 375892 267112 375898 267124
rect 552934 267112 552940 267124
rect 552992 267112 552998 267164
rect 300946 267044 300952 267096
rect 301004 267084 301010 267096
rect 354306 267084 354312 267096
rect 301004 267056 354312 267084
rect 301004 267044 301010 267056
rect 354306 267044 354312 267056
rect 354364 267044 354370 267096
rect 377122 267044 377128 267096
rect 377180 267084 377186 267096
rect 556430 267084 556436 267096
rect 377180 267056 556436 267084
rect 377180 267044 377186 267056
rect 556430 267044 556436 267056
rect 556488 267044 556494 267096
rect 302326 266976 302332 267028
rect 302384 267016 302390 267028
rect 357894 267016 357900 267028
rect 302384 266988 357900 267016
rect 302384 266976 302390 266988
rect 357894 266976 357900 266988
rect 357952 266976 357958 267028
rect 378502 266976 378508 267028
rect 378560 267016 378566 267028
rect 560018 267016 560024 267028
rect 378560 266988 560024 267016
rect 378560 266976 378566 266988
rect 560018 266976 560024 266988
rect 560076 266976 560082 267028
rect 303706 266908 303712 266960
rect 303764 266948 303770 266960
rect 361390 266948 361396 266960
rect 303764 266920 361396 266948
rect 303764 266908 303770 266920
rect 361390 266908 361396 266920
rect 361448 266908 361454 266960
rect 378870 266908 378876 266960
rect 378928 266948 378934 266960
rect 561214 266948 561220 266960
rect 378928 266920 561220 266948
rect 378928 266908 378934 266920
rect 561214 266908 561220 266920
rect 561272 266908 561278 266960
rect 304994 266840 305000 266892
rect 305052 266880 305058 266892
rect 364978 266880 364984 266892
rect 305052 266852 364984 266880
rect 305052 266840 305058 266852
rect 364978 266840 364984 266852
rect 365036 266840 365042 266892
rect 379790 266840 379796 266892
rect 379848 266880 379854 266892
rect 563514 266880 563520 266892
rect 379848 266852 563520 266880
rect 379848 266840 379854 266852
rect 563514 266840 563520 266852
rect 563572 266840 563578 266892
rect 306374 266772 306380 266824
rect 306432 266812 306438 266824
rect 368474 266812 368480 266824
rect 306432 266784 368480 266812
rect 306432 266772 306438 266784
rect 368474 266772 368480 266784
rect 368532 266772 368538 266824
rect 381630 266772 381636 266824
rect 381688 266812 381694 266824
rect 568298 266812 568304 266824
rect 381688 266784 568304 266812
rect 381688 266772 381694 266784
rect 568298 266772 568304 266784
rect 568356 266772 568362 266824
rect 307662 266704 307668 266756
rect 307720 266744 307726 266756
rect 372062 266744 372068 266756
rect 307720 266716 372068 266744
rect 307720 266704 307726 266716
rect 372062 266704 372068 266716
rect 372120 266704 372126 266756
rect 381170 266704 381176 266756
rect 381228 266744 381234 266756
rect 567102 266744 567108 266756
rect 381228 266716 567108 266744
rect 381228 266704 381234 266716
rect 567102 266704 567108 266716
rect 567160 266704 567166 266756
rect 309042 266636 309048 266688
rect 309100 266676 309106 266688
rect 375558 266676 375564 266688
rect 309100 266648 375564 266676
rect 309100 266636 309106 266648
rect 375558 266636 375564 266648
rect 375616 266636 375622 266688
rect 382458 266636 382464 266688
rect 382516 266676 382522 266688
rect 570690 266676 570696 266688
rect 382516 266648 570696 266676
rect 382516 266636 382522 266648
rect 570690 266636 570696 266648
rect 570748 266636 570754 266688
rect 123754 266568 123760 266620
rect 123812 266608 123818 266620
rect 214190 266608 214196 266620
rect 123812 266580 214196 266608
rect 123812 266568 123818 266580
rect 214190 266568 214196 266580
rect 214248 266568 214254 266620
rect 310330 266568 310336 266620
rect 310388 266608 310394 266620
rect 379146 266608 379152 266620
rect 310388 266580 379152 266608
rect 310388 266568 310394 266580
rect 379146 266568 379152 266580
rect 379204 266568 379210 266620
rect 384298 266568 384304 266620
rect 384356 266608 384362 266620
rect 575382 266608 575388 266620
rect 384356 266580 575388 266608
rect 384356 266568 384362 266580
rect 575382 266568 575388 266580
rect 575440 266568 575446 266620
rect 116670 266500 116676 266552
rect 116728 266540 116734 266552
rect 211522 266540 211528 266552
rect 116728 266512 211528 266540
rect 116728 266500 116734 266512
rect 211522 266500 211528 266512
rect 211580 266500 211586 266552
rect 311710 266500 311716 266552
rect 311768 266540 311774 266552
rect 382642 266540 382648 266552
rect 311768 266512 382648 266540
rect 311768 266500 311774 266512
rect 382642 266500 382648 266512
rect 382700 266500 382706 266552
rect 383838 266500 383844 266552
rect 383896 266540 383902 266552
rect 574186 266540 574192 266552
rect 383896 266512 574192 266540
rect 383896 266500 383902 266512
rect 574186 266500 574192 266512
rect 574244 266500 574250 266552
rect 72970 266432 72976 266484
rect 73028 266472 73034 266484
rect 195054 266472 195060 266484
rect 73028 266444 195060 266472
rect 73028 266432 73034 266444
rect 195054 266432 195060 266444
rect 195112 266432 195118 266484
rect 312998 266432 313004 266484
rect 313056 266472 313062 266484
rect 386230 266472 386236 266484
rect 313056 266444 386236 266472
rect 313056 266432 313062 266444
rect 386230 266432 386236 266444
rect 386288 266432 386294 266484
rect 389174 266432 389180 266484
rect 389232 266472 389238 266484
rect 588354 266472 588360 266484
rect 389232 266444 588360 266472
rect 389232 266432 389238 266444
rect 588354 266432 588360 266444
rect 588412 266432 588418 266484
rect 113174 266364 113180 266416
rect 113232 266404 113238 266416
rect 210142 266404 210148 266416
rect 113232 266376 210148 266404
rect 113232 266364 113238 266376
rect 210142 266364 210148 266376
rect 210200 266364 210206 266416
rect 315666 266364 315672 266416
rect 315724 266404 315730 266416
rect 315724 266376 391934 266404
rect 315724 266364 315730 266376
rect 68186 266296 68192 266348
rect 68244 266336 68250 266348
rect 193214 266336 193220 266348
rect 68244 266308 193220 266336
rect 68244 266296 68250 266308
rect 193214 266296 193220 266308
rect 193272 266296 193278 266348
rect 317046 266296 317052 266348
rect 317104 266336 317110 266348
rect 382182 266336 382188 266348
rect 317104 266308 382188 266336
rect 317104 266296 317110 266308
rect 382182 266296 382188 266308
rect 382240 266296 382246 266348
rect 391906 266336 391934 266376
rect 392302 266364 392308 266416
rect 392360 266404 392366 266416
rect 596634 266404 596640 266416
rect 392360 266376 596640 266404
rect 392360 266364 392366 266376
rect 596634 266364 596640 266376
rect 596692 266364 596698 266416
rect 393314 266336 393320 266348
rect 391906 266308 393320 266336
rect 393314 266296 393320 266308
rect 393372 266296 393378 266348
rect 394970 266296 394976 266348
rect 395028 266336 395034 266348
rect 603718 266336 603724 266348
rect 395028 266308 603724 266336
rect 395028 266296 395034 266308
rect 603718 266296 603724 266308
rect 603776 266296 603782 266348
rect 652938 266296 652944 266348
rect 652996 266336 653002 266348
rect 675662 266336 675668 266348
rect 652996 266308 675668 266336
rect 652996 266296 653002 266308
rect 675662 266296 675668 266308
rect 675720 266296 675726 266348
rect 357066 266228 357072 266280
rect 357124 266268 357130 266280
rect 503254 266268 503260 266280
rect 357124 266240 503260 266268
rect 357124 266228 357130 266240
rect 503254 266228 503260 266240
rect 503312 266228 503318 266280
rect 353110 266160 353116 266212
rect 353168 266200 353174 266212
rect 492582 266200 492588 266212
rect 353168 266172 492588 266200
rect 353168 266160 353174 266172
rect 492582 266160 492588 266172
rect 492640 266160 492646 266212
rect 351730 266092 351736 266144
rect 351788 266132 351794 266144
rect 489086 266132 489092 266144
rect 351788 266104 489092 266132
rect 351788 266092 351794 266104
rect 489086 266092 489092 266104
rect 489144 266092 489150 266144
rect 673270 266092 673276 266144
rect 673328 266132 673334 266144
rect 676214 266132 676220 266144
rect 673328 266104 676220 266132
rect 673328 266092 673334 266104
rect 676214 266092 676220 266104
rect 676272 266092 676278 266144
rect 347774 266024 347780 266076
rect 347832 266064 347838 266076
rect 478414 266064 478420 266076
rect 347832 266036 478420 266064
rect 347832 266024 347838 266036
rect 478414 266024 478420 266036
rect 478472 266024 478478 266076
rect 346394 265956 346400 266008
rect 346452 265996 346458 266008
rect 474918 265996 474924 266008
rect 346452 265968 474924 265996
rect 346452 265956 346458 265968
rect 474918 265956 474924 265968
rect 474976 265956 474982 266008
rect 339770 265888 339776 265940
rect 339828 265928 339834 265940
rect 457162 265928 457168 265940
rect 339828 265900 457168 265928
rect 339828 265888 339834 265900
rect 457162 265888 457168 265900
rect 457220 265888 457226 265940
rect 338390 265820 338396 265872
rect 338448 265860 338454 265872
rect 453574 265860 453580 265872
rect 338448 265832 453580 265860
rect 338448 265820 338454 265832
rect 453574 265820 453580 265832
rect 453632 265820 453638 265872
rect 317506 265752 317512 265804
rect 317564 265792 317570 265804
rect 382090 265792 382096 265804
rect 317564 265764 382096 265792
rect 317564 265752 317570 265764
rect 382090 265752 382096 265764
rect 382148 265752 382154 265804
rect 382182 265752 382188 265804
rect 382240 265792 382246 265804
rect 396902 265792 396908 265804
rect 382240 265764 396908 265792
rect 382240 265752 382246 265764
rect 396902 265752 396908 265764
rect 396960 265752 396966 265804
rect 397638 265752 397644 265804
rect 397696 265792 397702 265804
rect 511626 265792 511632 265804
rect 397696 265764 511632 265792
rect 397696 265752 397702 265764
rect 511626 265752 511632 265764
rect 511684 265752 511690 265804
rect 329466 265684 329472 265736
rect 329524 265724 329530 265736
rect 429930 265724 429936 265736
rect 329524 265696 353294 265724
rect 329524 265684 329530 265696
rect 353266 265656 353294 265696
rect 382200 265696 429936 265724
rect 382200 265656 382228 265696
rect 429930 265684 429936 265696
rect 429988 265684 429994 265736
rect 353266 265628 382228 265656
rect 382274 265616 382280 265668
rect 382332 265656 382338 265668
rect 398006 265656 398012 265668
rect 382332 265628 398012 265656
rect 382332 265616 382338 265628
rect 398006 265616 398012 265628
rect 398064 265616 398070 265668
rect 400306 265616 400312 265668
rect 400364 265656 400370 265668
rect 498838 265656 498844 265668
rect 400364 265628 498844 265656
rect 400364 265616 400370 265628
rect 498838 265616 498844 265628
rect 498896 265616 498902 265668
rect 325510 265548 325516 265600
rect 325568 265588 325574 265600
rect 419350 265588 419356 265600
rect 325568 265560 419356 265588
rect 325568 265548 325574 265560
rect 419350 265548 419356 265560
rect 419408 265548 419414 265600
rect 324130 265480 324136 265532
rect 324188 265520 324194 265532
rect 415762 265520 415768 265532
rect 324188 265492 415768 265520
rect 324188 265480 324194 265492
rect 415762 265480 415768 265492
rect 415820 265480 415826 265532
rect 322934 265412 322940 265464
rect 322992 265452 322998 265464
rect 412266 265452 412272 265464
rect 322992 265424 412272 265452
rect 322992 265412 322998 265424
rect 412266 265412 412272 265424
rect 412324 265412 412330 265464
rect 321462 265344 321468 265396
rect 321520 265384 321526 265396
rect 408678 265384 408684 265396
rect 321520 265356 408684 265384
rect 321520 265344 321526 265356
rect 408678 265344 408684 265356
rect 408736 265344 408742 265396
rect 674742 265344 674748 265396
rect 674800 265384 674806 265396
rect 676030 265384 676036 265396
rect 674800 265356 676036 265384
rect 674800 265344 674806 265356
rect 676030 265344 676036 265356
rect 676088 265344 676094 265396
rect 318334 265276 318340 265328
rect 318392 265316 318398 265328
rect 400398 265316 400404 265328
rect 318392 265288 400404 265316
rect 318392 265276 318398 265288
rect 400398 265276 400404 265288
rect 400456 265276 400462 265328
rect 402974 265276 402980 265328
rect 403032 265316 403038 265328
rect 471974 265316 471980 265328
rect 403032 265288 471980 265316
rect 403032 265276 403038 265288
rect 471974 265276 471980 265288
rect 472032 265276 472038 265328
rect 314378 265208 314384 265260
rect 314436 265248 314442 265260
rect 389726 265248 389732 265260
rect 314436 265220 389732 265248
rect 314436 265208 314442 265220
rect 389726 265208 389732 265220
rect 389784 265208 389790 265260
rect 319714 265140 319720 265192
rect 319772 265180 319778 265192
rect 403986 265180 403992 265192
rect 319772 265152 403992 265180
rect 319772 265140 319778 265152
rect 403986 265140 403992 265152
rect 404044 265140 404050 265192
rect 658274 265004 658280 265056
rect 658332 265044 658338 265056
rect 675754 265044 675760 265056
rect 658332 265016 675760 265044
rect 658332 265004 658338 265016
rect 675754 265004 675760 265016
rect 675812 265004 675818 265056
rect 671890 264936 671896 264988
rect 671948 264976 671954 264988
rect 676214 264976 676220 264988
rect 671948 264948 676220 264976
rect 671948 264936 671954 264948
rect 676214 264936 676220 264948
rect 676272 264936 676278 264988
rect 674190 263032 674196 263084
rect 674248 263072 674254 263084
rect 676030 263072 676036 263084
rect 674248 263044 676036 263072
rect 674248 263032 674254 263044
rect 676030 263032 676036 263044
rect 676088 263032 676094 263084
rect 674006 262488 674012 262540
rect 674064 262528 674070 262540
rect 676122 262528 676128 262540
rect 674064 262500 676128 262528
rect 674064 262488 674070 262500
rect 676122 262488 676128 262500
rect 676180 262488 676186 262540
rect 673730 262284 673736 262336
rect 673788 262324 673794 262336
rect 676122 262324 676128 262336
rect 673788 262296 676128 262324
rect 673788 262284 673794 262296
rect 676122 262284 676128 262296
rect 676180 262284 676186 262336
rect 416774 262216 416780 262268
rect 416832 262256 416838 262268
rect 571702 262256 571708 262268
rect 416832 262228 571708 262256
rect 416832 262216 416838 262228
rect 571702 262216 571708 262228
rect 571760 262216 571766 262268
rect 674282 262216 674288 262268
rect 674340 262256 674346 262268
rect 676030 262256 676036 262268
rect 674340 262228 676036 262256
rect 674340 262216 674346 262228
rect 676030 262216 676036 262228
rect 676088 262216 676094 262268
rect 674098 261808 674104 261860
rect 674156 261848 674162 261860
rect 676030 261848 676036 261860
rect 674156 261820 676036 261848
rect 674156 261808 674162 261820
rect 676030 261808 676036 261820
rect 676088 261808 676094 261860
rect 673454 260176 673460 260228
rect 673512 260216 673518 260228
rect 675570 260216 675576 260228
rect 673512 260188 675576 260216
rect 673512 260176 673518 260188
rect 675570 260176 675576 260188
rect 675628 260176 675634 260228
rect 673546 259700 673552 259752
rect 673604 259740 673610 259752
rect 675570 259740 675576 259752
rect 673604 259712 675576 259740
rect 673604 259700 673610 259712
rect 675570 259700 675576 259712
rect 675628 259700 675634 259752
rect 674466 259632 674472 259684
rect 674524 259672 674530 259684
rect 676122 259672 676128 259684
rect 674524 259644 676128 259672
rect 674524 259632 674530 259644
rect 676122 259632 676128 259644
rect 676180 259632 676186 259684
rect 674374 259564 674380 259616
rect 674432 259604 674438 259616
rect 675938 259604 675944 259616
rect 674432 259576 675944 259604
rect 674432 259564 674438 259576
rect 675938 259564 675944 259576
rect 675996 259564 676002 259616
rect 675018 259496 675024 259548
rect 675076 259536 675082 259548
rect 676122 259536 676128 259548
rect 675076 259508 676128 259536
rect 675076 259496 675082 259508
rect 676122 259496 676128 259508
rect 676180 259496 676186 259548
rect 675202 259428 675208 259480
rect 675260 259468 675266 259480
rect 676030 259468 676036 259480
rect 675260 259440 676036 259468
rect 675260 259428 675266 259440
rect 676030 259428 676036 259440
rect 676088 259428 676094 259480
rect 41506 258340 41512 258392
rect 41564 258380 41570 258392
rect 48406 258380 48412 258392
rect 41564 258352 48412 258380
rect 41564 258340 41570 258352
rect 48406 258340 48412 258352
rect 48464 258340 48470 258392
rect 41506 258000 41512 258052
rect 41564 258040 41570 258052
rect 53926 258040 53932 258052
rect 41564 258012 53932 258040
rect 41564 258000 41570 258012
rect 53926 258000 53932 258012
rect 53984 258000 53990 258052
rect 41506 257524 41512 257576
rect 41564 257564 41570 257576
rect 50982 257564 50988 257576
rect 41564 257536 50988 257564
rect 41564 257524 41570 257536
rect 50982 257524 50988 257536
rect 51040 257524 51046 257576
rect 41782 256844 41788 256896
rect 41840 256884 41846 256896
rect 45830 256884 45836 256896
rect 41840 256856 45836 256884
rect 41840 256844 41846 256856
rect 45830 256844 45836 256856
rect 45888 256844 45894 256896
rect 672810 256844 672816 256896
rect 672868 256884 672874 256896
rect 678974 256884 678980 256896
rect 672868 256856 678980 256884
rect 672868 256844 672874 256856
rect 678974 256844 678980 256856
rect 679032 256844 679038 256896
rect 673638 256776 673644 256828
rect 673696 256816 673702 256828
rect 676122 256816 676128 256828
rect 673696 256788 676128 256816
rect 673696 256776 673702 256788
rect 676122 256776 676128 256788
rect 676180 256776 676186 256828
rect 52270 256708 52276 256760
rect 52328 256748 52334 256760
rect 184934 256748 184940 256760
rect 52328 256720 184940 256748
rect 52328 256708 52334 256720
rect 184934 256708 184940 256720
rect 184992 256708 184998 256760
rect 416774 256708 416780 256760
rect 416832 256748 416838 256760
rect 571794 256748 571800 256760
rect 416832 256720 571800 256748
rect 416832 256708 416838 256720
rect 571794 256708 571800 256720
rect 571852 256708 571858 256760
rect 673822 256708 673828 256760
rect 673880 256748 673886 256760
rect 676030 256748 676036 256760
rect 673880 256720 676036 256748
rect 673880 256708 673886 256720
rect 676030 256708 676036 256720
rect 676088 256708 676094 256760
rect 674742 255280 674748 255332
rect 674800 255320 674806 255332
rect 675662 255320 675668 255332
rect 674800 255292 675668 255320
rect 674800 255280 674806 255292
rect 675662 255280 675668 255292
rect 675720 255280 675726 255332
rect 674650 255212 674656 255264
rect 674708 255252 674714 255264
rect 675754 255252 675760 255264
rect 674708 255224 675760 255252
rect 674708 255212 674714 255224
rect 675754 255212 675760 255224
rect 675812 255212 675818 255264
rect 416774 253920 416780 253972
rect 416832 253960 416838 253972
rect 571518 253960 571524 253972
rect 416832 253932 571524 253960
rect 416832 253920 416838 253932
rect 571518 253920 571524 253932
rect 571576 253920 571582 253972
rect 416774 251200 416780 251252
rect 416832 251240 416838 251252
rect 574094 251240 574100 251252
rect 416832 251212 574100 251240
rect 416832 251200 416838 251212
rect 574094 251200 574100 251212
rect 574152 251200 574158 251252
rect 675754 251200 675760 251252
rect 675812 251200 675818 251252
rect 675772 250980 675800 251200
rect 675754 250928 675760 250980
rect 675812 250928 675818 250980
rect 675202 250384 675208 250436
rect 675260 250424 675266 250436
rect 675478 250424 675484 250436
rect 675260 250396 675484 250424
rect 675260 250384 675266 250396
rect 675478 250384 675484 250396
rect 675536 250384 675542 250436
rect 33042 249772 33048 249824
rect 33100 249812 33106 249824
rect 43622 249812 43628 249824
rect 33100 249784 43628 249812
rect 33100 249772 33106 249784
rect 43622 249772 43628 249784
rect 43680 249772 43686 249824
rect 674190 249568 674196 249620
rect 674248 249608 674254 249620
rect 675386 249608 675392 249620
rect 674248 249580 675392 249608
rect 674248 249568 674254 249580
rect 675386 249568 675392 249580
rect 675444 249568 675450 249620
rect 416774 248412 416780 248464
rect 416832 248452 416838 248464
rect 574186 248452 574192 248464
rect 416832 248424 574192 248452
rect 416832 248412 416838 248424
rect 574186 248412 574192 248424
rect 574244 248412 574250 248464
rect 674282 247868 674288 247920
rect 674340 247908 674346 247920
rect 675478 247908 675484 247920
rect 674340 247880 675484 247908
rect 674340 247868 674346 247880
rect 675478 247868 675484 247880
rect 675536 247868 675542 247920
rect 41506 247664 41512 247716
rect 41564 247704 41570 247716
rect 45922 247704 45928 247716
rect 41564 247676 45928 247704
rect 41564 247664 41570 247676
rect 45922 247664 45928 247676
rect 45980 247664 45986 247716
rect 41506 247256 41512 247308
rect 41564 247296 41570 247308
rect 45830 247296 45836 247308
rect 41564 247268 45836 247296
rect 41564 247256 41570 247268
rect 45830 247256 45836 247268
rect 45888 247256 45894 247308
rect 674466 247256 674472 247308
rect 674524 247296 674530 247308
rect 675386 247296 675392 247308
rect 674524 247268 675392 247296
rect 674524 247256 674530 247268
rect 675386 247256 675392 247268
rect 675444 247256 675450 247308
rect 674374 246508 674380 246560
rect 674432 246548 674438 246560
rect 675386 246548 675392 246560
rect 674432 246520 675392 246548
rect 674432 246508 674438 246520
rect 675386 246508 675392 246520
rect 675444 246508 675450 246560
rect 41506 246440 41512 246492
rect 41564 246480 41570 246492
rect 45738 246480 45744 246492
rect 41564 246452 45744 246480
rect 41564 246440 41570 246452
rect 45738 246440 45744 246452
rect 45796 246440 45802 246492
rect 675110 246032 675116 246084
rect 675168 246072 675174 246084
rect 675386 246072 675392 246084
rect 675168 246044 675392 246072
rect 675168 246032 675174 246044
rect 675386 246032 675392 246044
rect 675444 246032 675450 246084
rect 52178 245624 52184 245676
rect 52236 245664 52242 245676
rect 184934 245664 184940 245676
rect 52236 245636 184940 245664
rect 52236 245624 52242 245636
rect 184934 245624 184940 245636
rect 184992 245624 184998 245676
rect 416774 245624 416780 245676
rect 416832 245664 416838 245676
rect 571610 245664 571616 245676
rect 416832 245636 571616 245664
rect 416832 245624 416838 245636
rect 571610 245624 571616 245636
rect 571668 245624 571674 245676
rect 42702 244468 42708 244520
rect 42760 244508 42766 244520
rect 43530 244508 43536 244520
rect 42760 244480 43536 244508
rect 42760 244468 42766 244480
rect 43530 244468 43536 244480
rect 43588 244468 43594 244520
rect 32950 244400 32956 244452
rect 33008 244440 33014 244452
rect 43070 244440 43076 244452
rect 33008 244412 43076 244440
rect 33008 244400 33014 244412
rect 43070 244400 43076 244412
rect 43128 244400 43134 244452
rect 33042 244332 33048 244384
rect 33100 244372 33106 244384
rect 42886 244372 42892 244384
rect 33100 244344 42892 244372
rect 33100 244332 33106 244344
rect 42886 244332 42892 244344
rect 42944 244332 42950 244384
rect 31662 244264 31668 244316
rect 31720 244304 31726 244316
rect 42702 244304 42708 244316
rect 31720 244276 42708 244304
rect 31720 244264 31726 244276
rect 42702 244264 42708 244276
rect 42760 244264 42766 244316
rect 32858 244196 32864 244248
rect 32916 244236 32922 244248
rect 42978 244236 42984 244248
rect 32916 244208 42984 244236
rect 32916 244196 32922 244208
rect 42978 244196 42984 244208
rect 43036 244196 43042 244248
rect 673730 243584 673736 243636
rect 673788 243624 673794 243636
rect 675294 243624 675300 243636
rect 673788 243596 675300 243624
rect 673788 243584 673794 243596
rect 675294 243584 675300 243596
rect 675352 243584 675358 243636
rect 42426 243312 42432 243364
rect 42484 243352 42490 243364
rect 43806 243352 43812 243364
rect 42484 243324 43812 243352
rect 42484 243312 42490 243324
rect 43806 243312 43812 243324
rect 43864 243312 43870 243364
rect 43346 243108 43352 243160
rect 43404 243148 43410 243160
rect 43622 243148 43628 243160
rect 43404 243120 43628 243148
rect 43404 243108 43410 243120
rect 43622 243108 43628 243120
rect 43680 243108 43686 243160
rect 42794 242972 42800 243024
rect 42852 243012 42858 243024
rect 43346 243012 43352 243024
rect 42852 242984 43352 243012
rect 42852 242972 42858 242984
rect 43346 242972 43352 242984
rect 43404 242972 43410 243024
rect 673822 242904 673828 242956
rect 673880 242944 673886 242956
rect 675294 242944 675300 242956
rect 673880 242916 675300 242944
rect 673880 242904 673886 242916
rect 675294 242904 675300 242916
rect 675352 242904 675358 242956
rect 38286 242836 38292 242888
rect 38344 242876 38350 242888
rect 42794 242876 42800 242888
rect 38344 242848 42800 242876
rect 38344 242836 38350 242848
rect 42794 242836 42800 242848
rect 42852 242836 42858 242888
rect 673546 242156 673552 242208
rect 673604 242196 673610 242208
rect 675386 242196 675392 242208
rect 673604 242168 675392 242196
rect 673604 242156 673610 242168
rect 675386 242156 675392 242168
rect 675444 242156 675450 242208
rect 674374 241884 674380 241936
rect 674432 241924 674438 241936
rect 675294 241924 675300 241936
rect 674432 241896 675300 241924
rect 674432 241884 674438 241896
rect 675294 241884 675300 241896
rect 675352 241884 675358 241936
rect 673638 241544 673644 241596
rect 673696 241584 673702 241596
rect 675386 241584 675392 241596
rect 673696 241556 675392 241584
rect 673696 241544 673702 241556
rect 675386 241544 675392 241556
rect 675444 241544 675450 241596
rect 673454 240524 673460 240576
rect 673512 240564 673518 240576
rect 675386 240564 675392 240576
rect 673512 240536 675392 240564
rect 673512 240524 673518 240536
rect 675386 240524 675392 240536
rect 675444 240524 675450 240576
rect 42150 240320 42156 240372
rect 42208 240360 42214 240372
rect 42426 240360 42432 240372
rect 42208 240332 42432 240360
rect 42208 240320 42214 240332
rect 42426 240320 42432 240332
rect 42484 240320 42490 240372
rect 42150 238416 42156 238468
rect 42208 238456 42214 238468
rect 42702 238456 42708 238468
rect 42208 238428 42708 238456
rect 42208 238416 42214 238428
rect 42702 238416 42708 238428
rect 42760 238416 42766 238468
rect 52086 237396 52092 237448
rect 52144 237436 52150 237448
rect 184934 237436 184940 237448
rect 52144 237408 184940 237436
rect 52144 237396 52150 237408
rect 184934 237396 184940 237408
rect 184992 237396 184998 237448
rect 674466 236852 674472 236904
rect 674524 236892 674530 236904
rect 675386 236892 675392 236904
rect 674524 236864 675392 236892
rect 674524 236852 674530 236864
rect 675386 236852 675392 236864
rect 675444 236852 675450 236904
rect 42150 236648 42156 236700
rect 42208 236688 42214 236700
rect 42886 236688 42892 236700
rect 42208 236660 42892 236688
rect 42208 236648 42214 236660
rect 42886 236648 42892 236660
rect 42944 236648 42950 236700
rect 674742 235560 674748 235612
rect 674800 235600 674806 235612
rect 675662 235600 675668 235612
rect 674800 235572 675668 235600
rect 674800 235560 674806 235572
rect 675662 235560 675668 235572
rect 675720 235560 675726 235612
rect 674650 235492 674656 235544
rect 674708 235532 674714 235544
rect 675754 235532 675760 235544
rect 674708 235504 675760 235532
rect 674708 235492 674714 235504
rect 675754 235492 675760 235504
rect 675812 235492 675818 235544
rect 42150 235356 42156 235408
rect 42208 235396 42214 235408
rect 42794 235396 42800 235408
rect 42208 235368 42800 235396
rect 42208 235356 42214 235368
rect 42794 235356 42800 235368
rect 42852 235356 42858 235408
rect 42150 234608 42156 234660
rect 42208 234648 42214 234660
rect 43254 234648 43260 234660
rect 42208 234620 43260 234648
rect 42208 234608 42214 234620
rect 43254 234608 43260 234620
rect 43312 234608 43318 234660
rect 42150 234200 42156 234252
rect 42208 234240 42214 234252
rect 43162 234240 43168 234252
rect 42208 234212 43168 234240
rect 42208 234200 42214 234212
rect 43162 234200 43168 234212
rect 43220 234200 43226 234252
rect 42150 233316 42156 233368
rect 42208 233356 42214 233368
rect 43714 233356 43720 233368
rect 42208 233328 43720 233356
rect 42208 233316 42214 233328
rect 43714 233316 43720 233328
rect 43772 233316 43778 233368
rect 42150 231072 42156 231124
rect 42208 231112 42214 231124
rect 43622 231112 43628 231124
rect 42208 231084 43628 231112
rect 42208 231072 42214 231084
rect 43622 231072 43628 231084
rect 43680 231072 43686 231124
rect 48866 231072 48872 231124
rect 48924 231112 48930 231124
rect 654134 231112 654140 231124
rect 48924 231084 654140 231112
rect 48924 231072 48930 231084
rect 654134 231072 654140 231084
rect 654192 231072 654198 231124
rect 48958 231004 48964 231056
rect 49016 231044 49022 231056
rect 656986 231044 656992 231056
rect 49016 231016 656992 231044
rect 49016 231004 49022 231016
rect 656986 231004 656992 231016
rect 657044 231004 657050 231056
rect 46658 230936 46664 230988
rect 46716 230976 46722 230988
rect 656894 230976 656900 230988
rect 46716 230948 656900 230976
rect 46716 230936 46722 230948
rect 656894 230936 656900 230948
rect 656952 230936 656958 230988
rect 46842 230868 46848 230920
rect 46900 230908 46906 230920
rect 659746 230908 659752 230920
rect 46900 230880 659752 230908
rect 46900 230868 46906 230880
rect 659746 230868 659752 230880
rect 659804 230868 659810 230920
rect 46198 230800 46204 230852
rect 46256 230840 46262 230852
rect 659654 230840 659660 230852
rect 46256 230812 659660 230840
rect 46256 230800 46262 230812
rect 659654 230800 659660 230812
rect 659712 230800 659718 230852
rect 46382 230732 46388 230784
rect 46440 230772 46446 230784
rect 662690 230772 662696 230784
rect 46440 230744 662696 230772
rect 46440 230732 46446 230744
rect 662690 230732 662696 230744
rect 662748 230732 662754 230784
rect 46106 230664 46112 230716
rect 46164 230704 46170 230716
rect 662414 230704 662420 230716
rect 46164 230676 662420 230704
rect 46164 230664 46170 230676
rect 662414 230664 662420 230676
rect 662472 230664 662478 230716
rect 45922 230596 45928 230648
rect 45980 230636 45986 230648
rect 662506 230636 662512 230648
rect 45980 230608 662512 230636
rect 45980 230596 45986 230608
rect 662506 230596 662512 230608
rect 662564 230596 662570 230648
rect 42150 230528 42156 230580
rect 42208 230568 42214 230580
rect 43070 230568 43076 230580
rect 42208 230540 43076 230568
rect 42208 230528 42214 230540
rect 43070 230528 43076 230540
rect 43128 230528 43134 230580
rect 45830 230528 45836 230580
rect 45888 230568 45894 230580
rect 662598 230568 662604 230580
rect 45888 230540 662604 230568
rect 45888 230528 45894 230540
rect 662598 230528 662604 230540
rect 662656 230528 662662 230580
rect 45738 230460 45744 230512
rect 45796 230500 45802 230512
rect 662782 230500 662788 230512
rect 45796 230472 662788 230500
rect 45796 230460 45802 230472
rect 662782 230460 662788 230472
rect 662840 230460 662846 230512
rect 45370 230392 45376 230444
rect 45428 230432 45434 230444
rect 662874 230432 662880 230444
rect 45428 230404 662880 230432
rect 45428 230392 45434 230404
rect 662874 230392 662880 230404
rect 662932 230392 662938 230444
rect 350166 230256 350172 230308
rect 350224 230296 350230 230308
rect 423858 230296 423864 230308
rect 350224 230268 423864 230296
rect 350224 230256 350230 230268
rect 423858 230256 423864 230268
rect 423916 230256 423922 230308
rect 351638 230188 351644 230240
rect 351696 230228 351702 230240
rect 427170 230228 427176 230240
rect 351696 230200 427176 230228
rect 351696 230188 351702 230200
rect 427170 230188 427176 230200
rect 427228 230188 427234 230240
rect 348786 230120 348792 230172
rect 348844 230160 348850 230172
rect 420454 230160 420460 230172
rect 348844 230132 420460 230160
rect 348844 230120 348850 230132
rect 420454 230120 420460 230132
rect 420512 230120 420518 230172
rect 347314 230052 347320 230104
rect 347372 230092 347378 230104
rect 417142 230092 417148 230104
rect 347372 230064 417148 230092
rect 347372 230052 347378 230064
rect 417142 230052 417148 230064
rect 417200 230052 417206 230104
rect 354490 229984 354496 230036
rect 354548 230024 354554 230036
rect 433886 230024 433892 230036
rect 354548 229996 433892 230024
rect 354548 229984 354554 229996
rect 433886 229984 433892 229996
rect 433944 229984 433950 230036
rect 355870 229916 355876 229968
rect 355928 229956 355934 229968
rect 437290 229956 437296 229968
rect 355928 229928 437296 229956
rect 355928 229916 355934 229928
rect 437290 229916 437296 229928
rect 437348 229916 437354 229968
rect 42150 229848 42156 229900
rect 42208 229888 42214 229900
rect 42978 229888 42984 229900
rect 42208 229860 42984 229888
rect 42208 229848 42214 229860
rect 42978 229848 42984 229860
rect 43036 229848 43042 229900
rect 357342 229848 357348 229900
rect 357400 229888 357406 229900
rect 440694 229888 440700 229900
rect 357400 229860 440700 229888
rect 357400 229848 357406 229860
rect 440694 229848 440700 229860
rect 440752 229848 440758 229900
rect 360194 229780 360200 229832
rect 360252 229820 360258 229832
rect 447410 229820 447416 229832
rect 360252 229792 447416 229820
rect 360252 229780 360258 229792
rect 447410 229780 447416 229792
rect 447468 229780 447474 229832
rect 364058 229712 364064 229764
rect 364116 229752 364122 229764
rect 455782 229752 455788 229764
rect 364116 229724 455788 229752
rect 364116 229712 364122 229724
rect 455782 229712 455788 229724
rect 455840 229712 455846 229764
rect 365530 229644 365536 229696
rect 365588 229684 365594 229696
rect 459186 229684 459192 229696
rect 365588 229656 459192 229684
rect 365588 229644 365594 229656
rect 459186 229644 459192 229656
rect 459244 229644 459250 229696
rect 368382 229576 368388 229628
rect 368440 229616 368446 229628
rect 465994 229616 466000 229628
rect 368440 229588 466000 229616
rect 368440 229576 368446 229588
rect 465994 229576 466000 229588
rect 466052 229576 466058 229628
rect 371602 229508 371608 229560
rect 371660 229548 371666 229560
rect 474274 229548 474280 229560
rect 371660 229520 474280 229548
rect 371660 229508 371666 229520
rect 474274 229508 474280 229520
rect 474332 229508 474338 229560
rect 370498 229440 370504 229492
rect 370556 229480 370562 229492
rect 473446 229480 473452 229492
rect 370556 229452 473452 229480
rect 370556 229440 370562 229452
rect 473446 229440 473452 229452
rect 473504 229440 473510 229492
rect 371234 229372 371240 229424
rect 371292 229412 371298 229424
rect 472618 229412 472624 229424
rect 371292 229384 472624 229412
rect 371292 229372 371298 229384
rect 472618 229372 472624 229384
rect 472676 229372 472682 229424
rect 374086 229304 374092 229356
rect 374144 229344 374150 229356
rect 479334 229344 479340 229356
rect 374144 229316 479340 229344
rect 374144 229304 374150 229316
rect 479334 229304 479340 229316
rect 479392 229304 479398 229356
rect 376202 229236 376208 229288
rect 376260 229276 376266 229288
rect 487154 229276 487160 229288
rect 376260 229248 487160 229276
rect 376260 229236 376266 229248
rect 487154 229236 487160 229248
rect 487212 229236 487218 229288
rect 393682 229168 393688 229220
rect 393740 229208 393746 229220
rect 528370 229208 528376 229220
rect 393740 229180 528376 229208
rect 393740 229168 393746 229180
rect 528370 229168 528376 229180
rect 528428 229168 528434 229220
rect 396902 229100 396908 229152
rect 396960 229140 396966 229152
rect 535546 229140 535552 229152
rect 396960 229112 535552 229140
rect 396960 229100 396966 229112
rect 535546 229100 535552 229112
rect 535604 229100 535610 229152
rect 42150 229032 42156 229084
rect 42208 229072 42214 229084
rect 43346 229072 43352 229084
rect 42208 229044 43352 229072
rect 42208 229032 42214 229044
rect 43346 229032 43352 229044
rect 43404 229032 43410 229084
rect 156138 229032 156144 229084
rect 156196 229072 156202 229084
rect 235350 229072 235356 229084
rect 156196 229044 235356 229072
rect 156196 229032 156202 229044
rect 235350 229032 235356 229044
rect 235408 229032 235414 229084
rect 247034 229032 247040 229084
rect 247092 229072 247098 229084
rect 273898 229072 273904 229084
rect 247092 229044 273904 229072
rect 247092 229032 247098 229044
rect 273898 229032 273904 229044
rect 273956 229032 273962 229084
rect 296346 229032 296352 229084
rect 296404 229072 296410 229084
rect 298462 229072 298468 229084
rect 296404 229044 298468 229072
rect 296404 229032 296410 229044
rect 298462 229032 298468 229044
rect 298520 229032 298526 229084
rect 304534 229032 304540 229084
rect 304592 229072 304598 229084
rect 316126 229072 316132 229084
rect 304592 229044 316132 229072
rect 304592 229032 304598 229044
rect 316126 229032 316132 229044
rect 316184 229032 316190 229084
rect 368014 229032 368020 229084
rect 368072 229072 368078 229084
rect 369762 229072 369768 229084
rect 368072 229044 369768 229072
rect 368072 229032 368078 229044
rect 369762 229032 369768 229044
rect 369820 229032 369826 229084
rect 386230 229032 386236 229084
rect 386288 229072 386294 229084
rect 460934 229072 460940 229084
rect 386288 229044 460940 229072
rect 386288 229032 386294 229044
rect 460934 229032 460940 229044
rect 460992 229032 460998 229084
rect 152826 228964 152832 229016
rect 152884 229004 152890 229016
rect 233970 229004 233976 229016
rect 152884 228976 233976 229004
rect 152884 228964 152890 228976
rect 233970 228964 233976 228976
rect 234028 228964 234034 229016
rect 239950 228964 239956 229016
rect 240008 229004 240014 229016
rect 265342 229004 265348 229016
rect 240008 228976 265348 229004
rect 240008 228964 240014 228976
rect 265342 228964 265348 228976
rect 265400 228964 265406 229016
rect 290734 228964 290740 229016
rect 290792 229004 290798 229016
rect 292390 229004 292396 229016
rect 290792 228976 292396 229004
rect 290792 228964 290798 228976
rect 292390 228964 292396 228976
rect 292448 228964 292454 229016
rect 293218 228964 293224 229016
rect 293276 229004 293282 229016
rect 294598 229004 294604 229016
rect 293276 228976 294604 229004
rect 293276 228964 293282 228976
rect 294598 228964 294604 228976
rect 294656 228964 294662 229016
rect 297450 228964 297456 229016
rect 297508 229004 297514 229016
rect 299382 229004 299388 229016
rect 297508 228976 299388 229004
rect 297508 228964 297514 228976
rect 299382 228964 299388 228976
rect 299440 228964 299446 229016
rect 304166 228964 304172 229016
rect 304224 229004 304230 229016
rect 314654 229004 314660 229016
rect 304224 228976 314660 229004
rect 304224 228964 304230 228976
rect 314654 228964 314660 228976
rect 314712 228964 314718 229016
rect 343450 228964 343456 229016
rect 343508 229004 343514 229016
rect 381078 229004 381084 229016
rect 343508 228976 381084 229004
rect 343508 228964 343514 228976
rect 381078 228964 381084 228976
rect 381136 228964 381142 229016
rect 395062 228964 395068 229016
rect 395120 229004 395126 229016
rect 477494 229004 477500 229016
rect 395120 228976 477500 229004
rect 395120 228964 395126 228976
rect 477494 228964 477500 228976
rect 477552 228964 477558 229016
rect 156966 228896 156972 228948
rect 157024 228936 157030 228948
rect 237190 228936 237196 228948
rect 157024 228908 237196 228936
rect 157024 228896 157030 228908
rect 237190 228896 237196 228908
rect 237248 228896 237254 228948
rect 239214 228896 239220 228948
rect 239272 228936 239278 228948
rect 266722 228936 266728 228948
rect 239272 228908 266728 228936
rect 239272 228896 239278 228908
rect 266722 228896 266728 228908
rect 266780 228896 266786 228948
rect 297818 228896 297824 228948
rect 297876 228936 297882 228948
rect 301866 228936 301872 228948
rect 297876 228908 301872 228936
rect 297876 228896 297882 228908
rect 301866 228896 301872 228908
rect 301924 228896 301930 228948
rect 305638 228896 305644 228948
rect 305696 228936 305702 228948
rect 317874 228936 317880 228948
rect 305696 228908 317880 228936
rect 305696 228896 305702 228908
rect 317874 228896 317880 228908
rect 317932 228896 317938 228948
rect 320266 228896 320272 228948
rect 320324 228936 320330 228948
rect 342162 228936 342168 228948
rect 320324 228908 342168 228936
rect 320324 228896 320330 228908
rect 342162 228896 342168 228908
rect 342220 228896 342226 228948
rect 342346 228896 342352 228948
rect 342404 228936 342410 228948
rect 383746 228936 383752 228948
rect 342404 228908 383752 228936
rect 342404 228896 342410 228908
rect 383746 228896 383752 228908
rect 383804 228896 383810 228948
rect 388714 228896 388720 228948
rect 388772 228936 388778 228948
rect 469858 228936 469864 228948
rect 388772 228908 469864 228936
rect 388772 228896 388778 228908
rect 469858 228896 469864 228908
rect 469916 228896 469922 228948
rect 150250 228828 150256 228880
rect 150308 228868 150314 228880
rect 234338 228868 234344 228880
rect 150308 228840 234344 228868
rect 150308 228828 150314 228840
rect 234338 228828 234344 228840
rect 234396 228828 234402 228880
rect 240686 228828 240692 228880
rect 240744 228868 240750 228880
rect 269574 228868 269580 228880
rect 240744 228840 269580 228868
rect 240744 228828 240750 228840
rect 269574 228828 269580 228840
rect 269632 228828 269638 228880
rect 308490 228828 308496 228880
rect 308548 228868 308554 228880
rect 324590 228868 324596 228880
rect 308548 228840 324596 228868
rect 308548 228828 308554 228840
rect 324590 228828 324596 228840
rect 324648 228828 324654 228880
rect 340598 228828 340604 228880
rect 340656 228868 340662 228880
rect 385218 228868 385224 228880
rect 340656 228840 385224 228868
rect 340656 228828 340662 228840
rect 385218 228828 385224 228840
rect 385276 228828 385282 228880
rect 392946 228828 392952 228880
rect 393004 228868 393010 228880
rect 474734 228868 474740 228880
rect 393004 228840 474740 228868
rect 393004 228828 393010 228840
rect 474734 228828 474740 228840
rect 474792 228828 474798 228880
rect 146018 228760 146024 228812
rect 146076 228800 146082 228812
rect 231118 228800 231124 228812
rect 146076 228772 231124 228800
rect 146076 228760 146082 228772
rect 231118 228760 231124 228772
rect 231176 228760 231182 228812
rect 245286 228760 245292 228812
rect 245344 228800 245350 228812
rect 273530 228800 273536 228812
rect 245344 228772 273536 228800
rect 245344 228760 245350 228772
rect 273530 228760 273536 228772
rect 273588 228760 273594 228812
rect 310606 228760 310612 228812
rect 310664 228800 310670 228812
rect 332134 228800 332140 228812
rect 310664 228772 332140 228800
rect 310664 228760 310670 228772
rect 332134 228760 332140 228772
rect 332192 228760 332198 228812
rect 340874 228760 340880 228812
rect 340932 228800 340938 228812
rect 383654 228800 383660 228812
rect 340932 228772 383660 228800
rect 340932 228760 340938 228772
rect 383654 228760 383660 228772
rect 383712 228760 383718 228812
rect 390830 228760 390836 228812
rect 390888 228800 390894 228812
rect 473262 228800 473268 228812
rect 390888 228772 473268 228800
rect 390888 228760 390894 228772
rect 473262 228760 473268 228772
rect 473320 228760 473326 228812
rect 151722 228692 151728 228744
rect 151780 228732 151786 228744
rect 234706 228732 234712 228744
rect 151780 228704 234712 228732
rect 151780 228692 151786 228704
rect 234706 228692 234712 228704
rect 234764 228692 234770 228744
rect 241974 228692 241980 228744
rect 242032 228732 242038 228744
rect 272150 228732 272156 228744
rect 242032 228704 272156 228732
rect 242032 228692 242038 228704
rect 272150 228692 272156 228704
rect 272208 228692 272214 228744
rect 298830 228692 298836 228744
rect 298888 228732 298894 228744
rect 302694 228732 302700 228744
rect 298888 228704 302700 228732
rect 298888 228692 298894 228704
rect 302694 228692 302700 228704
rect 302752 228692 302758 228744
rect 307386 228692 307392 228744
rect 307444 228732 307450 228744
rect 322934 228732 322940 228744
rect 307444 228704 322940 228732
rect 307444 228692 307450 228704
rect 322934 228692 322940 228704
rect 322992 228692 322998 228744
rect 336642 228692 336648 228744
rect 336700 228732 336706 228744
rect 380986 228732 380992 228744
rect 336700 228704 380992 228732
rect 336700 228692 336706 228704
rect 380986 228692 380992 228704
rect 381044 228692 381050 228744
rect 397270 228692 397276 228744
rect 397328 228732 397334 228744
rect 480254 228732 480260 228744
rect 397328 228704 480260 228732
rect 397328 228692 397334 228704
rect 480254 228692 480260 228704
rect 480312 228692 480318 228744
rect 143442 228624 143448 228676
rect 143500 228664 143506 228676
rect 231486 228664 231492 228676
rect 143500 228636 231492 228664
rect 143500 228624 143506 228636
rect 231486 228624 231492 228636
rect 231544 228624 231550 228676
rect 239858 228624 239864 228676
rect 239916 228664 239922 228676
rect 268194 228664 268200 228676
rect 239916 228636 268200 228664
rect 239916 228624 239922 228636
rect 268194 228624 268200 228636
rect 268252 228624 268258 228676
rect 306650 228624 306656 228676
rect 306708 228664 306714 228676
rect 323762 228664 323768 228676
rect 306708 228636 323768 228664
rect 306708 228624 306714 228636
rect 323762 228624 323768 228636
rect 323820 228624 323826 228676
rect 328822 228624 328828 228676
rect 328880 228664 328886 228676
rect 345382 228664 345388 228676
rect 328880 228636 345388 228664
rect 328880 228624 328886 228636
rect 345382 228624 345388 228636
rect 345440 228624 345446 228676
rect 376570 228624 376576 228676
rect 376628 228664 376634 228676
rect 465902 228664 465908 228676
rect 376628 228636 465908 228664
rect 376628 228624 376634 228636
rect 465902 228624 465908 228636
rect 465960 228624 465966 228676
rect 138474 228556 138480 228608
rect 138532 228596 138538 228608
rect 229002 228596 229008 228608
rect 138532 228568 229008 228596
rect 138532 228556 138538 228568
rect 229002 228556 229008 228568
rect 229060 228556 229066 228608
rect 240134 228556 240140 228608
rect 240192 228596 240198 228608
rect 271046 228596 271052 228608
rect 240192 228568 271052 228596
rect 240192 228556 240198 228568
rect 271046 228556 271052 228568
rect 271104 228556 271110 228608
rect 308122 228556 308128 228608
rect 308180 228596 308186 228608
rect 327074 228596 327080 228608
rect 308180 228568 327080 228596
rect 308180 228556 308186 228568
rect 327074 228556 327080 228568
rect 327132 228556 327138 228608
rect 337746 228556 337752 228608
rect 337804 228596 337810 228608
rect 383838 228596 383844 228608
rect 337804 228568 383844 228596
rect 337804 228556 337810 228568
rect 383838 228556 383844 228568
rect 383896 228556 383902 228608
rect 388346 228556 388352 228608
rect 388404 228596 388410 228608
rect 408310 228596 408316 228608
rect 388404 228568 408316 228596
rect 388404 228556 388410 228568
rect 408310 228556 408316 228568
rect 408368 228556 408374 228608
rect 410886 228556 410892 228608
rect 410944 228596 410950 228608
rect 411162 228596 411168 228608
rect 410944 228568 411168 228596
rect 410944 228556 410950 228568
rect 411162 228556 411168 228568
rect 411220 228556 411226 228608
rect 516226 228596 516232 228608
rect 417252 228568 516232 228596
rect 145190 228488 145196 228540
rect 145248 228528 145254 228540
rect 231854 228528 231860 228540
rect 145248 228500 231860 228528
rect 145248 228488 145254 228500
rect 231854 228488 231860 228500
rect 231912 228488 231918 228540
rect 238570 228488 238576 228540
rect 238628 228528 238634 228540
rect 270678 228528 270684 228540
rect 238628 228500 270684 228528
rect 238628 228488 238634 228500
rect 270678 228488 270684 228500
rect 270736 228488 270742 228540
rect 303522 228488 303528 228540
rect 303580 228528 303586 228540
rect 315298 228528 315304 228540
rect 303580 228500 315304 228528
rect 303580 228488 303586 228500
rect 315298 228488 315304 228500
rect 315356 228488 315362 228540
rect 317414 228488 317420 228540
rect 317472 228528 317478 228540
rect 338114 228528 338120 228540
rect 317472 228500 338120 228528
rect 317472 228488 317478 228500
rect 338114 228488 338120 228500
rect 338172 228488 338178 228540
rect 341978 228488 341984 228540
rect 342036 228528 342042 228540
rect 394602 228528 394608 228540
rect 342036 228500 394608 228528
rect 342036 228488 342042 228500
rect 394602 228488 394608 228500
rect 394660 228488 394666 228540
rect 409046 228488 409052 228540
rect 409104 228528 409110 228540
rect 417252 228528 417280 228568
rect 516226 228556 516232 228568
rect 516284 228556 516290 228608
rect 409104 228500 417280 228528
rect 409104 228488 409110 228500
rect 417326 228488 417332 228540
rect 417384 228528 417390 228540
rect 518894 228528 518900 228540
rect 417384 228500 518900 228528
rect 417384 228488 417390 228500
rect 518894 228488 518900 228500
rect 518952 228488 518958 228540
rect 136818 228420 136824 228472
rect 136876 228460 136882 228472
rect 228634 228460 228640 228472
rect 136876 228432 228640 228460
rect 136876 228420 136882 228432
rect 228634 228420 228640 228432
rect 228692 228420 228698 228472
rect 235258 228420 235264 228472
rect 235316 228460 235322 228472
rect 269298 228460 269304 228472
rect 235316 228432 269304 228460
rect 235316 228420 235322 228432
rect 269298 228420 269304 228432
rect 269356 228420 269362 228472
rect 306006 228420 306012 228472
rect 306064 228460 306070 228472
rect 319530 228460 319536 228472
rect 306064 228432 319536 228460
rect 306064 228420 306070 228432
rect 319530 228420 319536 228432
rect 319588 228420 319594 228472
rect 324866 228420 324872 228472
rect 324924 228460 324930 228472
rect 365806 228460 365812 228472
rect 324924 228432 365812 228460
rect 324924 228420 324930 228432
rect 365806 228420 365812 228432
rect 365864 228420 365870 228472
rect 380802 228420 380808 228472
rect 380860 228460 380866 228472
rect 497826 228460 497832 228472
rect 380860 228432 497832 228460
rect 380860 228420 380866 228432
rect 497826 228420 497832 228432
rect 497884 228420 497890 228472
rect 131758 228352 131764 228404
rect 131816 228392 131822 228404
rect 226150 228392 226156 228404
rect 131816 228364 226156 228392
rect 131816 228352 131822 228364
rect 226150 228352 226156 228364
rect 226208 228352 226214 228404
rect 227622 228352 227628 228404
rect 227680 228392 227686 228404
rect 267090 228392 267096 228404
rect 227680 228364 267096 228392
rect 227680 228352 227686 228364
rect 267090 228352 267096 228364
rect 267148 228352 267154 228404
rect 309502 228352 309508 228404
rect 309560 228392 309566 228404
rect 330478 228392 330484 228404
rect 309560 228364 330484 228392
rect 309560 228352 309566 228364
rect 330478 228352 330484 228364
rect 330536 228352 330542 228404
rect 338022 228352 338028 228404
rect 338080 228392 338086 228404
rect 378134 228392 378140 228404
rect 338080 228364 378140 228392
rect 338080 228352 338086 228364
rect 378134 228352 378140 228364
rect 378192 228352 378198 228404
rect 383378 228352 383384 228404
rect 383436 228392 383442 228404
rect 503714 228392 503720 228404
rect 383436 228364 503720 228392
rect 383436 228352 383442 228364
rect 503714 228352 503720 228364
rect 503772 228352 503778 228404
rect 125042 228284 125048 228336
rect 125100 228324 125106 228336
rect 223298 228324 223304 228336
rect 125100 228296 223304 228324
rect 125100 228284 125106 228296
rect 223298 228284 223304 228296
rect 223356 228284 223362 228336
rect 223482 228284 223488 228336
rect 223540 228324 223546 228336
rect 263870 228324 263876 228336
rect 223540 228296 263876 228324
rect 223540 228284 223546 228296
rect 263870 228284 263876 228296
rect 263928 228284 263934 228336
rect 307754 228284 307760 228336
rect 307812 228324 307818 228336
rect 325694 228324 325700 228336
rect 307812 228296 325700 228324
rect 307812 228284 307818 228296
rect 325694 228284 325700 228296
rect 325752 228284 325758 228336
rect 330570 228284 330576 228336
rect 330628 228324 330634 228336
rect 379238 228324 379244 228336
rect 330628 228296 379244 228324
rect 330628 228284 330634 228296
rect 379238 228284 379244 228296
rect 379296 228284 379302 228336
rect 385494 228284 385500 228336
rect 385552 228324 385558 228336
rect 508774 228324 508780 228336
rect 385552 228296 508780 228324
rect 385552 228284 385558 228296
rect 508774 228284 508780 228296
rect 508832 228284 508838 228336
rect 130102 228216 130108 228268
rect 130160 228256 130166 228268
rect 225782 228256 225788 228268
rect 130160 228228 225788 228256
rect 130160 228216 130166 228228
rect 225782 228216 225788 228228
rect 225840 228216 225846 228268
rect 229370 228216 229376 228268
rect 229428 228256 229434 228268
rect 267458 228256 267464 228268
rect 229428 228228 267464 228256
rect 229428 228216 229434 228228
rect 267458 228216 267464 228228
rect 267516 228216 267522 228268
rect 309226 228216 309232 228268
rect 309284 228256 309290 228268
rect 328822 228256 328828 228268
rect 309284 228228 328828 228256
rect 309284 228216 309290 228228
rect 328822 228216 328828 228228
rect 328880 228216 328886 228268
rect 333422 228216 333428 228268
rect 333480 228256 333486 228268
rect 385954 228256 385960 228268
rect 333480 228228 385960 228256
rect 333480 228216 333486 228228
rect 385954 228216 385960 228228
rect 386012 228216 386018 228268
rect 387610 228216 387616 228268
rect 387668 228256 387674 228268
rect 513834 228256 513840 228268
rect 387668 228228 513840 228256
rect 387668 228216 387674 228228
rect 513834 228216 513840 228228
rect 513892 228216 513898 228268
rect 123386 228148 123392 228200
rect 123444 228188 123450 228200
rect 222930 228188 222936 228200
rect 123444 228160 222936 228188
rect 123444 228148 123450 228160
rect 222930 228148 222936 228160
rect 222988 228148 222994 228200
rect 231670 228148 231676 228200
rect 231728 228188 231734 228200
rect 267826 228188 267832 228200
rect 231728 228160 267832 228188
rect 231728 228148 231734 228160
rect 267826 228148 267832 228160
rect 267884 228148 267890 228200
rect 300946 228148 300952 228200
rect 301004 228188 301010 228200
rect 310238 228188 310244 228200
rect 301004 228160 310244 228188
rect 301004 228148 301010 228160
rect 310238 228148 310244 228160
rect 310296 228148 310302 228200
rect 310514 228148 310520 228200
rect 310572 228188 310578 228200
rect 329650 228188 329656 228200
rect 310572 228160 329656 228188
rect 310572 228148 310578 228160
rect 329650 228148 329656 228160
rect 329708 228148 329714 228200
rect 339126 228148 339132 228200
rect 339184 228188 339190 228200
rect 391842 228188 391848 228200
rect 339184 228160 391848 228188
rect 339184 228148 339190 228160
rect 391842 228148 391848 228160
rect 391900 228148 391906 228200
rect 399386 228148 399392 228200
rect 399444 228188 399450 228200
rect 541618 228188 541624 228200
rect 399444 228160 541624 228188
rect 399444 228148 399450 228160
rect 541618 228148 541624 228160
rect 541676 228148 541682 228200
rect 108206 228080 108212 228132
rect 108264 228120 108270 228132
rect 216122 228120 216128 228132
rect 108264 228092 216128 228120
rect 108264 228080 108270 228092
rect 216122 228080 216128 228092
rect 216180 228080 216186 228132
rect 216674 228080 216680 228132
rect 216732 228120 216738 228132
rect 261018 228120 261024 228132
rect 216732 228092 261024 228120
rect 216732 228080 216738 228092
rect 261018 228080 261024 228092
rect 261076 228080 261082 228132
rect 308858 228080 308864 228132
rect 308916 228120 308922 228132
rect 326246 228120 326252 228132
rect 308916 228092 326252 228120
rect 308916 228080 308922 228092
rect 326246 228080 326252 228092
rect 326304 228080 326310 228132
rect 334894 228080 334900 228132
rect 334952 228120 334958 228132
rect 389082 228120 389088 228132
rect 334952 228092 389088 228120
rect 334952 228080 334958 228092
rect 389082 228080 389088 228092
rect 389140 228080 389146 228132
rect 407206 228080 407212 228132
rect 407264 228120 407270 228132
rect 417326 228120 417332 228132
rect 407264 228092 417332 228120
rect 407264 228080 407270 228092
rect 417326 228080 417332 228092
rect 417384 228080 417390 228132
rect 544102 228120 544108 228132
rect 417436 228092 544108 228120
rect 78766 228012 78772 228064
rect 78824 228052 78830 228064
rect 202598 228052 202604 228064
rect 78824 228024 202604 228052
rect 78824 228012 78830 228024
rect 202598 228012 202604 228024
rect 202656 228012 202662 228064
rect 209682 228012 209688 228064
rect 209740 228052 209746 228064
rect 258166 228052 258172 228064
rect 209740 228024 258172 228052
rect 209740 228012 209746 228024
rect 258166 228012 258172 228024
rect 258224 228012 258230 228064
rect 259362 228012 259368 228064
rect 259420 228052 259426 228064
rect 276014 228052 276020 228064
rect 259420 228024 276020 228052
rect 259420 228012 259426 228024
rect 276014 228012 276020 228024
rect 276072 228012 276078 228064
rect 311710 228012 311716 228064
rect 311768 228052 311774 228064
rect 332962 228052 332968 228064
rect 311768 228024 332968 228052
rect 311768 228012 311774 228024
rect 332962 228012 332968 228024
rect 333020 228012 333026 228064
rect 336274 228012 336280 228064
rect 336332 228052 336338 228064
rect 388990 228052 388996 228064
rect 336332 228024 388996 228052
rect 336332 228012 336338 228024
rect 388990 228012 388996 228024
rect 389048 228012 389054 228064
rect 400490 228012 400496 228064
rect 400548 228052 400554 228064
rect 417436 228052 417464 228092
rect 544102 228080 544108 228092
rect 544160 228080 544166 228132
rect 400548 228024 417464 228052
rect 400548 228012 400554 228024
rect 417510 228012 417516 228064
rect 417568 228052 417574 228064
rect 545206 228052 545212 228064
rect 417568 228024 545212 228052
rect 417568 228012 417574 228024
rect 545206 228012 545212 228024
rect 545264 228012 545270 228064
rect 65334 227944 65340 227996
rect 65392 227984 65398 227996
rect 196894 227984 196900 227996
rect 65392 227956 196900 227984
rect 65392 227944 65398 227956
rect 196894 227944 196900 227956
rect 196952 227944 196958 227996
rect 199010 227944 199016 227996
rect 199068 227984 199074 227996
rect 254302 227984 254308 227996
rect 199068 227956 254308 227984
rect 199068 227944 199074 227956
rect 254302 227944 254308 227956
rect 254360 227944 254366 227996
rect 254394 227944 254400 227996
rect 254452 227984 254458 227996
rect 275646 227984 275652 227996
rect 254452 227956 275652 227984
rect 254452 227944 254458 227956
rect 275646 227944 275652 227956
rect 275704 227944 275710 227996
rect 302786 227944 302792 227996
rect 302844 227984 302850 227996
rect 311158 227984 311164 227996
rect 302844 227956 311164 227984
rect 302844 227944 302850 227956
rect 311158 227944 311164 227956
rect 311216 227944 311222 227996
rect 311342 227944 311348 227996
rect 311400 227984 311406 227996
rect 331306 227984 331312 227996
rect 311400 227956 331312 227984
rect 311400 227944 311406 227956
rect 331306 227944 331312 227956
rect 331364 227944 331370 227996
rect 342714 227944 342720 227996
rect 342772 227984 342778 227996
rect 395154 227984 395160 227996
rect 342772 227956 395160 227984
rect 342772 227944 342778 227956
rect 395154 227944 395160 227956
rect 395212 227944 395218 227996
rect 402606 227944 402612 227996
rect 402664 227984 402670 227996
rect 549254 227984 549260 227996
rect 402664 227956 549260 227984
rect 402664 227944 402670 227956
rect 549254 227944 549260 227956
rect 549312 227944 549318 227996
rect 77938 227876 77944 227928
rect 77996 227916 78002 227928
rect 203058 227916 203064 227928
rect 77996 227888 203064 227916
rect 77996 227876 78002 227888
rect 203058 227876 203064 227888
rect 203116 227876 203122 227928
rect 203242 227876 203248 227928
rect 203300 227916 203306 227928
rect 255314 227916 255320 227928
rect 203300 227888 255320 227916
rect 203300 227876 203306 227888
rect 255314 227876 255320 227888
rect 255372 227876 255378 227928
rect 257246 227876 257252 227928
rect 257304 227916 257310 227928
rect 277486 227916 277492 227928
rect 257304 227888 277492 227916
rect 257304 227876 257310 227888
rect 277486 227876 277492 227888
rect 277544 227876 277550 227928
rect 301682 227876 301688 227928
rect 301740 227916 301746 227928
rect 309410 227916 309416 227928
rect 301740 227888 309416 227916
rect 301740 227876 301746 227888
rect 309410 227876 309416 227888
rect 309468 227876 309474 227928
rect 312722 227876 312728 227928
rect 312780 227916 312786 227928
rect 334710 227916 334716 227928
rect 312780 227888 334716 227916
rect 312780 227876 312786 227888
rect 334710 227876 334716 227888
rect 334768 227876 334774 227928
rect 338390 227876 338396 227928
rect 338448 227916 338454 227928
rect 395246 227916 395252 227928
rect 338448 227888 395252 227916
rect 338448 227876 338454 227888
rect 395246 227876 395252 227888
rect 395304 227876 395310 227928
rect 404722 227876 404728 227928
rect 404780 227916 404786 227928
rect 554222 227916 554228 227928
rect 404780 227888 554228 227916
rect 404780 227876 404786 227888
rect 554222 227876 554228 227888
rect 554280 227876 554286 227928
rect 72050 227808 72056 227860
rect 72108 227848 72114 227860
rect 199746 227848 199752 227860
rect 72108 227820 199752 227848
rect 72108 227808 72114 227820
rect 199746 227808 199752 227820
rect 199804 227808 199810 227860
rect 204070 227808 204076 227860
rect 204128 227848 204134 227860
rect 257154 227848 257160 227860
rect 204128 227820 257160 227848
rect 204128 227808 204134 227820
rect 257154 227808 257160 227820
rect 257212 227808 257218 227860
rect 261478 227808 261484 227860
rect 261536 227848 261542 227860
rect 278866 227848 278872 227860
rect 261536 227820 278872 227848
rect 261536 227808 261542 227820
rect 278866 227808 278872 227820
rect 278924 227808 278930 227860
rect 303798 227808 303804 227860
rect 303856 227848 303862 227860
rect 317414 227848 317420 227860
rect 303856 227820 317420 227848
rect 303856 227808 303862 227820
rect 317414 227808 317420 227820
rect 317472 227808 317478 227860
rect 318794 227808 318800 227860
rect 318852 227848 318858 227860
rect 318852 227820 322934 227848
rect 318852 227808 318858 227820
rect 64506 227740 64512 227792
rect 64564 227780 64570 227792
rect 197630 227780 197636 227792
rect 64564 227752 197636 227780
rect 64564 227740 64570 227752
rect 197630 227740 197636 227752
rect 197688 227740 197694 227792
rect 197722 227740 197728 227792
rect 197780 227780 197786 227792
rect 254026 227780 254032 227792
rect 197780 227752 254032 227780
rect 197780 227740 197786 227752
rect 254026 227740 254032 227752
rect 254084 227740 254090 227792
rect 254210 227740 254216 227792
rect 254268 227780 254274 227792
rect 277118 227780 277124 227792
rect 254268 227752 277124 227780
rect 254268 227740 254274 227752
rect 277118 227740 277124 227752
rect 277176 227740 277182 227792
rect 304902 227740 304908 227792
rect 304960 227780 304966 227792
rect 318702 227780 318708 227792
rect 304960 227752 318708 227780
rect 304960 227740 304966 227752
rect 318702 227740 318708 227752
rect 318760 227740 318766 227792
rect 322906 227780 322934 227820
rect 341242 227808 341248 227860
rect 341300 227848 341306 227860
rect 397638 227848 397644 227860
rect 341300 227820 397644 227848
rect 341300 227808 341306 227820
rect 397638 227808 397644 227820
rect 397696 227808 397702 227860
rect 406838 227808 406844 227860
rect 406896 227848 406902 227860
rect 559282 227848 559288 227860
rect 406896 227820 559288 227848
rect 406896 227808 406902 227820
rect 559282 227808 559288 227820
rect 559340 227808 559346 227860
rect 339770 227780 339776 227792
rect 322906 227752 339776 227780
rect 339770 227740 339776 227752
rect 339828 227740 339834 227792
rect 345934 227740 345940 227792
rect 345992 227780 345998 227792
rect 408218 227780 408224 227792
rect 345992 227752 408224 227780
rect 345992 227740 345998 227752
rect 408218 227740 408224 227752
rect 408276 227740 408282 227792
rect 409322 227740 409328 227792
rect 409380 227780 409386 227792
rect 565446 227780 565452 227792
rect 409380 227752 565452 227780
rect 409380 227740 409386 227752
rect 565446 227740 565452 227752
rect 565504 227740 565510 227792
rect 52730 227672 52736 227724
rect 52788 227712 52794 227724
rect 192938 227712 192944 227724
rect 52788 227684 192944 227712
rect 52788 227672 52794 227684
rect 192938 227672 192944 227684
rect 192996 227672 193002 227724
rect 193030 227672 193036 227724
rect 193088 227712 193094 227724
rect 251818 227712 251824 227724
rect 193088 227684 251824 227712
rect 193088 227672 193094 227684
rect 251818 227672 251824 227684
rect 251876 227672 251882 227724
rect 252002 227672 252008 227724
rect 252060 227712 252066 227724
rect 276382 227712 276388 227724
rect 252060 227684 276388 227712
rect 252060 227672 252066 227684
rect 276382 227672 276388 227684
rect 276440 227672 276446 227724
rect 312078 227672 312084 227724
rect 312136 227712 312142 227724
rect 335538 227712 335544 227724
rect 312136 227684 335544 227712
rect 312136 227672 312142 227684
rect 335538 227672 335544 227684
rect 335596 227672 335602 227724
rect 341610 227672 341616 227724
rect 341668 227712 341674 227724
rect 402146 227712 402152 227724
rect 341668 227684 402152 227712
rect 341668 227672 341674 227684
rect 402146 227672 402152 227684
rect 402204 227672 402210 227724
rect 410426 227672 410432 227724
rect 410484 227712 410490 227724
rect 567930 227712 567936 227724
rect 410484 227684 567936 227712
rect 410484 227672 410490 227684
rect 567930 227672 567936 227684
rect 567988 227672 567994 227724
rect 158714 227604 158720 227656
rect 158772 227644 158778 227656
rect 237558 227644 237564 227656
rect 158772 227616 237564 227644
rect 158772 227604 158778 227616
rect 237558 227604 237564 227616
rect 237616 227604 237622 227656
rect 243630 227604 243636 227656
rect 243688 227644 243694 227656
rect 272426 227644 272432 227656
rect 243688 227616 272432 227644
rect 243688 227604 243694 227616
rect 272426 227604 272432 227616
rect 272484 227604 272490 227656
rect 305270 227604 305276 227656
rect 305328 227644 305334 227656
rect 320358 227644 320364 227656
rect 305328 227616 320364 227644
rect 305328 227604 305334 227616
rect 320358 227604 320364 227616
rect 320416 227604 320422 227656
rect 320634 227604 320640 227656
rect 320692 227644 320698 227656
rect 320692 227616 322934 227644
rect 320692 227604 320698 227616
rect 165430 227536 165436 227588
rect 165488 227576 165494 227588
rect 240410 227576 240416 227588
rect 165488 227548 240416 227576
rect 165488 227536 165494 227548
rect 240410 227536 240416 227548
rect 240468 227536 240474 227588
rect 250346 227536 250352 227588
rect 250404 227576 250410 227588
rect 275278 227576 275284 227588
rect 250404 227548 275284 227576
rect 250404 227536 250410 227548
rect 275278 227536 275284 227548
rect 275336 227536 275342 227588
rect 307018 227536 307024 227588
rect 307076 227576 307082 227588
rect 321186 227576 321192 227588
rect 307076 227548 321192 227576
rect 307076 227536 307082 227548
rect 321186 227536 321192 227548
rect 321244 227536 321250 227588
rect 322906 227576 322934 227616
rect 332042 227604 332048 227656
rect 332100 227644 332106 227656
rect 369670 227644 369676 227656
rect 332100 227616 369676 227644
rect 332100 227604 332106 227616
rect 369670 227604 369676 227616
rect 369728 227604 369734 227656
rect 381906 227604 381912 227656
rect 381964 227644 381970 227656
rect 453666 227644 453672 227656
rect 381964 227616 453672 227644
rect 381964 227604 381970 227616
rect 453666 227604 453672 227616
rect 453724 227604 453730 227656
rect 356054 227576 356060 227588
rect 322906 227548 356060 227576
rect 356054 227536 356060 227548
rect 356112 227536 356118 227588
rect 356606 227536 356612 227588
rect 356664 227576 356670 227588
rect 372890 227576 372896 227588
rect 356664 227548 372896 227576
rect 356664 227536 356670 227548
rect 372890 227536 372896 227548
rect 372948 227536 372954 227588
rect 384022 227536 384028 227588
rect 384080 227576 384086 227588
rect 455414 227576 455420 227588
rect 384080 227548 455420 227576
rect 384080 227536 384086 227548
rect 455414 227536 455420 227548
rect 455472 227536 455478 227588
rect 162762 227468 162768 227520
rect 162820 227508 162826 227520
rect 238202 227508 238208 227520
rect 162820 227480 238208 227508
rect 162820 227468 162826 227480
rect 238202 227468 238208 227480
rect 238260 227468 238266 227520
rect 253658 227468 253664 227520
rect 253716 227508 253722 227520
rect 276750 227508 276756 227520
rect 253716 227480 276756 227508
rect 253716 227468 253722 227480
rect 276750 227468 276756 227480
rect 276808 227468 276814 227520
rect 303154 227468 303160 227520
rect 303212 227508 303218 227520
rect 312814 227508 312820 227520
rect 303212 227480 312820 227508
rect 303212 227468 303218 227480
rect 312814 227468 312820 227480
rect 312872 227468 312878 227520
rect 324498 227468 324504 227520
rect 324556 227508 324562 227520
rect 345290 227508 345296 227520
rect 324556 227480 345296 227508
rect 324556 227468 324562 227480
rect 345290 227468 345296 227480
rect 345348 227468 345354 227520
rect 353018 227468 353024 227520
rect 353076 227508 353082 227520
rect 410978 227508 410984 227520
rect 353076 227480 410984 227508
rect 353076 227468 353082 227480
rect 410978 227468 410984 227480
rect 411036 227468 411042 227520
rect 42058 227400 42064 227452
rect 42116 227440 42122 227452
rect 43530 227440 43536 227452
rect 42116 227412 43536 227440
rect 42116 227400 42122 227412
rect 43530 227400 43536 227412
rect 43588 227400 43594 227452
rect 163682 227400 163688 227452
rect 163740 227440 163746 227452
rect 240042 227440 240048 227452
rect 163740 227412 240048 227440
rect 163740 227400 163746 227412
rect 240042 227400 240048 227412
rect 240100 227400 240106 227452
rect 257338 227400 257344 227452
rect 257396 227440 257402 227452
rect 264606 227440 264612 227452
rect 257396 227412 264612 227440
rect 257396 227400 257402 227412
rect 264606 227400 264612 227412
rect 264664 227400 264670 227452
rect 264698 227400 264704 227452
rect 264756 227440 264762 227452
rect 275002 227440 275008 227452
rect 264756 227412 275008 227440
rect 264756 227400 264762 227412
rect 275002 227400 275008 227412
rect 275060 227400 275066 227452
rect 325970 227400 325976 227452
rect 326028 227440 326034 227452
rect 345106 227440 345112 227452
rect 326028 227412 345112 227440
rect 326028 227400 326034 227412
rect 345106 227400 345112 227412
rect 345164 227400 345170 227452
rect 372982 227400 372988 227452
rect 373040 227440 373046 227452
rect 433150 227440 433156 227452
rect 373040 227412 433156 227440
rect 373040 227400 373046 227412
rect 433150 227400 433156 227412
rect 433208 227400 433214 227452
rect 167086 227332 167092 227384
rect 167144 227372 167150 227384
rect 241422 227372 241428 227384
rect 167144 227344 241428 227372
rect 167144 227332 167150 227344
rect 241422 227332 241428 227344
rect 241480 227332 241486 227384
rect 251266 227332 251272 227384
rect 251324 227372 251330 227384
rect 271414 227372 271420 227384
rect 251324 227344 271420 227372
rect 251324 227332 251330 227344
rect 271414 227332 271420 227344
rect 271472 227332 271478 227384
rect 323118 227332 323124 227384
rect 323176 227372 323182 227384
rect 342806 227372 342812 227384
rect 323176 227344 342812 227372
rect 323176 227332 323182 227344
rect 342806 227332 342812 227344
rect 342864 227332 342870 227384
rect 358722 227332 358728 227384
rect 358780 227372 358786 227384
rect 415302 227372 415308 227384
rect 358780 227344 415308 227372
rect 358780 227332 358786 227344
rect 415302 227332 415308 227344
rect 415360 227332 415366 227384
rect 172146 227264 172152 227316
rect 172204 227304 172210 227316
rect 243262 227304 243268 227316
rect 172204 227276 243268 227304
rect 172204 227264 172210 227276
rect 243262 227264 243268 227276
rect 243320 227264 243326 227316
rect 248506 227264 248512 227316
rect 248564 227304 248570 227316
rect 268562 227304 268568 227316
rect 248564 227276 268568 227304
rect 248564 227264 248570 227276
rect 268562 227264 268568 227276
rect 268620 227264 268626 227316
rect 295242 227264 295248 227316
rect 295300 227304 295306 227316
rect 296806 227304 296812 227316
rect 295300 227276 296812 227304
rect 295300 227264 295306 227276
rect 296806 227264 296812 227276
rect 296864 227264 296870 227316
rect 298738 227264 298744 227316
rect 298796 227304 298802 227316
rect 301038 227304 301044 227316
rect 298796 227276 301044 227304
rect 298796 227264 298802 227276
rect 301038 227264 301044 227276
rect 301096 227264 301102 227316
rect 302418 227264 302424 227316
rect 302476 227304 302482 227316
rect 313642 227304 313648 227316
rect 302476 227276 313648 227304
rect 302476 227264 302482 227276
rect 313642 227264 313648 227276
rect 313700 227264 313706 227316
rect 374822 227264 374828 227316
rect 374880 227304 374886 227316
rect 433242 227304 433248 227316
rect 374880 227276 433248 227304
rect 374880 227264 374886 227276
rect 433242 227264 433248 227276
rect 433300 227264 433306 227316
rect 169570 227196 169576 227248
rect 169628 227236 169634 227248
rect 241054 227236 241060 227248
rect 169628 227208 241060 227236
rect 169628 227196 169634 227208
rect 241054 227196 241060 227208
rect 241112 227196 241118 227248
rect 251174 227196 251180 227248
rect 251232 227236 251238 227248
rect 272794 227236 272800 227248
rect 251232 227208 272800 227236
rect 251232 227196 251238 227208
rect 272794 227196 272800 227208
rect 272852 227196 272858 227248
rect 302050 227196 302056 227248
rect 302108 227236 302114 227248
rect 311986 227236 311992 227248
rect 302108 227208 311992 227236
rect 302108 227196 302114 227208
rect 311986 227196 311992 227208
rect 312044 227196 312050 227248
rect 370130 227196 370136 227248
rect 370188 227236 370194 227248
rect 428366 227236 428372 227248
rect 370188 227208 428372 227236
rect 370188 227196 370194 227208
rect 428366 227196 428372 227208
rect 428424 227196 428430 227248
rect 173618 227128 173624 227180
rect 173676 227168 173682 227180
rect 244274 227168 244280 227180
rect 173676 227140 244280 227168
rect 173676 227128 173682 227140
rect 244274 227128 244280 227140
rect 244332 227128 244338 227180
rect 248598 227128 248604 227180
rect 248656 227168 248662 227180
rect 269942 227168 269948 227180
rect 248656 227140 269948 227168
rect 248656 227128 248662 227140
rect 269942 227128 269948 227140
rect 270000 227128 270006 227180
rect 333054 227128 333060 227180
rect 333112 227168 333118 227180
rect 347774 227168 347780 227180
rect 333112 227140 347780 227168
rect 333112 227128 333118 227140
rect 347774 227128 347780 227140
rect 347832 227128 347838 227180
rect 367278 227128 367284 227180
rect 367336 227168 367342 227180
rect 422294 227168 422300 227180
rect 367336 227140 422300 227168
rect 367336 227128 367342 227140
rect 422294 227128 422300 227140
rect 422352 227128 422358 227180
rect 178862 227060 178868 227112
rect 178920 227100 178926 227112
rect 246114 227100 246120 227112
rect 178920 227072 246120 227100
rect 178920 227060 178926 227072
rect 246114 227060 246120 227072
rect 246172 227060 246178 227112
rect 254118 227060 254124 227112
rect 254176 227100 254182 227112
rect 274266 227100 274272 227112
rect 254176 227072 274272 227100
rect 254176 227060 254182 227072
rect 274266 227060 274272 227072
rect 274324 227060 274330 227112
rect 331674 227060 331680 227112
rect 331732 227100 331738 227112
rect 347866 227100 347872 227112
rect 331732 227072 347872 227100
rect 331732 227060 331738 227072
rect 347866 227060 347872 227072
rect 347924 227060 347930 227112
rect 364426 227060 364432 227112
rect 364484 227100 364490 227112
rect 416774 227100 416780 227112
rect 364484 227072 416780 227100
rect 364484 227060 364490 227072
rect 416774 227060 416780 227072
rect 416832 227060 416838 227112
rect 176378 226992 176384 227044
rect 176436 227032 176442 227044
rect 243906 227032 243912 227044
rect 176436 227004 243912 227032
rect 176436 226992 176442 227004
rect 243906 226992 243912 227004
rect 243964 226992 243970 227044
rect 248414 226992 248420 227044
rect 248472 227032 248478 227044
rect 265710 227032 265716 227044
rect 248472 227004 265716 227032
rect 248472 226992 248478 227004
rect 265710 226992 265716 227004
rect 265768 226992 265774 227044
rect 322014 226992 322020 227044
rect 322072 227032 322078 227044
rect 359090 227032 359096 227044
rect 322072 227004 359096 227032
rect 322072 226992 322078 227004
rect 359090 226992 359096 227004
rect 359148 226992 359154 227044
rect 361574 226992 361580 227044
rect 361632 227032 361638 227044
rect 415486 227032 415492 227044
rect 361632 227004 415492 227032
rect 361632 226992 361638 227004
rect 415486 226992 415492 227004
rect 415544 226992 415550 227044
rect 180518 226924 180524 226976
rect 180576 226964 180582 226976
rect 247126 226964 247132 226976
rect 180576 226936 247132 226964
rect 180576 226924 180582 226936
rect 247126 226924 247132 226936
rect 247184 226924 247190 226976
rect 254302 226924 254308 226976
rect 254360 226964 254366 226976
rect 271782 226964 271788 226976
rect 254360 226936 271788 226964
rect 254360 226924 254366 226936
rect 271782 226924 271788 226936
rect 271840 226924 271846 226976
rect 345198 226924 345204 226976
rect 345256 226964 345262 226976
rect 376662 226964 376668 226976
rect 345256 226936 376668 226964
rect 345256 226924 345262 226936
rect 376662 226924 376668 226936
rect 376720 226924 376726 226976
rect 379054 226924 379060 226976
rect 379112 226964 379118 226976
rect 387518 226964 387524 226976
rect 379112 226936 387524 226964
rect 379112 226924 379118 226936
rect 387518 226924 387524 226936
rect 387576 226924 387582 226976
rect 399018 226924 399024 226976
rect 399076 226964 399082 226976
rect 438854 226964 438860 226976
rect 399076 226936 438860 226964
rect 399076 226924 399082 226936
rect 438854 226924 438860 226936
rect 438912 226924 438918 226976
rect 190362 226856 190368 226908
rect 190420 226896 190426 226908
rect 251450 226896 251456 226908
rect 190420 226868 251456 226896
rect 190420 226856 190426 226868
rect 251450 226856 251456 226868
rect 251508 226856 251514 226908
rect 257798 226856 257804 226908
rect 257856 226896 257862 226908
rect 274634 226896 274640 226908
rect 257856 226868 274640 226896
rect 257856 226856 257862 226868
rect 274634 226856 274640 226868
rect 274692 226856 274698 226908
rect 300670 226856 300676 226908
rect 300728 226896 300734 226908
rect 308582 226896 308588 226908
rect 300728 226868 308588 226896
rect 300728 226856 300734 226868
rect 308582 226856 308588 226868
rect 308640 226856 308646 226908
rect 359826 226856 359832 226908
rect 359884 226896 359890 226908
rect 400214 226896 400220 226908
rect 359884 226868 400220 226896
rect 359884 226856 359890 226868
rect 400214 226856 400220 226868
rect 400272 226856 400278 226908
rect 400766 226856 400772 226908
rect 400824 226896 400830 226908
rect 417510 226896 417516 226908
rect 400824 226868 417516 226896
rect 400824 226856 400830 226868
rect 417510 226856 417516 226868
rect 417568 226856 417574 226908
rect 449618 226896 449624 226908
rect 417620 226868 449624 226896
rect 42150 226788 42156 226840
rect 42208 226828 42214 226840
rect 43898 226828 43904 226840
rect 42208 226800 43904 226828
rect 42208 226788 42214 226800
rect 43898 226788 43904 226800
rect 43956 226788 43962 226840
rect 185578 226788 185584 226840
rect 185636 226828 185642 226840
rect 185636 226800 234016 226828
rect 185636 226788 185642 226800
rect 186406 226720 186412 226772
rect 186464 226760 186470 226772
rect 233878 226760 233884 226772
rect 186464 226732 233884 226760
rect 186464 226720 186470 226732
rect 233878 226720 233884 226732
rect 233936 226720 233942 226772
rect 192938 226652 192944 226704
rect 192996 226692 193002 226704
rect 233988 226692 234016 226800
rect 234062 226788 234068 226840
rect 234120 226828 234126 226840
rect 248230 226828 248236 226840
rect 234120 226800 248236 226828
rect 234120 226788 234126 226800
rect 248230 226788 248236 226800
rect 248288 226788 248294 226840
rect 248690 226788 248696 226840
rect 248748 226828 248754 226840
rect 264698 226828 264704 226840
rect 248748 226800 264704 226828
rect 248748 226788 248754 226800
rect 264698 226788 264704 226800
rect 264756 226788 264762 226840
rect 299566 226788 299572 226840
rect 299624 226828 299630 226840
rect 306926 226828 306932 226840
rect 299624 226800 306932 226828
rect 299624 226788 299630 226800
rect 306926 226788 306932 226800
rect 306984 226788 306990 226840
rect 323486 226788 323492 226840
rect 323544 226828 323550 226840
rect 362402 226828 362408 226840
rect 323544 226800 362408 226828
rect 323544 226788 323550 226800
rect 362402 226788 362408 226800
rect 362460 226788 362466 226840
rect 363046 226788 363052 226840
rect 363104 226828 363110 226840
rect 371510 226828 371516 226840
rect 363104 226800 371516 226828
rect 363104 226788 363110 226800
rect 371510 226788 371516 226800
rect 371568 226788 371574 226840
rect 373350 226788 373356 226840
rect 373408 226828 373414 226840
rect 395982 226828 395988 226840
rect 373408 226800 395988 226828
rect 373408 226788 373414 226800
rect 395982 226788 395988 226800
rect 396040 226788 396046 226840
rect 407574 226788 407580 226840
rect 407632 226828 407638 226840
rect 417620 226828 417648 226868
rect 449618 226856 449624 226868
rect 449676 226856 449682 226908
rect 407632 226800 417648 226828
rect 407632 226788 407638 226800
rect 417694 226788 417700 226840
rect 417752 226828 417758 226840
rect 441614 226828 441620 226840
rect 417752 226800 441620 226828
rect 417752 226788 417758 226800
rect 441614 226788 441620 226800
rect 441672 226788 441678 226840
rect 258442 226720 258448 226772
rect 258500 226760 258506 226772
rect 273162 226760 273168 226772
rect 258500 226732 273168 226760
rect 258500 226720 258506 226732
rect 273162 226720 273168 226732
rect 273220 226720 273226 226772
rect 299198 226720 299204 226772
rect 299256 226760 299262 226772
rect 305270 226760 305276 226772
rect 299256 226732 305276 226760
rect 299256 226720 299262 226732
rect 305270 226720 305276 226732
rect 305328 226720 305334 226772
rect 306374 226720 306380 226772
rect 306432 226760 306438 226772
rect 322014 226760 322020 226772
rect 306432 226732 322020 226760
rect 306432 226720 306438 226732
rect 322014 226720 322020 226732
rect 322072 226720 322078 226772
rect 371970 226720 371976 226772
rect 372028 226760 372034 226772
rect 400398 226760 400404 226772
rect 372028 226732 400404 226760
rect 372028 226720 372034 226732
rect 400398 226720 400404 226732
rect 400456 226720 400462 226772
rect 405458 226720 405464 226772
rect 405516 226760 405522 226772
rect 444558 226760 444564 226772
rect 405516 226732 444564 226760
rect 405516 226720 405522 226732
rect 444558 226720 444564 226732
rect 444616 226720 444622 226772
rect 248966 226692 248972 226704
rect 192996 226664 207014 226692
rect 233988 226664 248972 226692
rect 192996 226652 193002 226664
rect 206986 226556 207014 226664
rect 248966 226652 248972 226664
rect 249024 226652 249030 226704
rect 298094 226652 298100 226704
rect 298152 226692 298158 226704
rect 303614 226692 303620 226704
rect 298152 226664 303620 226692
rect 298152 226652 298158 226664
rect 303614 226652 303620 226664
rect 303672 226652 303678 226704
rect 369578 226652 369584 226704
rect 369636 226692 369642 226704
rect 402974 226692 402980 226704
rect 369636 226664 402980 226692
rect 369636 226652 369642 226664
rect 402974 226652 402980 226664
rect 403032 226652 403038 226704
rect 409690 226652 409696 226704
rect 409748 226692 409754 226704
rect 451182 226692 451188 226704
rect 409748 226664 451188 226692
rect 409748 226652 409754 226664
rect 451182 226652 451188 226664
rect 451240 226652 451246 226704
rect 237282 226584 237288 226636
rect 237340 226624 237346 226636
rect 256786 226624 256792 226636
rect 237340 226596 256792 226624
rect 237340 226584 237346 226596
rect 256786 226584 256792 226596
rect 256844 226584 256850 226636
rect 296714 226584 296720 226636
rect 296772 226624 296778 226636
rect 300210 226624 300216 226636
rect 296772 226596 300216 226624
rect 296772 226584 296778 226596
rect 300210 226584 300216 226596
rect 300268 226584 300274 226636
rect 300302 226584 300308 226636
rect 300360 226624 300366 226636
rect 306374 226624 306380 226636
rect 300360 226596 306380 226624
rect 300360 226584 300366 226596
rect 306374 226584 306380 226596
rect 306432 226584 306438 226636
rect 395798 226584 395804 226636
rect 395856 226624 395862 226636
rect 434622 226624 434628 226636
rect 395856 226596 434628 226624
rect 395856 226584 395862 226596
rect 434622 226584 434628 226596
rect 434680 226584 434686 226636
rect 251082 226556 251088 226568
rect 206986 226528 251088 226556
rect 251082 226516 251088 226528
rect 251140 226516 251146 226568
rect 254026 226516 254032 226568
rect 254084 226556 254090 226568
rect 270310 226556 270316 226568
rect 254084 226528 270316 226556
rect 254084 226516 254090 226528
rect 270310 226516 270316 226528
rect 270368 226516 270374 226568
rect 301314 226516 301320 226568
rect 301372 226556 301378 226568
rect 307754 226556 307760 226568
rect 301372 226528 307760 226556
rect 301372 226516 301378 226528
rect 307754 226516 307760 226528
rect 307812 226516 307818 226568
rect 334526 226516 334532 226568
rect 334584 226556 334590 226568
rect 351914 226556 351920 226568
rect 334584 226528 351920 226556
rect 334584 226516 334590 226528
rect 351914 226516 351920 226528
rect 351972 226516 351978 226568
rect 378686 226516 378692 226568
rect 378744 226556 378750 226568
rect 397454 226556 397460 226568
rect 378744 226528 397460 226556
rect 378744 226516 378750 226528
rect 397454 226516 397460 226528
rect 397512 226516 397518 226568
rect 401134 226516 401140 226568
rect 401192 226556 401198 226568
rect 417694 226556 417700 226568
rect 401192 226528 417700 226556
rect 401192 226516 401198 226528
rect 417694 226516 417700 226528
rect 417752 226516 417758 226568
rect 246298 226448 246304 226500
rect 246356 226488 246362 226500
rect 258534 226488 258540 226500
rect 246356 226460 258540 226488
rect 246356 226448 246362 226460
rect 258534 226448 258540 226460
rect 258592 226448 258598 226500
rect 389358 226448 389364 226500
rect 389416 226488 389422 226500
rect 408402 226488 408408 226500
rect 389416 226460 408408 226488
rect 389416 226448 389422 226460
rect 408402 226448 408408 226460
rect 408460 226448 408466 226500
rect 394786 226380 394792 226432
rect 394844 226420 394850 226432
rect 411162 226420 411168 226432
rect 394844 226392 411168 226420
rect 394844 226380 394850 226392
rect 411162 226380 411168 226392
rect 411220 226380 411226 226432
rect 197906 226312 197912 226364
rect 197964 226352 197970 226364
rect 207934 226352 207940 226364
rect 197964 226324 207940 226352
rect 197964 226312 197970 226324
rect 207934 226312 207940 226324
rect 207992 226312 207998 226364
rect 253934 226312 253940 226364
rect 253992 226352 253998 226364
rect 268930 226352 268936 226364
rect 253992 226324 268936 226352
rect 253992 226312 253998 226324
rect 268930 226312 268936 226324
rect 268988 226312 268994 226364
rect 299934 226312 299940 226364
rect 299992 226352 299998 226364
rect 304350 226352 304356 226364
rect 299992 226324 304356 226352
rect 299992 226312 299998 226324
rect 304350 226312 304356 226324
rect 304408 226312 304414 226364
rect 309870 226312 309876 226364
rect 309928 226352 309934 226364
rect 327902 226352 327908 226364
rect 309928 226324 327908 226352
rect 309928 226312 309934 226324
rect 327902 226312 327908 226324
rect 327960 226312 327966 226364
rect 151078 226244 151084 226296
rect 151136 226284 151142 226296
rect 233602 226284 233608 226296
rect 151136 226256 233608 226284
rect 151136 226244 151142 226256
rect 233602 226244 233608 226256
rect 233660 226244 233666 226296
rect 353754 226244 353760 226296
rect 353812 226284 353818 226296
rect 434806 226284 434812 226296
rect 353812 226256 434812 226284
rect 353812 226244 353818 226256
rect 434806 226244 434812 226256
rect 434864 226244 434870 226296
rect 154482 226176 154488 226228
rect 154540 226216 154546 226228
rect 235074 226216 235080 226228
rect 154540 226188 235080 226216
rect 154540 226176 154546 226188
rect 235074 226176 235080 226188
rect 235132 226176 235138 226228
rect 352282 226176 352288 226228
rect 352340 226216 352346 226228
rect 431402 226216 431408 226228
rect 352340 226188 431408 226216
rect 352340 226176 352346 226188
rect 431402 226176 431408 226188
rect 431460 226176 431466 226228
rect 433242 226176 433248 226228
rect 433300 226216 433306 226228
rect 483014 226216 483020 226228
rect 433300 226188 483020 226216
rect 433300 226176 433306 226188
rect 483014 226176 483020 226188
rect 483072 226176 483078 226228
rect 144362 226108 144368 226160
rect 144420 226148 144426 226160
rect 230750 226148 230756 226160
rect 144420 226120 230756 226148
rect 144420 226108 144426 226120
rect 230750 226108 230756 226120
rect 230808 226108 230814 226160
rect 355134 226108 355140 226160
rect 355192 226148 355198 226160
rect 438118 226148 438124 226160
rect 355192 226120 438124 226148
rect 355192 226108 355198 226120
rect 438118 226108 438124 226120
rect 438176 226108 438182 226160
rect 147766 226040 147772 226092
rect 147824 226080 147830 226092
rect 232222 226080 232228 226092
rect 147824 226052 232228 226080
rect 147824 226040 147830 226052
rect 232222 226040 232228 226052
rect 232280 226040 232286 226092
rect 359458 226040 359464 226092
rect 359516 226080 359522 226092
rect 448238 226080 448244 226092
rect 359516 226052 448244 226080
rect 359516 226040 359522 226052
rect 448238 226040 448244 226052
rect 448296 226040 448302 226092
rect 465902 226040 465908 226092
rect 465960 226080 465966 226092
rect 487798 226080 487804 226092
rect 465960 226052 487804 226080
rect 465960 226040 465966 226052
rect 487798 226040 487804 226052
rect 487856 226040 487862 226092
rect 141050 225972 141056 226024
rect 141108 226012 141114 226024
rect 229094 226012 229100 226024
rect 141108 225984 229100 226012
rect 141108 225972 141114 225984
rect 229094 225972 229100 225984
rect 229152 225972 229158 226024
rect 362310 225972 362316 226024
rect 362368 226012 362374 226024
rect 362368 225984 453620 226012
rect 362368 225972 362374 225984
rect 137646 225904 137652 225956
rect 137704 225944 137710 225956
rect 227898 225944 227904 225956
rect 137704 225916 227904 225944
rect 137704 225904 137710 225916
rect 227898 225904 227904 225916
rect 227956 225904 227962 225956
rect 362678 225904 362684 225956
rect 362736 225944 362742 225956
rect 452654 225944 452660 225956
rect 362736 225916 452660 225944
rect 362736 225904 362742 225916
rect 452654 225904 452660 225916
rect 452712 225904 452718 225956
rect 453592 225944 453620 225984
rect 453666 225972 453672 226024
rect 453724 226012 453730 226024
rect 500678 226012 500684 226024
rect 453724 225984 500684 226012
rect 453724 225972 453730 225984
rect 500678 225972 500684 225984
rect 500736 225972 500742 226024
rect 454954 225944 454960 225956
rect 453592 225916 454960 225944
rect 454954 225904 454960 225916
rect 455012 225904 455018 225956
rect 455414 225904 455420 225956
rect 455472 225944 455478 225956
rect 505738 225944 505744 225956
rect 455472 225916 505744 225944
rect 455472 225904 455478 225916
rect 505738 225904 505744 225916
rect 505796 225904 505802 225956
rect 516410 225944 516416 225956
rect 516106 225916 516416 225944
rect 134242 225836 134248 225888
rect 134300 225876 134306 225888
rect 226518 225876 226524 225888
rect 134300 225848 226524 225876
rect 134300 225836 134306 225848
rect 226518 225836 226524 225848
rect 226576 225836 226582 225888
rect 366910 225836 366916 225888
rect 366968 225876 366974 225888
rect 462498 225876 462504 225888
rect 366968 225848 462504 225876
rect 366968 225836 366974 225848
rect 462498 225836 462504 225848
rect 462556 225836 462562 225888
rect 469858 225836 469864 225888
rect 469916 225876 469922 225888
rect 516106 225876 516134 225916
rect 516410 225904 516416 225916
rect 516468 225904 516474 225956
rect 518894 225904 518900 225956
rect 518952 225944 518958 225956
rect 560386 225944 560392 225956
rect 518952 225916 560392 225944
rect 518952 225904 518958 225916
rect 560386 225904 560392 225916
rect 560444 225904 560450 225956
rect 469916 225848 516134 225876
rect 469916 225836 469922 225848
rect 516226 225836 516232 225888
rect 516284 225876 516290 225888
rect 564342 225876 564348 225888
rect 516284 225848 564348 225876
rect 516284 225836 516290 225848
rect 564342 225836 564348 225848
rect 564400 225836 564406 225888
rect 130930 225768 130936 225820
rect 130988 225808 130994 225820
rect 225046 225808 225052 225820
rect 130988 225780 225052 225808
rect 130988 225768 130994 225780
rect 225046 225768 225052 225780
rect 225104 225768 225110 225820
rect 365162 225768 365168 225820
rect 365220 225808 365226 225820
rect 461670 225808 461676 225820
rect 365220 225780 461676 225808
rect 365220 225768 365226 225780
rect 461670 225768 461676 225780
rect 461728 225768 461734 225820
rect 474734 225768 474740 225820
rect 474792 225808 474798 225820
rect 526438 225808 526444 225820
rect 474792 225780 526444 225808
rect 474792 225768 474798 225780
rect 526438 225768 526444 225780
rect 526496 225768 526502 225820
rect 127526 225700 127532 225752
rect 127584 225740 127590 225752
rect 223666 225740 223672 225752
rect 127584 225712 223672 225740
rect 127584 225700 127590 225712
rect 223666 225700 223672 225712
rect 223724 225700 223730 225752
rect 230106 225700 230112 225752
rect 230164 225740 230170 225752
rect 249610 225740 249616 225752
rect 230164 225712 249616 225740
rect 230164 225700 230170 225712
rect 249610 225700 249616 225712
rect 249668 225700 249674 225752
rect 363690 225700 363696 225752
rect 363748 225740 363754 225752
rect 458450 225740 458456 225752
rect 363748 225712 458456 225740
rect 363748 225700 363754 225712
rect 458450 225700 458456 225712
rect 458508 225700 458514 225752
rect 460934 225700 460940 225752
rect 460992 225740 460998 225752
rect 510706 225740 510712 225752
rect 460992 225712 510712 225740
rect 460992 225700 460998 225712
rect 510706 225700 510712 225712
rect 510764 225700 510770 225752
rect 516134 225700 516140 225752
rect 516192 225740 516198 225752
rect 566826 225740 566832 225752
rect 516192 225712 566832 225740
rect 516192 225700 516198 225712
rect 566826 225700 566832 225712
rect 566884 225700 566890 225752
rect 119154 225632 119160 225684
rect 119212 225672 119218 225684
rect 219710 225672 219716 225684
rect 119212 225644 219716 225672
rect 119212 225632 119218 225644
rect 219710 225632 219716 225644
rect 219768 225632 219774 225684
rect 230290 225632 230296 225684
rect 230348 225672 230354 225684
rect 249978 225672 249984 225684
rect 230348 225644 249984 225672
rect 230348 225632 230354 225644
rect 249978 225632 249984 225644
rect 250036 225632 250042 225684
rect 344462 225632 344468 225684
rect 344520 225672 344526 225684
rect 369578 225672 369584 225684
rect 344520 225644 369584 225672
rect 344520 225632 344526 225644
rect 369578 225632 369584 225644
rect 369636 225632 369642 225684
rect 369762 225632 369768 225684
rect 369820 225672 369826 225684
rect 468386 225672 468392 225684
rect 369820 225644 468392 225672
rect 369820 225632 369826 225644
rect 468386 225632 468392 225644
rect 468444 225632 468450 225684
rect 473262 225632 473268 225684
rect 473320 225672 473326 225684
rect 521654 225672 521660 225684
rect 473320 225644 521660 225672
rect 473320 225632 473326 225644
rect 521654 225632 521660 225644
rect 521712 225632 521718 225684
rect 124122 225564 124128 225616
rect 124180 225604 124186 225616
rect 222194 225604 222200 225616
rect 124180 225576 222200 225604
rect 124180 225564 124186 225576
rect 222194 225564 222200 225576
rect 222252 225564 222258 225616
rect 234522 225564 234528 225616
rect 234580 225604 234586 225616
rect 253842 225604 253848 225616
rect 234580 225576 253848 225604
rect 234580 225564 234586 225576
rect 253842 225564 253848 225576
rect 253900 225564 253906 225616
rect 366542 225564 366548 225616
rect 366600 225604 366606 225616
rect 465074 225604 465080 225616
rect 366600 225576 465080 225604
rect 366600 225564 366606 225576
rect 465074 225564 465080 225576
rect 465132 225564 465138 225616
rect 477494 225564 477500 225616
rect 477552 225604 477558 225616
rect 531498 225604 531504 225616
rect 477552 225576 531504 225604
rect 477552 225564 477558 225576
rect 531498 225564 531504 225576
rect 531556 225564 531562 225616
rect 114094 225496 114100 225548
rect 114152 225536 114158 225548
rect 217962 225536 217968 225548
rect 114152 225508 217968 225536
rect 114152 225496 114158 225508
rect 217962 225496 217968 225508
rect 218020 225496 218026 225548
rect 218054 225496 218060 225548
rect 218112 225536 218118 225548
rect 245378 225536 245384 225548
rect 218112 225508 245384 225536
rect 218112 225496 218118 225508
rect 245378 225496 245384 225508
rect 245436 225496 245442 225548
rect 355502 225496 355508 225548
rect 355560 225536 355566 225548
rect 433518 225536 433524 225548
rect 355560 225508 433524 225536
rect 355560 225496 355566 225508
rect 433518 225496 433524 225508
rect 433576 225496 433582 225548
rect 434622 225496 434628 225548
rect 434680 225536 434686 225548
rect 532786 225536 532792 225548
rect 434680 225508 532792 225536
rect 434680 225496 434686 225508
rect 532786 225496 532792 225508
rect 532844 225496 532850 225548
rect 117498 225428 117504 225480
rect 117556 225468 117562 225480
rect 219342 225468 219348 225480
rect 117556 225440 219348 225468
rect 117556 225428 117562 225440
rect 219342 225428 219348 225440
rect 219400 225428 219406 225480
rect 228450 225428 228456 225480
rect 228508 225468 228514 225480
rect 266446 225468 266452 225480
rect 228508 225440 266452 225468
rect 228508 225428 228514 225440
rect 266446 225428 266452 225440
rect 266504 225428 266510 225480
rect 339862 225428 339868 225480
rect 339920 225468 339926 225480
rect 371234 225468 371240 225480
rect 339920 225440 371240 225468
rect 339920 225428 339926 225440
rect 371234 225428 371240 225440
rect 371292 225428 371298 225480
rect 372614 225428 372620 225480
rect 372672 225468 372678 225480
rect 476022 225468 476028 225480
rect 372672 225440 476028 225468
rect 372672 225428 372678 225440
rect 476022 225428 476028 225440
rect 476080 225428 476086 225480
rect 480254 225428 480260 225480
rect 480312 225468 480318 225480
rect 536558 225468 536564 225480
rect 480312 225440 536564 225468
rect 480312 225428 480318 225440
rect 536558 225428 536564 225440
rect 536616 225428 536622 225480
rect 107378 225360 107384 225412
rect 107436 225400 107442 225412
rect 215110 225400 215116 225412
rect 107436 225372 215116 225400
rect 107436 225360 107442 225372
rect 215110 225360 215116 225372
rect 215168 225360 215174 225412
rect 218422 225360 218428 225412
rect 218480 225400 218486 225412
rect 262122 225400 262128 225412
rect 218480 225372 262128 225400
rect 218480 225360 218486 225372
rect 262122 225360 262128 225372
rect 262180 225360 262186 225412
rect 356974 225360 356980 225412
rect 357032 225400 357038 225412
rect 357032 225372 429148 225400
rect 357032 225360 357038 225372
rect 105722 225292 105728 225344
rect 105780 225332 105786 225344
rect 214006 225332 214012 225344
rect 105780 225304 214012 225332
rect 105780 225292 105786 225304
rect 214006 225292 214012 225304
rect 214064 225292 214070 225344
rect 221734 225292 221740 225344
rect 221792 225332 221798 225344
rect 263594 225332 263600 225344
rect 221792 225304 263600 225332
rect 221792 225292 221798 225304
rect 263594 225292 263600 225304
rect 263652 225292 263658 225344
rect 358354 225292 358360 225344
rect 358412 225332 358418 225344
rect 429010 225332 429016 225344
rect 358412 225304 429016 225332
rect 358412 225292 358418 225304
rect 429010 225292 429016 225304
rect 429068 225292 429074 225344
rect 429120 225332 429148 225372
rect 438854 225360 438860 225412
rect 438912 225400 438918 225412
rect 541434 225400 541440 225412
rect 438912 225372 541440 225400
rect 438912 225360 438918 225372
rect 541434 225360 541440 225372
rect 541492 225360 541498 225412
rect 439038 225332 439044 225344
rect 429120 225304 439044 225332
rect 439038 225292 439044 225304
rect 439096 225292 439102 225344
rect 441614 225292 441620 225344
rect 441672 225332 441678 225344
rect 545758 225332 545764 225344
rect 441672 225304 545764 225332
rect 441672 225292 441678 225304
rect 545758 225292 545764 225304
rect 545816 225292 545822 225344
rect 90542 225224 90548 225276
rect 90600 225264 90606 225276
rect 197906 225264 197912 225276
rect 90600 225236 197912 225264
rect 90600 225224 90606 225236
rect 197906 225224 197912 225236
rect 197964 225224 197970 225276
rect 198182 225224 198188 225276
rect 198240 225264 198246 225276
rect 253566 225264 253572 225276
rect 198240 225236 253572 225264
rect 198240 225224 198246 225236
rect 253566 225224 253572 225236
rect 253624 225224 253630 225276
rect 357986 225224 357992 225276
rect 358044 225264 358050 225276
rect 358044 225236 444328 225264
rect 358044 225224 358050 225236
rect 100662 225156 100668 225208
rect 100720 225196 100726 225208
rect 212258 225196 212264 225208
rect 100720 225168 212264 225196
rect 100720 225156 100726 225168
rect 212258 225156 212264 225168
rect 212316 225156 212322 225208
rect 225138 225156 225144 225208
rect 225196 225196 225202 225208
rect 264974 225196 264980 225208
rect 225196 225168 264980 225196
rect 225196 225156 225202 225168
rect 264974 225156 264980 225168
rect 265032 225156 265038 225208
rect 317782 225156 317788 225208
rect 317840 225196 317846 225208
rect 348970 225196 348976 225208
rect 317840 225168 348976 225196
rect 317840 225156 317846 225168
rect 348970 225156 348976 225168
rect 349028 225156 349034 225208
rect 361206 225156 361212 225208
rect 361264 225196 361270 225208
rect 444300 225196 444328 225236
rect 444558 225224 444564 225276
rect 444616 225264 444622 225276
rect 557442 225264 557448 225276
rect 444616 225236 557448 225264
rect 444616 225224 444622 225236
rect 557442 225224 557448 225236
rect 557500 225224 557506 225276
rect 444834 225196 444840 225208
rect 361264 225168 444236 225196
rect 444300 225168 444840 225196
rect 361264 225156 361270 225168
rect 103974 225088 103980 225140
rect 104032 225128 104038 225140
rect 213638 225128 213644 225140
rect 104032 225100 213644 225128
rect 104032 225088 104038 225100
rect 213638 225088 213644 225100
rect 213696 225088 213702 225140
rect 215018 225088 215024 225140
rect 215076 225128 215082 225140
rect 260742 225128 260748 225140
rect 215076 225100 260748 225128
rect 215076 225088 215082 225100
rect 260742 225088 260748 225100
rect 260800 225088 260806 225140
rect 319162 225088 319168 225140
rect 319220 225128 319226 225140
rect 352374 225128 352380 225140
rect 319220 225100 352380 225128
rect 319220 225088 319226 225100
rect 352374 225088 352380 225100
rect 352432 225088 352438 225140
rect 360838 225088 360844 225140
rect 360896 225128 360902 225140
rect 444098 225128 444104 225140
rect 360896 225100 444104 225128
rect 360896 225088 360902 225100
rect 444098 225088 444104 225100
rect 444156 225088 444162 225140
rect 444208 225128 444236 225168
rect 444834 225156 444840 225168
rect 444892 225156 444898 225208
rect 449618 225156 449624 225208
rect 449676 225196 449682 225208
rect 561214 225196 561220 225208
rect 449676 225168 561220 225196
rect 449676 225156 449682 225168
rect 561214 225156 561220 225168
rect 561272 225156 561278 225208
rect 449066 225128 449072 225140
rect 444208 225100 449072 225128
rect 449066 225088 449072 225100
rect 449124 225088 449130 225140
rect 451182 225088 451188 225140
rect 451240 225128 451246 225140
rect 565998 225128 566004 225140
rect 451240 225100 566004 225128
rect 451240 225088 451246 225100
rect 565998 225088 566004 225100
rect 566056 225088 566062 225140
rect 95602 225020 95608 225072
rect 95660 225060 95666 225072
rect 209498 225060 209504 225072
rect 95660 225032 209504 225060
rect 95660 225020 95666 225032
rect 209498 225020 209504 225032
rect 209556 225020 209562 225072
rect 211706 225020 211712 225072
rect 211764 225060 211770 225072
rect 259270 225060 259276 225072
rect 211764 225032 259276 225060
rect 211764 225020 211770 225032
rect 259270 225020 259276 225032
rect 259328 225020 259334 225072
rect 313458 225020 313464 225072
rect 313516 225060 313522 225072
rect 338850 225060 338856 225072
rect 313516 225032 338856 225060
rect 313516 225020 313522 225032
rect 338850 225020 338856 225032
rect 338908 225020 338914 225072
rect 344094 225020 344100 225072
rect 344152 225060 344158 225072
rect 408678 225060 408684 225072
rect 344152 225032 408684 225060
rect 344152 225020 344158 225032
rect 408678 225020 408684 225032
rect 408736 225020 408742 225072
rect 408954 225020 408960 225072
rect 409012 225060 409018 225072
rect 563698 225060 563704 225072
rect 409012 225032 563704 225060
rect 409012 225020 409018 225032
rect 563698 225020 563704 225032
rect 563756 225020 563762 225072
rect 88886 224952 88892 225004
rect 88944 224992 88950 225004
rect 206830 224992 206836 225004
rect 88944 224964 206836 224992
rect 88944 224952 88950 224964
rect 206830 224952 206836 224964
rect 206888 224952 206894 225004
rect 208302 224952 208308 225004
rect 208360 224992 208366 225004
rect 257890 224992 257896 225004
rect 208360 224964 257896 224992
rect 208360 224952 208366 224964
rect 257890 224952 257896 224964
rect 257948 224952 257954 225004
rect 316310 224952 316316 225004
rect 316368 224992 316374 225004
rect 345658 224992 345664 225004
rect 316368 224964 345664 224992
rect 316368 224952 316374 224964
rect 345658 224952 345664 224964
rect 345716 224952 345722 225004
rect 345842 224952 345848 225004
rect 345900 224992 345906 225004
rect 410794 224992 410800 225004
rect 345900 224964 410800 224992
rect 345900 224952 345906 224964
rect 410794 224952 410800 224964
rect 410852 224952 410858 225004
rect 411162 224992 411168 225004
rect 410996 224964 411168 224992
rect 73706 224884 73712 224936
rect 73764 224924 73770 224936
rect 200850 224924 200856 224936
rect 73764 224896 200856 224924
rect 73764 224884 73770 224896
rect 200850 224884 200856 224896
rect 200908 224884 200914 224936
rect 201402 224884 201408 224936
rect 201460 224924 201466 224936
rect 255038 224924 255044 224936
rect 201460 224896 255044 224924
rect 201460 224884 201466 224896
rect 255038 224884 255044 224896
rect 255096 224884 255102 224936
rect 314930 224884 314936 224936
rect 314988 224924 314994 224936
rect 342438 224924 342444 224936
rect 314988 224896 342444 224924
rect 314988 224884 314994 224896
rect 342438 224884 342444 224896
rect 342496 224884 342502 224936
rect 343726 224884 343732 224936
rect 343784 224924 343790 224936
rect 410996 224924 411024 224964
rect 411162 224952 411168 224964
rect 411220 224952 411226 225004
rect 411530 224952 411536 225004
rect 411588 224992 411594 225004
rect 570230 224992 570236 225004
rect 411588 224964 570236 224992
rect 411588 224952 411594 224964
rect 570230 224952 570236 224964
rect 570288 224952 570294 225004
rect 343784 224896 411024 224924
rect 343784 224884 343790 224896
rect 411070 224884 411076 224936
rect 411128 224924 411134 224936
rect 568574 224924 568580 224936
rect 411128 224896 568580 224924
rect 411128 224884 411134 224896
rect 568574 224884 568580 224896
rect 568632 224884 568638 224936
rect 161198 224816 161204 224868
rect 161256 224856 161262 224868
rect 237926 224856 237932 224868
rect 161256 224828 237932 224856
rect 161256 224816 161262 224828
rect 237926 224816 237932 224828
rect 237984 224816 237990 224868
rect 354122 224816 354128 224868
rect 354180 224856 354186 224868
rect 432230 224856 432236 224868
rect 354180 224828 432236 224856
rect 354180 224816 354186 224828
rect 432230 224816 432236 224828
rect 432288 224816 432294 224868
rect 433150 224816 433156 224868
rect 433208 224856 433214 224868
rect 477770 224856 477776 224868
rect 433208 224828 477776 224856
rect 433208 224816 433214 224828
rect 477770 224816 477776 224828
rect 477828 224816 477834 224868
rect 157794 224748 157800 224800
rect 157852 224788 157858 224800
rect 236454 224788 236460 224800
rect 157852 224760 236460 224788
rect 157852 224748 157858 224760
rect 236454 224748 236460 224760
rect 236512 224748 236518 224800
rect 349430 224748 349436 224800
rect 349488 224788 349494 224800
rect 425054 224788 425060 224800
rect 349488 224760 425060 224788
rect 349488 224748 349494 224760
rect 425054 224748 425060 224760
rect 425112 224748 425118 224800
rect 428366 224748 428372 224800
rect 428424 224788 428430 224800
rect 470962 224788 470968 224800
rect 428424 224760 470968 224788
rect 428424 224748 428430 224760
rect 470962 224748 470968 224760
rect 471020 224748 471026 224800
rect 167914 224680 167920 224732
rect 167972 224720 167978 224732
rect 240778 224720 240784 224732
rect 167972 224692 240784 224720
rect 167972 224680 167978 224692
rect 240778 224680 240784 224692
rect 240836 224680 240842 224732
rect 352650 224680 352656 224732
rect 352708 224720 352714 224732
rect 428918 224720 428924 224732
rect 352708 224692 428924 224720
rect 352708 224680 352714 224692
rect 428918 224680 428924 224692
rect 428976 224680 428982 224732
rect 429010 224680 429016 224732
rect 429068 224720 429074 224732
rect 442350 224720 442356 224732
rect 429068 224692 442356 224720
rect 429068 224680 429074 224692
rect 442350 224680 442356 224692
rect 442408 224680 442414 224732
rect 444098 224680 444104 224732
rect 444156 224720 444162 224732
rect 451550 224720 451556 224732
rect 444156 224692 451556 224720
rect 444156 224680 444162 224692
rect 451550 224680 451556 224692
rect 451608 224680 451614 224732
rect 164602 224612 164608 224664
rect 164660 224652 164666 224664
rect 239306 224652 239312 224664
rect 164660 224624 239312 224652
rect 164660 224612 164666 224624
rect 239306 224612 239312 224624
rect 239364 224612 239370 224664
rect 350902 224612 350908 224664
rect 350960 224652 350966 224664
rect 427998 224652 428004 224664
rect 350960 224624 428004 224652
rect 350960 224612 350966 224624
rect 427998 224612 428004 224624
rect 428056 224612 428062 224664
rect 170950 224544 170956 224596
rect 171008 224584 171014 224596
rect 242158 224584 242164 224596
rect 171008 224556 242164 224584
rect 171008 224544 171014 224556
rect 242158 224544 242164 224556
rect 242216 224544 242222 224596
rect 349798 224544 349804 224596
rect 349856 224584 349862 224596
rect 409690 224584 409696 224596
rect 349856 224556 409696 224584
rect 349856 224544 349862 224556
rect 409690 224544 409696 224556
rect 409748 224544 409754 224596
rect 421282 224584 421288 224596
rect 409984 224556 421288 224584
rect 174630 224476 174636 224528
rect 174688 224516 174694 224528
rect 243354 224516 243360 224528
rect 174688 224488 243360 224516
rect 174688 224476 174694 224488
rect 243354 224476 243360 224488
rect 243412 224476 243418 224528
rect 346578 224476 346584 224528
rect 346636 224516 346642 224528
rect 409598 224516 409604 224528
rect 346636 224488 409604 224516
rect 346636 224476 346642 224488
rect 409598 224476 409604 224488
rect 409656 224476 409662 224528
rect 181346 224408 181352 224460
rect 181404 224448 181410 224460
rect 246482 224448 246488 224460
rect 181404 224420 246488 224448
rect 181404 224408 181410 224420
rect 246482 224408 246488 224420
rect 246540 224408 246546 224460
rect 348050 224408 348056 224460
rect 348108 224448 348114 224460
rect 409984 224448 410012 224556
rect 421282 224544 421288 224556
rect 421340 224544 421346 224596
rect 422294 224544 422300 224596
rect 422352 224584 422358 224596
rect 464246 224584 464252 224596
rect 422352 224556 464252 224584
rect 422352 224544 422358 224556
rect 464246 224544 464252 224556
rect 464304 224544 464310 224596
rect 416774 224476 416780 224528
rect 416832 224516 416838 224528
rect 457438 224516 457444 224528
rect 416832 224488 457444 224516
rect 416832 224476 416838 224488
rect 457438 224476 457444 224488
rect 457496 224476 457502 224528
rect 348108 224420 410012 224448
rect 348108 224408 348114 224420
rect 410794 224408 410800 224460
rect 410852 224448 410858 224460
rect 412082 224448 412088 224460
rect 410852 224420 412088 224448
rect 410852 224408 410858 224420
rect 412082 224408 412088 224420
rect 412140 224408 412146 224460
rect 178034 224340 178040 224392
rect 178092 224380 178098 224392
rect 245010 224380 245016 224392
rect 178092 224352 245016 224380
rect 178092 224340 178098 224352
rect 245010 224340 245016 224352
rect 245068 224340 245074 224392
rect 340230 224340 340236 224392
rect 340288 224380 340294 224392
rect 371142 224380 371148 224392
rect 340288 224352 371148 224380
rect 340288 224340 340294 224352
rect 371142 224340 371148 224352
rect 371200 224340 371206 224392
rect 372890 224340 372896 224392
rect 372948 224380 372954 224392
rect 441614 224380 441620 224392
rect 372948 224352 441620 224380
rect 372948 224340 372954 224352
rect 441614 224340 441620 224352
rect 441672 224340 441678 224392
rect 184750 224272 184756 224324
rect 184808 224312 184814 224324
rect 247862 224312 247868 224324
rect 184808 224284 247868 224312
rect 184808 224272 184814 224284
rect 247862 224272 247868 224284
rect 247920 224272 247926 224324
rect 348418 224272 348424 224324
rect 348476 224312 348482 224324
rect 418798 224312 418804 224324
rect 348476 224284 418804 224312
rect 348476 224272 348482 224284
rect 418798 224272 418804 224284
rect 418856 224272 418862 224324
rect 188154 224204 188160 224256
rect 188212 224244 188218 224256
rect 249334 224244 249340 224256
rect 188212 224216 249340 224244
rect 188212 224204 188218 224216
rect 249334 224204 249340 224216
rect 249392 224204 249398 224256
rect 346946 224204 346952 224256
rect 347004 224244 347010 224256
rect 415394 224244 415400 224256
rect 347004 224216 415400 224244
rect 347004 224204 347010 224216
rect 415394 224204 415400 224216
rect 415452 224204 415458 224256
rect 415486 224204 415492 224256
rect 415544 224244 415550 224256
rect 450722 224244 450728 224256
rect 415544 224216 450728 224244
rect 415544 224204 415550 224216
rect 450722 224204 450728 224216
rect 450780 224204 450786 224256
rect 191466 224136 191472 224188
rect 191524 224176 191530 224188
rect 250714 224176 250720 224188
rect 191524 224148 250720 224176
rect 191524 224136 191530 224148
rect 250714 224136 250720 224148
rect 250772 224136 250778 224188
rect 339494 224136 339500 224188
rect 339552 224176 339558 224188
rect 394786 224176 394792 224188
rect 339552 224148 394792 224176
rect 339552 224136 339558 224148
rect 394786 224136 394792 224148
rect 394844 224136 394850 224188
rect 402974 224136 402980 224188
rect 403032 224176 403038 224188
rect 469214 224176 469220 224188
rect 403032 224148 469220 224176
rect 403032 224136 403038 224148
rect 469214 224136 469220 224148
rect 469272 224136 469278 224188
rect 139302 224068 139308 224120
rect 139360 224108 139366 224120
rect 194870 224108 194876 224120
rect 139360 224080 194876 224108
rect 139360 224068 139366 224080
rect 194870 224068 194876 224080
rect 194928 224068 194934 224120
rect 194962 224068 194968 224120
rect 195020 224108 195026 224120
rect 252186 224108 252192 224120
rect 195020 224080 252192 224108
rect 195020 224068 195026 224080
rect 252186 224068 252192 224080
rect 252244 224068 252250 224120
rect 335170 224068 335176 224120
rect 335228 224108 335234 224120
rect 391014 224108 391020 224120
rect 335228 224080 391020 224108
rect 335228 224068 335234 224080
rect 391014 224068 391020 224080
rect 391072 224068 391078 224120
rect 400214 224068 400220 224120
rect 400272 224108 400278 224120
rect 445662 224108 445668 224120
rect 400272 224080 445668 224108
rect 400272 224068 400278 224080
rect 445662 224068 445668 224080
rect 445720 224068 445726 224120
rect 155862 224000 155868 224052
rect 155920 224040 155926 224052
rect 155920 224012 189672 224040
rect 155920 224000 155926 224012
rect 189644 223768 189672 224012
rect 209590 224000 209596 224052
rect 209648 224040 209654 224052
rect 236822 224040 236828 224052
rect 209648 224012 236828 224040
rect 209648 224000 209654 224012
rect 236822 224000 236828 224012
rect 236880 224000 236886 224052
rect 343082 224000 343088 224052
rect 343140 224040 343146 224052
rect 368106 224040 368112 224052
rect 343140 224012 368112 224040
rect 343140 224000 343146 224012
rect 368106 224000 368112 224012
rect 368164 224000 368170 224052
rect 376662 224000 376668 224052
rect 376720 224040 376726 224052
rect 376720 224012 409644 224040
rect 376720 224000 376726 224012
rect 204898 223932 204904 223984
rect 204956 223972 204962 223984
rect 256418 223972 256424 223984
rect 204956 223944 256424 223972
rect 204956 223932 204962 223944
rect 256418 223932 256424 223944
rect 256476 223932 256482 223984
rect 383746 223932 383752 223984
rect 383804 223972 383810 223984
rect 407850 223972 407856 223984
rect 383804 223944 407856 223972
rect 383804 223932 383810 223944
rect 407850 223932 407856 223944
rect 407908 223932 407914 223984
rect 409616 223972 409644 224012
rect 409690 224000 409696 224052
rect 409748 224040 409754 224052
rect 422294 224040 422300 224052
rect 409748 224012 422300 224040
rect 409748 224000 409754 224012
rect 422294 224000 422300 224012
rect 422352 224000 422358 224052
rect 414566 223972 414572 223984
rect 409616 223944 414572 223972
rect 414566 223932 414572 223944
rect 414624 223932 414630 223984
rect 204254 223864 204260 223916
rect 204312 223904 204318 223916
rect 252462 223904 252468 223916
rect 204312 223876 252468 223904
rect 204312 223864 204318 223876
rect 252462 223864 252468 223876
rect 252520 223864 252526 223916
rect 383654 223864 383660 223916
rect 383712 223904 383718 223916
rect 404446 223904 404452 223916
rect 383712 223876 404452 223904
rect 383712 223864 383718 223876
rect 404446 223864 404452 223876
rect 404504 223864 404510 223916
rect 415302 223864 415308 223916
rect 415360 223904 415366 223916
rect 444374 223904 444380 223916
rect 415360 223876 444380 223904
rect 415360 223864 415366 223876
rect 444374 223864 444380 223876
rect 444432 223864 444438 223916
rect 189718 223796 189724 223848
rect 189776 223836 189782 223848
rect 232498 223836 232504 223848
rect 189776 223808 232504 223836
rect 189776 223796 189782 223808
rect 232498 223796 232504 223808
rect 232556 223796 232562 223848
rect 395154 223796 395160 223848
rect 395212 223836 395218 223848
rect 405734 223836 405740 223848
rect 395212 223808 405740 223836
rect 395212 223796 395218 223808
rect 405734 223796 405740 223808
rect 405792 223796 405798 223848
rect 410978 223796 410984 223848
rect 411036 223836 411042 223848
rect 430574 223836 430580 223848
rect 411036 223808 430580 223836
rect 411036 223796 411042 223808
rect 430574 223796 430580 223808
rect 430632 223796 430638 223848
rect 209406 223768 209412 223780
rect 189644 223740 209412 223768
rect 209406 223728 209412 223740
rect 209464 223728 209470 223780
rect 213086 223728 213092 223780
rect 213144 223768 213150 223780
rect 242526 223768 242532 223780
rect 213144 223740 242532 223768
rect 213144 223728 213150 223740
rect 242526 223728 242532 223740
rect 242584 223728 242590 223780
rect 409598 223728 409604 223780
rect 409656 223768 409662 223780
rect 417970 223768 417976 223780
rect 409656 223740 417976 223768
rect 409656 223728 409662 223740
rect 417970 223728 417976 223740
rect 418028 223728 418034 223780
rect 171042 223660 171048 223712
rect 171100 223700 171106 223712
rect 206554 223700 206560 223712
rect 171100 223672 206560 223700
rect 171100 223660 171106 223672
rect 206554 223660 206560 223672
rect 206612 223660 206618 223712
rect 215202 223660 215208 223712
rect 215260 223700 215266 223712
rect 239674 223700 239680 223712
rect 215260 223672 239680 223700
rect 215260 223660 215266 223672
rect 239674 223660 239680 223672
rect 239732 223660 239738 223712
rect 182174 223592 182180 223644
rect 182232 223632 182238 223644
rect 192294 223632 192300 223644
rect 182232 223604 192300 223632
rect 182232 223592 182238 223604
rect 192294 223592 192300 223604
rect 192352 223592 192358 223644
rect 230014 223632 230020 223644
rect 218072 223604 230020 223632
rect 140130 223524 140136 223576
rect 140188 223564 140194 223576
rect 218072 223564 218100 223604
rect 230014 223592 230020 223604
rect 230072 223592 230078 223644
rect 348142 223632 348148 223644
rect 347700 223604 348148 223632
rect 140188 223536 218100 223564
rect 140188 223524 140194 223536
rect 278682 223524 278688 223576
rect 278740 223564 278746 223576
rect 287790 223564 287796 223576
rect 278740 223536 287796 223564
rect 278740 223524 278746 223536
rect 287790 223524 287796 223536
rect 287848 223524 287854 223576
rect 318426 223524 318432 223576
rect 318484 223564 318490 223576
rect 347700 223564 347728 223604
rect 348142 223592 348148 223604
rect 348200 223592 348206 223644
rect 408218 223592 408224 223644
rect 408276 223632 408282 223644
rect 414014 223632 414020 223644
rect 408276 223604 414020 223632
rect 408276 223592 408282 223604
rect 414014 223592 414020 223604
rect 414072 223592 414078 223644
rect 433518 223592 433524 223644
rect 433576 223632 433582 223644
rect 435634 223632 435640 223644
rect 433576 223604 435640 223632
rect 433576 223592 433582 223604
rect 435634 223592 435640 223604
rect 435692 223592 435698 223644
rect 318484 223536 347728 223564
rect 318484 223524 318490 223536
rect 347774 223524 347780 223576
rect 347832 223564 347838 223576
rect 383654 223564 383660 223576
rect 347832 223536 383660 223564
rect 347832 223524 347838 223536
rect 383654 223524 383660 223536
rect 383712 223524 383718 223576
rect 386506 223524 386512 223576
rect 386564 223564 386570 223576
rect 511350 223564 511356 223576
rect 386564 223536 511356 223564
rect 386564 223524 386570 223536
rect 511350 223524 511356 223536
rect 511408 223524 511414 223576
rect 674558 223524 674564 223576
rect 674616 223564 674622 223576
rect 675846 223564 675852 223576
rect 674616 223536 675852 223564
rect 674616 223524 674622 223536
rect 675846 223524 675852 223536
rect 675904 223524 675910 223576
rect 153654 223456 153660 223508
rect 153712 223496 153718 223508
rect 235718 223496 235724 223508
rect 153712 223468 235724 223496
rect 153712 223456 153718 223468
rect 235718 223456 235724 223468
rect 235776 223456 235782 223508
rect 322382 223456 322388 223508
rect 322440 223496 322446 223508
rect 360746 223496 360752 223508
rect 322440 223468 360752 223496
rect 322440 223456 322446 223468
rect 360746 223456 360752 223468
rect 360804 223456 360810 223508
rect 495802 223456 495808 223508
rect 495860 223496 495866 223508
rect 607582 223496 607588 223508
rect 495860 223468 607588 223496
rect 495860 223456 495866 223468
rect 607582 223456 607588 223468
rect 607640 223456 607646 223508
rect 87138 223388 87144 223440
rect 87196 223428 87202 223440
rect 171042 223428 171048 223440
rect 87196 223400 171048 223428
rect 87196 223388 87202 223400
rect 171042 223388 171048 223400
rect 171100 223388 171106 223440
rect 177206 223388 177212 223440
rect 177264 223428 177270 223440
rect 245746 223428 245752 223440
rect 177264 223400 245752 223428
rect 177264 223388 177270 223400
rect 245746 223388 245752 223400
rect 245804 223388 245810 223440
rect 333946 223400 343588 223428
rect 146938 223320 146944 223372
rect 146996 223360 147002 223372
rect 232866 223360 232872 223372
rect 146996 223332 232872 223360
rect 146996 223320 147002 223332
rect 232866 223320 232872 223332
rect 232924 223320 232930 223372
rect 326982 223320 326988 223372
rect 327040 223360 327046 223372
rect 333946 223360 333974 223400
rect 327040 223332 333974 223360
rect 343560 223360 343588 223400
rect 343634 223388 343640 223440
rect 343692 223428 343698 223440
rect 361758 223428 361764 223440
rect 343692 223400 361764 223428
rect 343692 223388 343698 223400
rect 361758 223388 361764 223400
rect 361816 223388 361822 223440
rect 387242 223388 387248 223440
rect 387300 223428 387306 223440
rect 513374 223428 513380 223440
rect 387300 223400 513380 223428
rect 387300 223388 387306 223400
rect 513374 223388 513380 223400
rect 513432 223388 513438 223440
rect 368290 223360 368296 223372
rect 343560 223332 368296 223360
rect 327040 223320 327046 223332
rect 368290 223320 368296 223332
rect 368348 223320 368354 223372
rect 389726 223320 389732 223372
rect 389784 223360 389790 223372
rect 518894 223360 518900 223372
rect 389784 223332 518900 223360
rect 389784 223320 389790 223332
rect 518894 223320 518900 223332
rect 518952 223320 518958 223372
rect 543550 223320 543556 223372
rect 543608 223360 543614 223372
rect 616414 223360 616420 223372
rect 543608 223332 616420 223360
rect 543608 223320 543614 223332
rect 616414 223320 616420 223332
rect 616472 223320 616478 223372
rect 148594 223252 148600 223304
rect 148652 223292 148658 223304
rect 233234 223292 233240 223304
rect 148652 223264 233240 223292
rect 148652 223252 148658 223264
rect 233234 223252 233240 223264
rect 233292 223252 233298 223304
rect 246666 223252 246672 223304
rect 246724 223292 246730 223304
rect 256050 223292 256056 223304
rect 246724 223264 256056 223292
rect 246724 223252 246730 223264
rect 256050 223252 256056 223264
rect 256108 223252 256114 223304
rect 269666 223252 269672 223304
rect 269724 223292 269730 223304
rect 284570 223292 284576 223304
rect 269724 223264 284576 223292
rect 269724 223252 269730 223264
rect 284570 223252 284576 223264
rect 284628 223252 284634 223304
rect 324130 223252 324136 223304
rect 324188 223292 324194 223304
rect 343450 223292 343456 223304
rect 324188 223264 343456 223292
rect 324188 223252 324194 223264
rect 343450 223252 343456 223264
rect 343508 223252 343514 223304
rect 343542 223252 343548 223304
rect 343600 223292 343606 223304
rect 364334 223292 364340 223304
rect 343600 223264 364340 223292
rect 343600 223252 343606 223264
rect 364334 223252 364340 223264
rect 364392 223252 364398 223304
rect 391934 223252 391940 223304
rect 391992 223292 391998 223304
rect 523954 223292 523960 223304
rect 391992 223264 523960 223292
rect 391992 223252 391998 223264
rect 523954 223252 523960 223264
rect 524012 223252 524018 223304
rect 552014 223252 552020 223304
rect 552072 223292 552078 223304
rect 553670 223292 553676 223304
rect 552072 223264 553676 223292
rect 552072 223252 552078 223264
rect 553670 223252 553676 223264
rect 553728 223292 553734 223304
rect 618254 223292 618260 223304
rect 553728 223264 618260 223292
rect 553728 223252 553734 223264
rect 618254 223252 618260 223264
rect 618312 223252 618318 223304
rect 60274 223184 60280 223236
rect 60332 223224 60338 223236
rect 139302 223224 139308 223236
rect 60332 223196 139308 223224
rect 60332 223184 60338 223196
rect 139302 223184 139308 223196
rect 139360 223184 139366 223236
rect 141878 223184 141884 223236
rect 141936 223224 141942 223236
rect 230382 223224 230388 223236
rect 141936 223196 230388 223224
rect 141936 223184 141942 223196
rect 230382 223184 230388 223196
rect 230440 223184 230446 223236
rect 248506 223224 248512 223236
rect 237346 223196 248512 223224
rect 135162 223116 135168 223168
rect 135220 223156 135226 223168
rect 227530 223156 227536 223168
rect 135220 223128 227536 223156
rect 135220 223116 135226 223128
rect 227530 223116 227536 223128
rect 227588 223116 227594 223168
rect 133414 223048 133420 223100
rect 133472 223088 133478 223100
rect 227162 223088 227168 223100
rect 133472 223060 227168 223088
rect 133472 223048 133478 223060
rect 227162 223048 227168 223060
rect 227220 223048 227226 223100
rect 231026 223048 231032 223100
rect 231084 223088 231090 223100
rect 237346 223088 237374 223196
rect 248506 223184 248512 223196
rect 248564 223184 248570 223236
rect 326338 223184 326344 223236
rect 326396 223224 326402 223236
rect 369118 223224 369124 223236
rect 326396 223196 369124 223224
rect 326396 223184 326402 223196
rect 369118 223184 369124 223196
rect 369176 223184 369182 223236
rect 394050 223184 394056 223236
rect 394108 223224 394114 223236
rect 529014 223224 529020 223236
rect 394108 223196 529020 223224
rect 394108 223184 394114 223196
rect 529014 223184 529020 223196
rect 529072 223184 529078 223236
rect 545758 223184 545764 223236
rect 545816 223224 545822 223236
rect 616874 223224 616880 223236
rect 545816 223196 616880 223224
rect 545816 223184 545822 223196
rect 616874 223184 616880 223196
rect 616932 223184 616938 223236
rect 242802 223116 242808 223168
rect 242860 223156 242866 223168
rect 258442 223156 258448 223168
rect 242860 223128 258448 223156
rect 242860 223116 242866 223128
rect 258442 223116 258448 223128
rect 258500 223116 258506 223168
rect 328454 223116 328460 223168
rect 328512 223156 328518 223168
rect 371694 223156 371700 223168
rect 328512 223128 371700 223156
rect 328512 223116 328518 223128
rect 371694 223116 371700 223128
rect 371752 223116 371758 223168
rect 396166 223116 396172 223168
rect 396224 223156 396230 223168
rect 533982 223156 533988 223168
rect 396224 223128 533988 223156
rect 396224 223116 396230 223128
rect 533982 223116 533988 223128
rect 534040 223116 534046 223168
rect 535546 223116 535552 223168
rect 535604 223156 535610 223168
rect 536098 223156 536104 223168
rect 535604 223128 536104 223156
rect 535604 223116 535610 223128
rect 536098 223116 536104 223128
rect 536156 223156 536162 223168
rect 615034 223156 615040 223168
rect 536156 223128 615040 223156
rect 536156 223116 536162 223128
rect 615034 223116 615040 223128
rect 615092 223116 615098 223168
rect 231084 223060 237374 223088
rect 231084 223048 231090 223060
rect 246758 223048 246764 223100
rect 246816 223088 246822 223100
rect 248414 223088 248420 223100
rect 246816 223060 248420 223088
rect 246816 223048 246822 223060
rect 248414 223048 248420 223060
rect 248472 223048 248478 223100
rect 271414 223048 271420 223100
rect 271472 223088 271478 223100
rect 285674 223088 285680 223100
rect 271472 223060 285680 223088
rect 271472 223048 271478 223060
rect 285674 223048 285680 223060
rect 285732 223048 285738 223100
rect 325602 223048 325608 223100
rect 325660 223088 325666 223100
rect 364978 223088 364984 223100
rect 325660 223060 364984 223088
rect 325660 223048 325666 223060
rect 364978 223048 364984 223060
rect 365036 223048 365042 223100
rect 398650 223048 398656 223100
rect 398708 223088 398714 223100
rect 539870 223088 539876 223100
rect 398708 223060 539876 223088
rect 398708 223048 398714 223060
rect 539870 223048 539876 223060
rect 539928 223048 539934 223100
rect 560202 223048 560208 223100
rect 560260 223088 560266 223100
rect 619174 223088 619180 223100
rect 560260 223060 619180 223088
rect 560260 223048 560266 223060
rect 619174 223048 619180 223060
rect 619232 223048 619238 223100
rect 128354 222980 128360 223032
rect 128412 223020 128418 223032
rect 224678 223020 224684 223032
rect 128412 222992 224684 223020
rect 128412 222980 128418 222992
rect 224678 222980 224684 222992
rect 224736 222980 224742 223032
rect 236086 222980 236092 223032
rect 236144 223020 236150 223032
rect 254026 223020 254032 223032
rect 236144 222992 254032 223020
rect 236144 222980 236150 222992
rect 254026 222980 254032 222992
rect 254084 222980 254090 223032
rect 263778 222980 263784 223032
rect 263836 223020 263842 223032
rect 280982 223020 280988 223032
rect 263836 222992 280988 223020
rect 263836 222980 263842 222992
rect 280982 222980 280988 222992
rect 281040 222980 281046 223032
rect 324038 222980 324044 223032
rect 324096 223020 324102 223032
rect 343542 223020 343548 223032
rect 324096 222992 343548 223020
rect 324096 222980 324102 222992
rect 343542 222980 343548 222992
rect 343600 222980 343606 223032
rect 343634 222980 343640 223032
rect 343692 223020 343698 223032
rect 367462 223020 367468 223032
rect 343692 222992 367468 223020
rect 343692 222980 343698 222992
rect 367462 222980 367468 222992
rect 367520 222980 367526 223032
rect 398282 222980 398288 223032
rect 398340 223020 398346 223032
rect 539042 223020 539048 223032
rect 398340 222992 539048 223020
rect 398340 222980 398346 222992
rect 539042 222980 539048 222992
rect 539100 222980 539106 223032
rect 541434 222980 541440 223032
rect 541492 223020 541498 223032
rect 615954 223020 615960 223032
rect 541492 222992 615960 223020
rect 541492 222980 541498 222992
rect 615954 222980 615960 222992
rect 616012 222980 616018 223032
rect 126698 222912 126704 222964
rect 126756 222952 126762 222964
rect 224034 222952 224040 222964
rect 126756 222924 224040 222952
rect 126756 222912 126762 222924
rect 224034 222912 224040 222924
rect 224092 222912 224098 222964
rect 232682 222912 232688 222964
rect 232740 222952 232746 222964
rect 253934 222952 253940 222964
rect 232740 222924 253940 222952
rect 232740 222912 232746 222924
rect 253934 222912 253940 222924
rect 253992 222912 253998 222964
rect 266354 222912 266360 222964
rect 266412 222952 266418 222964
rect 283190 222952 283196 222964
rect 266412 222924 283196 222952
rect 266412 222912 266418 222924
rect 283190 222912 283196 222924
rect 283248 222912 283254 222964
rect 326614 222912 326620 222964
rect 326672 222952 326678 222964
rect 370866 222952 370872 222964
rect 326672 222924 370872 222952
rect 326672 222912 326678 222924
rect 370866 222912 370872 222924
rect 370924 222912 370930 222964
rect 371234 222912 371240 222964
rect 371292 222952 371298 222964
rect 398558 222952 398564 222964
rect 371292 222924 398564 222952
rect 371292 222912 371298 222924
rect 398558 222912 398564 222924
rect 398616 222912 398622 222964
rect 399754 222912 399760 222964
rect 399812 222952 399818 222964
rect 543090 222952 543096 222964
rect 399812 222924 543096 222952
rect 399812 222912 399818 222924
rect 543090 222912 543096 222924
rect 543148 222912 543154 222964
rect 119982 222844 119988 222896
rect 120040 222884 120046 222896
rect 221458 222884 221464 222896
rect 120040 222856 221464 222884
rect 120040 222844 120046 222856
rect 221458 222844 221464 222856
rect 221516 222844 221522 222896
rect 224310 222844 224316 222896
rect 224368 222884 224374 222896
rect 246758 222884 246764 222896
rect 224368 222856 246764 222884
rect 224368 222844 224374 222856
rect 246758 222844 246764 222856
rect 246816 222844 246822 222896
rect 246850 222844 246856 222896
rect 246908 222884 246914 222896
rect 256694 222884 256700 222896
rect 246908 222856 256700 222884
rect 246908 222844 246914 222856
rect 256694 222844 256700 222856
rect 256752 222844 256758 222896
rect 257062 222844 257068 222896
rect 257120 222884 257126 222896
rect 278130 222884 278136 222896
rect 257120 222856 278136 222884
rect 257120 222844 257126 222856
rect 278130 222844 278136 222856
rect 278188 222844 278194 222896
rect 327350 222844 327356 222896
rect 327408 222884 327414 222896
rect 370038 222884 370044 222896
rect 327408 222856 370044 222884
rect 327408 222844 327414 222856
rect 370038 222844 370044 222856
rect 370096 222844 370102 222896
rect 371142 222844 371148 222896
rect 371200 222884 371206 222896
rect 400398 222884 400404 222896
rect 371200 222856 400404 222884
rect 371200 222844 371206 222856
rect 400398 222844 400404 222856
rect 400456 222844 400462 222896
rect 401870 222844 401876 222896
rect 401928 222884 401934 222896
rect 547506 222884 547512 222896
rect 401928 222856 547512 222884
rect 401928 222844 401934 222856
rect 547506 222844 547512 222856
rect 547564 222844 547570 222896
rect 565998 222844 566004 222896
rect 566056 222884 566062 222896
rect 620554 222884 620560 222896
rect 566056 222856 620560 222884
rect 566056 222844 566062 222856
rect 620554 222844 620560 222856
rect 620612 222844 620618 222896
rect 116578 222776 116584 222828
rect 116636 222816 116642 222828
rect 220078 222816 220084 222828
rect 116636 222788 220084 222816
rect 116636 222776 116642 222788
rect 220078 222776 220084 222788
rect 220136 222776 220142 222828
rect 222562 222776 222568 222828
rect 222620 222816 222626 222828
rect 257338 222816 257344 222828
rect 222620 222788 231854 222816
rect 222620 222776 222626 222788
rect 91370 222708 91376 222760
rect 91428 222748 91434 222760
rect 209038 222748 209044 222760
rect 91428 222720 209044 222748
rect 91428 222708 91434 222720
rect 209038 222708 209044 222720
rect 209096 222708 209102 222760
rect 231826 222748 231854 222788
rect 251146 222788 257344 222816
rect 251146 222748 251174 222788
rect 257338 222776 257344 222788
rect 257396 222776 257402 222828
rect 261294 222776 261300 222828
rect 261352 222816 261358 222828
rect 281350 222816 281356 222828
rect 261352 222788 281356 222816
rect 261352 222776 261358 222788
rect 281350 222776 281356 222788
rect 281408 222776 281414 222828
rect 330202 222776 330208 222828
rect 330260 222816 330266 222828
rect 376754 222816 376760 222828
rect 330260 222788 376760 222816
rect 330260 222776 330266 222788
rect 376754 222776 376760 222788
rect 376812 222776 376818 222828
rect 401502 222776 401508 222828
rect 401560 222816 401566 222828
rect 546678 222816 546684 222828
rect 401560 222788 546684 222816
rect 401560 222776 401566 222788
rect 546678 222776 546684 222788
rect 546736 222776 546742 222828
rect 549346 222776 549352 222828
rect 549404 222816 549410 222828
rect 551094 222816 551100 222828
rect 549404 222788 551100 222816
rect 549404 222776 549410 222788
rect 551094 222776 551100 222788
rect 551152 222816 551158 222828
rect 617794 222816 617800 222828
rect 551152 222788 617800 222816
rect 551152 222776 551158 222788
rect 617794 222776 617800 222788
rect 617852 222776 617858 222828
rect 258902 222748 258908 222760
rect 231826 222720 251174 222748
rect 256666 222720 258908 222748
rect 82170 222640 82176 222692
rect 82228 222680 82234 222692
rect 203978 222680 203984 222692
rect 82228 222652 203984 222680
rect 82228 222640 82234 222652
rect 203978 222640 203984 222652
rect 204036 222640 204042 222692
rect 215846 222640 215852 222692
rect 215904 222680 215910 222692
rect 246850 222680 246856 222692
rect 215904 222652 246856 222680
rect 215904 222640 215910 222652
rect 246850 222640 246856 222652
rect 246908 222640 246914 222692
rect 256666 222680 256694 222720
rect 258902 222708 258908 222720
rect 258960 222708 258966 222760
rect 262950 222708 262956 222760
rect 263008 222748 263014 222760
rect 281718 222748 281724 222760
rect 263008 222720 281724 222748
rect 263008 222708 263014 222720
rect 281718 222708 281724 222720
rect 281776 222708 281782 222760
rect 328086 222708 328092 222760
rect 328144 222748 328150 222760
rect 374178 222748 374184 222760
rect 328144 222720 374184 222748
rect 328144 222708 328150 222720
rect 374178 222708 374184 222720
rect 374236 222708 374242 222760
rect 402238 222708 402244 222760
rect 402296 222748 402302 222760
rect 548334 222748 548340 222760
rect 402296 222720 548340 222748
rect 402296 222708 402302 222720
rect 548334 222708 548340 222720
rect 548392 222708 548398 222760
rect 567930 222708 567936 222760
rect 567988 222748 567994 222760
rect 635458 222748 635464 222760
rect 567988 222720 635464 222748
rect 567988 222708 567994 222720
rect 635458 222708 635464 222720
rect 635516 222708 635522 222760
rect 246960 222652 256694 222680
rect 85482 222572 85488 222624
rect 85540 222612 85546 222624
rect 205450 222612 205456 222624
rect 85540 222584 205456 222612
rect 85540 222572 85546 222584
rect 205450 222572 205456 222584
rect 205508 222572 205514 222624
rect 209130 222572 209136 222624
rect 209188 222612 209194 222624
rect 246960 222612 246988 222652
rect 260466 222640 260472 222692
rect 260524 222680 260530 222692
rect 279602 222680 279608 222692
rect 260524 222652 279608 222680
rect 260524 222640 260530 222652
rect 279602 222640 279608 222652
rect 279660 222640 279666 222692
rect 329466 222640 329472 222692
rect 329524 222680 329530 222692
rect 377582 222680 377588 222692
rect 329524 222652 377588 222680
rect 329524 222640 329530 222652
rect 377582 222640 377588 222652
rect 377640 222640 377646 222692
rect 403618 222640 403624 222692
rect 403676 222680 403682 222692
rect 552014 222680 552020 222692
rect 403676 222652 552020 222680
rect 403676 222640 403682 222652
rect 552014 222640 552020 222652
rect 552072 222640 552078 222692
rect 568574 222640 568580 222692
rect 568632 222680 568638 222692
rect 621014 222680 621020 222692
rect 568632 222652 621020 222680
rect 568632 222640 568638 222652
rect 621014 222640 621020 222652
rect 621072 222640 621078 222692
rect 257522 222612 257528 222624
rect 209188 222584 246988 222612
rect 256666 222584 257528 222612
rect 209188 222572 209194 222584
rect 75362 222504 75368 222556
rect 75420 222544 75426 222556
rect 201126 222544 201132 222556
rect 75420 222516 201132 222544
rect 75420 222504 75426 222516
rect 201126 222504 201132 222516
rect 201184 222504 201190 222556
rect 205818 222504 205824 222556
rect 205876 222544 205882 222556
rect 256666 222544 256694 222584
rect 257522 222572 257528 222584
rect 257580 222572 257586 222624
rect 262122 222572 262128 222624
rect 262180 222612 262186 222624
rect 280706 222612 280712 222624
rect 262180 222584 280712 222612
rect 262180 222572 262186 222584
rect 280706 222572 280712 222584
rect 280764 222572 280770 222624
rect 284938 222612 284944 222624
rect 282932 222584 284944 222612
rect 205876 222516 246988 222544
rect 205876 222504 205882 222516
rect 68646 222436 68652 222488
rect 68704 222476 68710 222488
rect 198274 222476 198280 222488
rect 68704 222448 198280 222476
rect 68704 222436 68710 222448
rect 198274 222436 198280 222448
rect 198332 222436 198338 222488
rect 202414 222436 202420 222488
rect 202472 222476 202478 222488
rect 246666 222476 246672 222488
rect 202472 222448 246672 222476
rect 202472 222436 202478 222448
rect 246666 222436 246672 222448
rect 246724 222436 246730 222488
rect 53558 222368 53564 222420
rect 53616 222408 53622 222420
rect 182174 222408 182180 222420
rect 53616 222380 182180 222408
rect 53616 222368 53622 222380
rect 182174 222368 182180 222380
rect 182232 222368 182238 222420
rect 188982 222368 188988 222420
rect 189040 222408 189046 222420
rect 246960 222408 246988 222516
rect 247236 222516 256694 222544
rect 247236 222408 247264 222516
rect 264606 222504 264612 222556
rect 264664 222544 264670 222556
rect 282822 222544 282828 222556
rect 264664 222516 282828 222544
rect 264664 222504 264670 222516
rect 282822 222504 282828 222516
rect 282880 222504 282886 222556
rect 249518 222436 249524 222488
rect 249576 222476 249582 222488
rect 259362 222476 259368 222488
rect 249576 222448 259368 222476
rect 249576 222436 249582 222448
rect 259362 222436 259368 222448
rect 259420 222436 259426 222488
rect 272242 222436 272248 222488
rect 272300 222476 272306 222488
rect 282932 222476 282960 222584
rect 284938 222572 284944 222584
rect 284996 222572 285002 222624
rect 331582 222572 331588 222624
rect 331640 222612 331646 222624
rect 378410 222612 378416 222624
rect 331640 222584 378416 222612
rect 331640 222572 331646 222584
rect 378410 222572 378416 222584
rect 378468 222572 378474 222624
rect 405826 222572 405832 222624
rect 405884 222612 405890 222624
rect 556706 222612 556712 222624
rect 405884 222584 556712 222612
rect 405884 222572 405890 222584
rect 556706 222572 556712 222584
rect 556764 222572 556770 222624
rect 557442 222572 557448 222624
rect 557500 222612 557506 222624
rect 618714 222612 618720 222624
rect 557500 222584 618720 222612
rect 557500 222572 557506 222584
rect 618714 222572 618720 222584
rect 618772 222572 618778 222624
rect 283190 222504 283196 222556
rect 283248 222544 283254 222556
rect 290274 222544 290280 222556
rect 283248 222516 290280 222544
rect 283248 222504 283254 222516
rect 290274 222504 290280 222516
rect 290332 222504 290338 222556
rect 343634 222544 343640 222556
rect 333946 222516 343640 222544
rect 272300 222448 282960 222476
rect 272300 222436 272306 222448
rect 325234 222436 325240 222488
rect 325292 222476 325298 222488
rect 333946 222476 333974 222516
rect 343634 222504 343640 222516
rect 343692 222504 343698 222556
rect 343726 222504 343732 222556
rect 343784 222544 343790 222556
rect 375374 222544 375380 222556
rect 343784 222516 375380 222544
rect 343784 222504 343790 222516
rect 375374 222504 375380 222516
rect 375432 222504 375438 222556
rect 380986 222504 380992 222556
rect 381044 222544 381050 222556
rect 394694 222544 394700 222556
rect 381044 222516 394700 222544
rect 381044 222504 381050 222516
rect 394694 222504 394700 222516
rect 394752 222504 394758 222556
rect 403986 222504 403992 222556
rect 404044 222544 404050 222556
rect 552106 222544 552112 222556
rect 404044 222516 552112 222544
rect 404044 222504 404050 222516
rect 552106 222504 552112 222516
rect 552164 222504 552170 222556
rect 556522 222504 556528 222556
rect 556580 222544 556586 222556
rect 557460 222544 557488 222572
rect 556580 222516 557488 222544
rect 556580 222504 556586 222516
rect 561214 222504 561220 222556
rect 561272 222544 561278 222556
rect 561272 222516 563560 222544
rect 561272 222504 561278 222516
rect 372614 222476 372620 222488
rect 325292 222448 333974 222476
rect 341812 222448 372620 222476
rect 325292 222436 325298 222448
rect 189040 222380 243860 222408
rect 246960 222380 247264 222408
rect 189040 222368 189046 222380
rect 66162 222300 66168 222352
rect 66220 222340 66226 222352
rect 198642 222340 198648 222352
rect 66220 222312 198648 222340
rect 66220 222300 66226 222312
rect 198642 222300 198648 222312
rect 198700 222300 198706 222352
rect 200758 222300 200764 222352
rect 200816 222340 200822 222352
rect 243722 222340 243728 222352
rect 200816 222312 243728 222340
rect 200816 222300 200822 222312
rect 243722 222300 243728 222312
rect 243780 222300 243786 222352
rect 243832 222340 243860 222380
rect 247862 222368 247868 222420
rect 247920 222408 247926 222420
rect 254394 222408 254400 222420
rect 247920 222380 254400 222408
rect 247920 222368 247926 222380
rect 254394 222368 254400 222380
rect 254452 222368 254458 222420
rect 254578 222368 254584 222420
rect 254636 222408 254642 222420
rect 278498 222408 278504 222420
rect 254636 222380 278504 222408
rect 254636 222368 254642 222380
rect 278498 222368 278504 222380
rect 278556 222368 278562 222420
rect 327718 222368 327724 222420
rect 327776 222408 327782 222420
rect 341812 222408 341840 222448
rect 372614 222436 372620 222448
rect 372672 222436 372678 222488
rect 382274 222436 382280 222488
rect 382332 222476 382338 222488
rect 396258 222476 396264 222488
rect 382332 222448 396264 222476
rect 382332 222436 382338 222448
rect 396258 222436 396264 222448
rect 396316 222436 396322 222488
rect 406470 222436 406476 222488
rect 406528 222476 406534 222488
rect 558822 222476 558828 222488
rect 406528 222448 558828 222476
rect 406528 222436 406534 222448
rect 558822 222436 558828 222448
rect 558880 222476 558886 222488
rect 560202 222476 560208 222488
rect 558880 222448 560208 222476
rect 558880 222436 558886 222448
rect 560202 222436 560208 222448
rect 560260 222436 560266 222488
rect 560386 222436 560392 222488
rect 560444 222476 560450 222488
rect 560444 222448 563468 222476
rect 560444 222436 560450 222448
rect 327776 222380 341840 222408
rect 327776 222368 327782 222380
rect 343542 222368 343548 222420
rect 343600 222408 343606 222420
rect 375926 222408 375932 222420
rect 343600 222380 375932 222408
rect 343600 222368 343606 222380
rect 375926 222368 375932 222380
rect 375984 222368 375990 222420
rect 378134 222368 378140 222420
rect 378192 222408 378198 222420
rect 397730 222408 397736 222420
rect 378192 222380 397736 222408
rect 378192 222368 378198 222380
rect 397730 222368 397736 222380
rect 397788 222368 397794 222420
rect 406194 222368 406200 222420
rect 406252 222368 406258 222420
rect 407942 222368 407948 222420
rect 408000 222408 408006 222420
rect 561766 222408 561772 222420
rect 408000 222380 561772 222408
rect 408000 222368 408006 222380
rect 561766 222368 561772 222380
rect 561824 222368 561830 222420
rect 250070 222340 250076 222352
rect 243832 222312 250076 222340
rect 250070 222300 250076 222312
rect 250128 222300 250134 222352
rect 259362 222300 259368 222352
rect 259420 222340 259426 222352
rect 280338 222340 280344 222352
rect 259420 222312 280344 222340
rect 259420 222300 259426 222312
rect 280338 222300 280344 222312
rect 280396 222300 280402 222352
rect 310974 222300 310980 222352
rect 311032 222340 311038 222352
rect 333974 222340 333980 222352
rect 311032 222312 333980 222340
rect 311032 222300 311038 222312
rect 333974 222300 333980 222312
rect 334032 222300 334038 222352
rect 339770 222300 339776 222352
rect 339828 222340 339834 222352
rect 349798 222340 349804 222352
rect 339828 222312 349804 222340
rect 339828 222300 339834 222312
rect 349798 222300 349804 222312
rect 349856 222300 349862 222352
rect 349890 222300 349896 222352
rect 349948 222340 349954 222352
rect 385126 222340 385132 222352
rect 349948 222312 385132 222340
rect 349948 222300 349954 222312
rect 385126 222300 385132 222312
rect 385184 222300 385190 222352
rect 385218 222300 385224 222352
rect 385276 222340 385282 222352
rect 402974 222340 402980 222352
rect 385276 222312 402980 222340
rect 385276 222300 385282 222312
rect 402974 222300 402980 222312
rect 403032 222300 403038 222352
rect 406212 222340 406240 222368
rect 557534 222340 557540 222352
rect 406212 222312 557540 222340
rect 557534 222300 557540 222312
rect 557592 222300 557598 222352
rect 563440 222340 563468 222448
rect 563532 222408 563560 222516
rect 563698 222436 563704 222488
rect 563756 222476 563762 222488
rect 620094 222476 620100 222488
rect 563756 222448 620100 222476
rect 563756 222436 563762 222448
rect 620094 222436 620100 222448
rect 620152 222436 620158 222488
rect 619634 222408 619640 222420
rect 563532 222380 619640 222408
rect 619634 222368 619640 222380
rect 619692 222368 619698 222420
rect 634078 222340 634084 222352
rect 563440 222312 634084 222340
rect 634078 222300 634084 222312
rect 634136 222300 634142 222352
rect 61930 222232 61936 222284
rect 61988 222272 61994 222284
rect 195422 222272 195428 222284
rect 61988 222244 195428 222272
rect 61988 222232 61994 222244
rect 195422 222232 195428 222244
rect 195480 222232 195486 222284
rect 195698 222232 195704 222284
rect 195756 222272 195762 222284
rect 253198 222272 253204 222284
rect 195756 222244 253204 222272
rect 195756 222232 195762 222244
rect 253198 222232 253204 222244
rect 253256 222232 253262 222284
rect 314194 222232 314200 222284
rect 314252 222272 314258 222284
rect 338022 222272 338028 222284
rect 314252 222244 338028 222272
rect 314252 222232 314258 222244
rect 338022 222232 338028 222244
rect 338080 222232 338086 222284
rect 338114 222232 338120 222284
rect 338172 222272 338178 222284
rect 346486 222272 346492 222284
rect 338172 222244 346492 222272
rect 338172 222232 338178 222244
rect 346486 222232 346492 222244
rect 346544 222232 346550 222284
rect 393590 222272 393596 222284
rect 346596 222244 393596 222272
rect 59170 222164 59176 222216
rect 59228 222204 59234 222216
rect 195790 222204 195796 222216
rect 59228 222176 195796 222204
rect 59228 222164 59234 222176
rect 195790 222164 195796 222176
rect 195848 222164 195854 222216
rect 207474 222164 207480 222216
rect 207532 222204 207538 222216
rect 246298 222204 246304 222216
rect 207532 222176 246304 222204
rect 207532 222164 207538 222176
rect 246298 222164 246304 222176
rect 246356 222164 246362 222216
rect 257890 222164 257896 222216
rect 257948 222204 257954 222216
rect 279970 222204 279976 222216
rect 257948 222176 279976 222204
rect 257948 222164 257954 222176
rect 279970 222164 279976 222176
rect 280028 222164 280034 222216
rect 281442 222164 281448 222216
rect 281500 222204 281506 222216
rect 289906 222204 289912 222216
rect 281500 222176 289912 222204
rect 281500 222164 281506 222176
rect 289906 222164 289912 222176
rect 289964 222164 289970 222216
rect 313090 222164 313096 222216
rect 313148 222204 313154 222216
rect 336734 222204 336740 222216
rect 313148 222176 336740 222204
rect 313148 222164 313154 222176
rect 336734 222164 336740 222176
rect 336792 222164 336798 222216
rect 337378 222164 337384 222216
rect 337436 222204 337442 222216
rect 346596 222204 346624 222244
rect 393590 222232 393596 222244
rect 393648 222232 393654 222284
rect 394602 222232 394608 222284
rect 394660 222272 394666 222284
rect 406194 222272 406200 222284
rect 394660 222244 406200 222272
rect 394660 222232 394666 222244
rect 406194 222232 406200 222244
rect 406252 222232 406258 222284
rect 408126 222232 408132 222284
rect 408184 222272 408190 222284
rect 562870 222272 562876 222284
rect 408184 222244 562876 222272
rect 408184 222232 408190 222244
rect 562870 222232 562876 222244
rect 562928 222232 562934 222284
rect 565446 222232 565452 222284
rect 565504 222272 565510 222284
rect 634998 222272 635004 222284
rect 565504 222244 635004 222272
rect 565504 222232 565510 222244
rect 634998 222232 635004 222244
rect 635056 222232 635062 222284
rect 337436 222176 346624 222204
rect 337436 222164 337442 222176
rect 346670 222164 346676 222216
rect 346728 222204 346734 222216
rect 391934 222204 391940 222216
rect 346728 222176 391940 222204
rect 346728 222164 346734 222176
rect 391934 222164 391940 222176
rect 391992 222164 391998 222216
rect 397638 222164 397644 222216
rect 397696 222204 397702 222216
rect 401962 222204 401968 222216
rect 397696 222176 401968 222204
rect 397696 222164 397702 222176
rect 401962 222164 401968 222176
rect 402020 222164 402026 222216
rect 410886 222164 410892 222216
rect 410944 222204 410950 222216
rect 569310 222204 569316 222216
rect 410944 222176 569316 222204
rect 410944 222164 410950 222176
rect 569310 222164 569316 222176
rect 569368 222164 569374 222216
rect 652846 222164 652852 222216
rect 652904 222204 652910 222216
rect 674650 222204 674656 222216
rect 652904 222176 674656 222204
rect 652904 222164 652910 222176
rect 674650 222164 674656 222176
rect 674708 222204 674714 222216
rect 675754 222204 675760 222216
rect 674708 222176 675760 222204
rect 674708 222164 674714 222176
rect 675754 222164 675760 222176
rect 675812 222164 675818 222216
rect 155310 222096 155316 222148
rect 155368 222136 155374 222148
rect 235810 222136 235816 222148
rect 155368 222108 235816 222136
rect 155368 222096 155374 222108
rect 235810 222096 235816 222108
rect 235868 222096 235874 222148
rect 244642 222136 244648 222148
rect 237346 222108 244648 222136
rect 93762 222028 93768 222080
rect 93820 222068 93826 222080
rect 155862 222068 155868 222080
rect 93820 222040 155868 222068
rect 93820 222028 93826 222040
rect 155862 222028 155868 222040
rect 155920 222028 155926 222080
rect 232590 222028 232596 222080
rect 232648 222068 232654 222080
rect 237346 222068 237374 222108
rect 244642 222096 244648 222108
rect 244700 222096 244706 222148
rect 251082 222096 251088 222148
rect 251140 222136 251146 222148
rect 254210 222136 254216 222148
rect 251140 222108 254216 222136
rect 251140 222096 251146 222108
rect 254210 222096 254216 222108
rect 254268 222096 254274 222148
rect 273070 222096 273076 222148
rect 273128 222136 273134 222148
rect 286042 222136 286048 222148
rect 273128 222108 286048 222136
rect 273128 222096 273134 222108
rect 286042 222096 286048 222108
rect 286100 222096 286106 222148
rect 321646 222096 321652 222148
rect 321704 222136 321710 222148
rect 356514 222136 356520 222148
rect 321704 222108 356520 222136
rect 321704 222096 321710 222108
rect 356514 222096 356520 222108
rect 356572 222096 356578 222148
rect 383010 222096 383016 222148
rect 383068 222136 383074 222148
rect 503530 222136 503536 222148
rect 383068 222108 503536 222136
rect 383068 222096 383074 222108
rect 503530 222096 503536 222108
rect 503588 222096 503594 222148
rect 538858 222096 538864 222148
rect 538916 222136 538922 222148
rect 615494 222136 615500 222148
rect 538916 222108 615500 222136
rect 538916 222096 538922 222108
rect 615494 222096 615500 222108
rect 615552 222096 615558 222148
rect 238294 222068 238300 222080
rect 232648 222040 237374 222068
rect 237668 222040 238300 222068
rect 232648 222028 232654 222040
rect 160370 221960 160376 222012
rect 160428 222000 160434 222012
rect 237668 222000 237696 222040
rect 238294 222028 238300 222040
rect 238352 222028 238358 222080
rect 243722 222028 243728 222080
rect 243780 222068 243786 222080
rect 255682 222068 255688 222080
rect 243780 222040 255688 222068
rect 243780 222028 243786 222040
rect 255682 222028 255688 222040
rect 255740 222028 255746 222080
rect 320910 222028 320916 222080
rect 320968 222068 320974 222080
rect 357342 222068 357348 222080
rect 320968 222040 357348 222068
rect 320968 222028 320974 222040
rect 357342 222028 357348 222040
rect 357400 222028 357406 222080
rect 384390 222028 384396 222080
rect 384448 222068 384454 222080
rect 506290 222068 506296 222080
rect 384448 222040 506296 222068
rect 384448 222028 384454 222040
rect 506290 222028 506296 222040
rect 506348 222028 506354 222080
rect 555050 222028 555056 222080
rect 555108 222068 555114 222080
rect 633158 222068 633164 222080
rect 555108 222040 633164 222068
rect 555108 222028 555114 222040
rect 633158 222028 633164 222040
rect 633216 222028 633222 222080
rect 160428 221972 237696 222000
rect 160428 221960 160434 221972
rect 237742 221960 237748 222012
rect 237800 222000 237806 222012
rect 251266 222000 251272 222012
rect 237800 221972 251272 222000
rect 237800 221960 237806 221972
rect 251266 221960 251272 221972
rect 251324 221960 251330 222012
rect 322750 221960 322756 222012
rect 322808 222000 322814 222012
rect 358262 222000 358268 222012
rect 322808 221972 358268 222000
rect 322808 221960 322814 221972
rect 358262 221960 358268 221972
rect 358320 221960 358326 222012
rect 380526 221960 380532 222012
rect 380584 222000 380590 222012
rect 497366 222000 497372 222012
rect 380584 221972 497372 222000
rect 380584 221960 380590 221972
rect 497366 221960 497372 221972
rect 497424 222000 497430 222012
rect 499022 222000 499028 222012
rect 497424 221972 499028 222000
rect 497424 221960 497430 221972
rect 499022 221960 499028 221972
rect 499080 221960 499086 222012
rect 552106 221960 552112 222012
rect 552164 222000 552170 222012
rect 552842 222000 552848 222012
rect 552164 221972 552848 222000
rect 552164 221960 552170 221972
rect 552842 221960 552848 221972
rect 552900 222000 552906 222012
rect 632698 222000 632704 222012
rect 552900 221972 632704 222000
rect 552900 221960 552906 221972
rect 632698 221960 632704 221972
rect 632756 221960 632762 222012
rect 170490 221892 170496 221944
rect 170548 221932 170554 221944
rect 242894 221932 242900 221944
rect 170548 221904 242900 221932
rect 170548 221892 170554 221904
rect 242894 221892 242900 221904
rect 242952 221892 242958 221944
rect 319806 221892 319812 221944
rect 319864 221932 319870 221944
rect 354030 221932 354036 221944
rect 319864 221904 354036 221932
rect 319864 221892 319870 221904
rect 354030 221892 354036 221904
rect 354088 221892 354094 221944
rect 387518 221892 387524 221944
rect 387576 221932 387582 221944
rect 396166 221932 396172 221944
rect 387576 221904 396172 221932
rect 387576 221892 387582 221904
rect 396166 221892 396172 221904
rect 396224 221892 396230 221944
rect 396258 221892 396264 221944
rect 396316 221932 396322 221944
rect 501230 221932 501236 221944
rect 396316 221904 501236 221932
rect 396316 221892 396322 221904
rect 501230 221892 501236 221904
rect 501288 221892 501294 221944
rect 532786 221892 532792 221944
rect 532844 221932 532850 221944
rect 533430 221932 533436 221944
rect 532844 221904 533436 221932
rect 532844 221892 532850 221904
rect 533430 221892 533436 221904
rect 533488 221932 533494 221944
rect 614574 221932 614580 221944
rect 533488 221904 614580 221932
rect 533488 221892 533494 221904
rect 614574 221892 614580 221904
rect 614632 221892 614638 221944
rect 168742 221824 168748 221876
rect 168800 221864 168806 221876
rect 241790 221864 241796 221876
rect 168800 221836 241796 221864
rect 168800 221824 168806 221836
rect 241790 221824 241796 221836
rect 241848 221824 241854 221876
rect 244458 221824 244464 221876
rect 244516 221864 244522 221876
rect 254118 221864 254124 221876
rect 244516 221836 254124 221864
rect 244516 221824 244522 221836
rect 254118 221824 254124 221836
rect 254176 221824 254182 221876
rect 274726 221824 274732 221876
rect 274784 221864 274790 221876
rect 287054 221864 287060 221876
rect 274784 221836 287060 221864
rect 274784 221824 274790 221836
rect 287054 221824 287060 221836
rect 287112 221824 287118 221876
rect 287146 221824 287152 221876
rect 287204 221864 287210 221876
rect 289262 221864 289268 221876
rect 287204 221836 289268 221864
rect 287204 221824 287210 221836
rect 289262 221824 289268 221836
rect 289320 221824 289326 221876
rect 318058 221824 318064 221876
rect 318116 221864 318122 221876
rect 350626 221864 350632 221876
rect 318116 221836 350632 221864
rect 318116 221824 318122 221836
rect 350626 221824 350632 221836
rect 350684 221824 350690 221876
rect 377950 221824 377956 221876
rect 378008 221864 378014 221876
rect 491294 221864 491300 221876
rect 378008 221836 491300 221864
rect 378008 221824 378014 221836
rect 491294 221824 491300 221836
rect 491352 221824 491358 221876
rect 547506 221824 547512 221876
rect 547564 221864 547570 221876
rect 631778 221864 631784 221876
rect 547564 221836 631784 221864
rect 547564 221824 547570 221836
rect 631778 221824 631784 221836
rect 631836 221824 631842 221876
rect 175458 221756 175464 221808
rect 175516 221796 175522 221808
rect 232590 221796 232596 221808
rect 175516 221768 232596 221796
rect 175516 221756 175522 221768
rect 232590 221756 232596 221768
rect 232648 221756 232654 221808
rect 234338 221756 234344 221808
rect 234396 221796 234402 221808
rect 248598 221796 248604 221808
rect 234396 221768 248604 221796
rect 234396 221756 234402 221768
rect 248598 221756 248604 221768
rect 248656 221756 248662 221808
rect 255406 221756 255412 221808
rect 255464 221796 255470 221808
rect 277854 221796 277860 221808
rect 255464 221768 277860 221796
rect 255464 221756 255470 221768
rect 277854 221756 277860 221768
rect 277912 221756 277918 221808
rect 285306 221796 285312 221808
rect 279344 221768 285312 221796
rect 182082 221688 182088 221740
rect 182140 221728 182146 221740
rect 182140 221700 235948 221728
rect 182140 221688 182146 221700
rect 183922 221620 183928 221672
rect 183980 221660 183986 221672
rect 235920 221660 235948 221700
rect 239398 221688 239404 221740
rect 239456 221728 239462 221740
rect 254302 221728 254308 221740
rect 239456 221700 254308 221728
rect 239456 221688 239462 221700
rect 254302 221688 254308 221700
rect 254360 221688 254366 221740
rect 258810 221688 258816 221740
rect 258868 221728 258874 221740
rect 279234 221728 279240 221740
rect 258868 221700 279240 221728
rect 258868 221688 258874 221700
rect 279234 221688 279240 221700
rect 279292 221688 279298 221740
rect 240962 221660 240968 221672
rect 183980 221632 235810 221660
rect 235920 221632 240968 221660
rect 183980 221620 183986 221632
rect 183094 221552 183100 221604
rect 183152 221592 183158 221604
rect 235626 221592 235632 221604
rect 183152 221564 235632 221592
rect 183152 221552 183158 221564
rect 235626 221552 235632 221564
rect 235684 221552 235690 221604
rect 159542 221484 159548 221536
rect 159600 221524 159606 221536
rect 209590 221524 209596 221536
rect 159600 221496 209596 221524
rect 159600 221484 159606 221496
rect 209590 221484 209596 221496
rect 209648 221484 209654 221536
rect 214190 221484 214196 221536
rect 214248 221524 214254 221536
rect 235782 221524 235810 221632
rect 240962 221620 240968 221632
rect 241020 221620 241026 221672
rect 246574 221660 246580 221672
rect 241072 221632 246580 221660
rect 235902 221552 235908 221604
rect 235960 221592 235966 221604
rect 241072 221592 241100 221632
rect 246574 221620 246580 221632
rect 246632 221620 246638 221672
rect 273898 221620 273904 221672
rect 273956 221660 273962 221672
rect 279344 221660 279372 221768
rect 285306 221756 285312 221768
rect 285364 221756 285370 221808
rect 321278 221756 321284 221808
rect 321336 221796 321342 221808
rect 354858 221796 354864 221808
rect 321336 221768 354864 221796
rect 321336 221756 321342 221768
rect 354858 221756 354864 221768
rect 354916 221756 354922 221808
rect 379422 221756 379428 221808
rect 379480 221796 379486 221808
rect 494514 221796 494520 221808
rect 379480 221768 494520 221796
rect 379480 221756 379486 221768
rect 494514 221756 494520 221768
rect 494572 221756 494578 221808
rect 530670 221756 530676 221808
rect 530728 221796 530734 221808
rect 614022 221796 614028 221808
rect 530728 221768 614028 221796
rect 530728 221756 530734 221768
rect 614022 221756 614028 221768
rect 614080 221756 614086 221808
rect 283926 221688 283932 221740
rect 283984 221728 283990 221740
rect 289538 221728 289544 221740
rect 283984 221700 289544 221728
rect 283984 221688 283990 221700
rect 289538 221688 289544 221700
rect 289596 221688 289602 221740
rect 319898 221688 319904 221740
rect 319956 221728 319962 221740
rect 351454 221728 351460 221740
rect 319956 221700 351460 221728
rect 319956 221688 319962 221700
rect 351454 221688 351460 221700
rect 351512 221688 351518 221740
rect 377674 221688 377680 221740
rect 377732 221728 377738 221740
rect 490282 221728 490288 221740
rect 377732 221700 490288 221728
rect 377732 221688 377738 221700
rect 490282 221688 490288 221700
rect 490340 221688 490346 221740
rect 545206 221688 545212 221740
rect 545264 221728 545270 221740
rect 631318 221728 631324 221740
rect 545264 221700 631324 221728
rect 545264 221688 545270 221700
rect 631318 221688 631324 221700
rect 631376 221688 631382 221740
rect 273956 221632 279372 221660
rect 273956 221620 273962 221632
rect 287054 221620 287060 221672
rect 287112 221660 287118 221672
rect 288526 221660 288532 221672
rect 287112 221632 288532 221660
rect 287112 221620 287118 221632
rect 288526 221620 288532 221632
rect 288584 221620 288590 221672
rect 316678 221620 316684 221672
rect 316736 221660 316742 221672
rect 347314 221660 347320 221672
rect 316736 221632 347320 221660
rect 316736 221620 316742 221632
rect 347314 221620 347320 221632
rect 347372 221620 347378 221672
rect 351914 221620 351920 221672
rect 351972 221660 351978 221672
rect 383746 221660 383752 221672
rect 351972 221632 383752 221660
rect 351972 221620 351978 221632
rect 383746 221620 383752 221632
rect 383804 221620 383810 221672
rect 383838 221620 383844 221672
rect 383896 221660 383902 221672
rect 396074 221660 396080 221672
rect 383896 221632 396080 221660
rect 383896 221620 383902 221632
rect 396074 221620 396080 221632
rect 396132 221620 396138 221672
rect 396166 221620 396172 221672
rect 396224 221660 396230 221672
rect 494146 221660 494152 221672
rect 396224 221632 494152 221660
rect 396224 221620 396230 221632
rect 494146 221620 494152 221632
rect 494204 221660 494210 221672
rect 495802 221660 495808 221672
rect 494204 221632 495808 221660
rect 494204 221620 494210 221632
rect 495802 221620 495808 221632
rect 495860 221620 495866 221672
rect 528370 221620 528376 221672
rect 528428 221660 528434 221672
rect 613562 221660 613568 221672
rect 528428 221632 613568 221660
rect 528428 221620 528434 221632
rect 613562 221620 613568 221632
rect 613620 221620 613626 221672
rect 235960 221564 241100 221592
rect 235960 221552 235966 221564
rect 241146 221552 241152 221604
rect 241204 221592 241210 221604
rect 251174 221592 251180 221604
rect 241204 221564 251180 221592
rect 241204 221552 241210 221564
rect 251174 221552 251180 221564
rect 251232 221552 251238 221604
rect 268838 221552 268844 221604
rect 268896 221592 268902 221604
rect 283558 221592 283564 221604
rect 268896 221564 283564 221592
rect 268896 221552 268902 221564
rect 283558 221552 283564 221564
rect 283616 221552 283622 221604
rect 313826 221552 313832 221604
rect 313884 221592 313890 221604
rect 340598 221592 340604 221604
rect 313884 221564 340604 221592
rect 313884 221552 313890 221564
rect 340598 221552 340604 221564
rect 340656 221552 340662 221604
rect 345382 221552 345388 221604
rect 345440 221592 345446 221604
rect 373350 221592 373356 221604
rect 345440 221564 373356 221592
rect 345440 221552 345446 221564
rect 373350 221552 373356 221564
rect 373408 221552 373414 221604
rect 375466 221552 375472 221604
rect 375524 221592 375530 221604
rect 484394 221592 484400 221604
rect 375524 221564 484400 221592
rect 375524 221552 375530 221564
rect 484394 221552 484400 221564
rect 484452 221552 484458 221604
rect 543090 221552 543096 221604
rect 543148 221592 543154 221604
rect 630858 221592 630864 221604
rect 543148 221564 630864 221592
rect 543148 221552 543154 221564
rect 630858 221552 630864 221564
rect 630916 221552 630922 221604
rect 214248 221496 233740 221524
rect 235782 221496 240916 221524
rect 214248 221484 214254 221496
rect 166258 221416 166264 221468
rect 166316 221456 166322 221468
rect 215202 221456 215208 221468
rect 166316 221428 215208 221456
rect 166316 221416 166322 221428
rect 215202 221416 215208 221428
rect 215260 221416 215266 221468
rect 220078 221416 220084 221468
rect 220136 221456 220142 221468
rect 233712 221456 233740 221496
rect 240888 221456 240916 221496
rect 240962 221484 240968 221536
rect 241020 221524 241026 221536
rect 247494 221524 247500 221536
rect 241020 221496 247500 221524
rect 241020 221484 241026 221496
rect 247494 221484 247500 221496
rect 247552 221484 247558 221536
rect 270402 221484 270408 221536
rect 270460 221524 270466 221536
rect 283834 221524 283840 221536
rect 270460 221496 283840 221524
rect 270460 221484 270466 221496
rect 283834 221484 283840 221496
rect 283892 221484 283898 221536
rect 284846 221484 284852 221536
rect 284904 221524 284910 221536
rect 291378 221524 291384 221536
rect 284904 221496 291384 221524
rect 284904 221484 284910 221496
rect 291378 221484 291384 221496
rect 291436 221484 291442 221536
rect 317046 221484 317052 221536
rect 317104 221524 317110 221536
rect 345014 221524 345020 221536
rect 317104 221496 345020 221524
rect 317104 221484 317110 221496
rect 345014 221484 345020 221496
rect 345072 221484 345078 221536
rect 345106 221484 345112 221536
rect 345164 221524 345170 221536
rect 366634 221524 366640 221536
rect 345164 221496 366640 221524
rect 345164 221484 345170 221496
rect 366634 221484 366640 221496
rect 366692 221484 366698 221536
rect 374454 221484 374460 221536
rect 374512 221524 374518 221536
rect 480990 221524 480996 221536
rect 374512 221496 480996 221524
rect 374512 221484 374518 221496
rect 480990 221484 480996 221496
rect 481048 221484 481054 221536
rect 532694 221484 532700 221536
rect 532752 221524 532758 221536
rect 532970 221524 532976 221536
rect 532752 221496 532976 221524
rect 532752 221484 532758 221496
rect 532970 221484 532976 221496
rect 533028 221524 533034 221536
rect 628926 221524 628932 221536
rect 533028 221496 628932 221524
rect 533028 221484 533034 221496
rect 628926 221484 628932 221496
rect 628984 221484 628990 221536
rect 248782 221456 248788 221468
rect 220136 221428 230980 221456
rect 233712 221428 240824 221456
rect 240888 221428 248788 221456
rect 220136 221416 220142 221428
rect 187234 221348 187240 221400
rect 187292 221388 187298 221400
rect 230290 221388 230296 221400
rect 187292 221360 230296 221388
rect 187292 221348 187298 221360
rect 230290 221348 230296 221360
rect 230348 221348 230354 221400
rect 230952 221388 230980 221428
rect 235534 221388 235540 221400
rect 230952 221360 235540 221388
rect 235534 221348 235540 221360
rect 235592 221348 235598 221400
rect 236914 221348 236920 221400
rect 236972 221388 236978 221400
rect 240686 221388 240692 221400
rect 236972 221360 240692 221388
rect 236972 221348 236978 221360
rect 240686 221348 240692 221360
rect 240744 221348 240750 221400
rect 240796 221388 240824 221428
rect 248782 221416 248788 221428
rect 248840 221416 248846 221468
rect 275554 221416 275560 221468
rect 275612 221456 275618 221468
rect 286410 221456 286416 221468
rect 275612 221428 286416 221456
rect 275612 221416 275618 221428
rect 286410 221416 286416 221428
rect 286468 221416 286474 221468
rect 286502 221416 286508 221468
rect 286560 221456 286566 221468
rect 291746 221456 291752 221468
rect 286560 221428 291752 221456
rect 286560 221416 286566 221428
rect 291746 221416 291752 221428
rect 291804 221416 291810 221468
rect 315206 221416 315212 221468
rect 315264 221456 315270 221468
rect 343910 221456 343916 221468
rect 315264 221428 343916 221456
rect 315264 221416 315270 221428
rect 343910 221416 343916 221428
rect 343968 221416 343974 221468
rect 345290 221416 345296 221468
rect 345348 221456 345354 221468
rect 363230 221456 363236 221468
rect 345348 221428 363236 221456
rect 345348 221416 345354 221428
rect 363230 221416 363236 221428
rect 363288 221416 363294 221468
rect 368750 221416 368756 221468
rect 368808 221456 368814 221468
rect 467558 221456 467564 221468
rect 368808 221428 467564 221456
rect 368808 221416 368814 221428
rect 467558 221416 467564 221428
rect 467616 221416 467622 221468
rect 535454 221416 535460 221468
rect 535512 221456 535518 221468
rect 538030 221456 538036 221468
rect 535512 221428 538036 221456
rect 535512 221416 535518 221428
rect 538030 221416 538036 221428
rect 538088 221456 538094 221468
rect 629938 221456 629944 221468
rect 538088 221428 629944 221456
rect 538088 221416 538094 221428
rect 629938 221416 629944 221428
rect 629996 221416 630002 221468
rect 246942 221388 246948 221400
rect 240796 221360 246948 221388
rect 246942 221348 246948 221360
rect 247000 221348 247006 221400
rect 256234 221348 256240 221400
rect 256292 221388 256298 221400
rect 261478 221388 261484 221400
rect 256292 221360 261484 221388
rect 256292 221348 256298 221360
rect 261478 221348 261484 221360
rect 261536 221348 261542 221400
rect 267182 221348 267188 221400
rect 267240 221388 267246 221400
rect 282454 221388 282460 221400
rect 267240 221360 282460 221388
rect 267240 221348 267246 221360
rect 282454 221348 282460 221360
rect 282512 221348 282518 221400
rect 289078 221348 289084 221400
rect 289136 221388 289142 221400
rect 292114 221388 292120 221400
rect 289136 221360 292120 221388
rect 289136 221348 289142 221360
rect 292114 221348 292120 221360
rect 292172 221348 292178 221400
rect 292390 221348 292396 221400
rect 292448 221388 292454 221400
rect 293494 221388 293500 221400
rect 292448 221360 293500 221388
rect 292448 221348 292454 221360
rect 293494 221348 293500 221360
rect 293552 221348 293558 221400
rect 314562 221348 314568 221400
rect 314620 221388 314626 221400
rect 339678 221388 339684 221400
rect 314620 221360 339684 221388
rect 314620 221348 314626 221360
rect 339678 221348 339684 221360
rect 339736 221348 339742 221400
rect 342806 221348 342812 221400
rect 342864 221388 342870 221400
rect 359918 221388 359924 221400
rect 342864 221360 359924 221388
rect 342864 221348 342870 221360
rect 359918 221348 359924 221360
rect 359976 221348 359982 221400
rect 365898 221348 365904 221400
rect 365956 221388 365962 221400
rect 460934 221388 460940 221400
rect 365956 221360 460940 221388
rect 365956 221348 365962 221360
rect 460934 221348 460940 221360
rect 460992 221348 460998 221400
rect 507946 221348 507952 221400
rect 508004 221388 508010 221400
rect 609882 221388 609888 221400
rect 508004 221360 609888 221388
rect 508004 221348 508010 221360
rect 609882 221348 609888 221360
rect 609940 221348 609946 221400
rect 172974 221280 172980 221332
rect 173032 221320 173038 221332
rect 213086 221320 213092 221332
rect 173032 221292 213092 221320
rect 173032 221280 173038 221292
rect 213086 221280 213092 221292
rect 213144 221280 213150 221332
rect 233510 221280 233516 221332
rect 233568 221320 233574 221332
rect 239858 221320 239864 221332
rect 233568 221292 239864 221320
rect 233568 221280 233574 221292
rect 239858 221280 239864 221292
rect 239916 221280 239922 221332
rect 280614 221280 280620 221332
rect 280672 221320 280678 221332
rect 288158 221320 288164 221332
rect 280672 221292 288164 221320
rect 280672 221280 280678 221292
rect 288158 221280 288164 221292
rect 288216 221280 288222 221332
rect 289722 221280 289728 221332
rect 289780 221320 289786 221332
rect 293126 221320 293132 221332
rect 289780 221292 293132 221320
rect 289780 221280 289786 221292
rect 293126 221280 293132 221292
rect 293184 221280 293190 221332
rect 294966 221280 294972 221332
rect 295024 221320 295030 221332
rect 295610 221320 295616 221332
rect 295024 221292 295616 221320
rect 295024 221280 295030 221292
rect 295610 221280 295616 221292
rect 295668 221280 295674 221332
rect 315942 221280 315948 221332
rect 316000 221320 316006 221332
rect 343082 221320 343088 221332
rect 316000 221292 343088 221320
rect 316000 221280 316006 221292
rect 343082 221280 343088 221292
rect 343140 221280 343146 221332
rect 371510 221280 371516 221332
rect 371568 221320 371574 221332
rect 454126 221320 454132 221332
rect 371568 221292 454132 221320
rect 371568 221280 371574 221292
rect 454126 221280 454132 221292
rect 454184 221280 454190 221332
rect 510706 221280 510712 221332
rect 510764 221320 510770 221332
rect 610342 221320 610348 221332
rect 510764 221292 610348 221320
rect 510764 221280 510770 221292
rect 610342 221280 610348 221292
rect 610400 221280 610406 221332
rect 192294 221212 192300 221264
rect 192352 221252 192358 221264
rect 193030 221252 193036 221264
rect 192352 221224 193036 221252
rect 192352 221212 192358 221224
rect 193030 221212 193036 221224
rect 193088 221212 193094 221264
rect 230106 221252 230112 221264
rect 193232 221224 230112 221252
rect 149422 221144 149428 221196
rect 149480 221184 149486 221196
rect 189718 221184 189724 221196
rect 149480 221156 189724 221184
rect 149480 221144 149486 221156
rect 189718 221144 189724 221156
rect 189776 221144 189782 221196
rect 189810 221144 189816 221196
rect 189868 221184 189874 221196
rect 193232 221184 193260 221224
rect 230106 221212 230112 221224
rect 230164 221212 230170 221264
rect 230198 221212 230204 221264
rect 230256 221252 230262 221264
rect 239214 221252 239220 221264
rect 230256 221224 239220 221252
rect 230256 221212 230262 221224
rect 239214 221212 239220 221224
rect 239272 221212 239278 221264
rect 277302 221212 277308 221264
rect 277360 221252 277366 221264
rect 286686 221252 286692 221264
rect 277360 221224 286692 221252
rect 277360 221212 277366 221224
rect 286686 221212 286692 221224
rect 286744 221212 286750 221264
rect 315574 221212 315580 221264
rect 315632 221252 315638 221264
rect 341426 221252 341432 221264
rect 315632 221224 341432 221252
rect 315632 221212 315638 221224
rect 341426 221212 341432 221224
rect 341484 221212 341490 221264
rect 342162 221212 342168 221264
rect 342220 221252 342226 221264
rect 342220 221224 346808 221252
rect 342220 221212 342226 221224
rect 189868 221156 193260 221184
rect 189868 221144 189874 221156
rect 199930 221144 199936 221196
rect 199988 221184 199994 221196
rect 234522 221184 234528 221196
rect 199988 221156 234528 221184
rect 199988 221144 199994 221156
rect 234522 221144 234528 221156
rect 234580 221144 234586 221196
rect 246114 221144 246120 221196
rect 246172 221184 246178 221196
rect 257798 221184 257804 221196
rect 246172 221156 257804 221184
rect 246172 221144 246178 221156
rect 257798 221144 257804 221156
rect 257856 221144 257862 221196
rect 279786 221144 279792 221196
rect 279844 221184 279850 221196
rect 288894 221184 288900 221196
rect 279844 221156 288900 221184
rect 279844 221144 279850 221156
rect 288894 221144 288900 221156
rect 288952 221144 288958 221196
rect 312354 221144 312360 221196
rect 312412 221184 312418 221196
rect 337194 221184 337200 221196
rect 312412 221156 337200 221184
rect 312412 221144 312418 221156
rect 337194 221144 337200 221156
rect 337252 221144 337258 221196
rect 337286 221144 337292 221196
rect 337344 221184 337350 221196
rect 346670 221184 346676 221196
rect 337344 221156 346676 221184
rect 337344 221144 337350 221156
rect 346670 221144 346676 221156
rect 346728 221144 346734 221196
rect 346780 221184 346808 221224
rect 347866 221212 347872 221264
rect 347924 221252 347930 221264
rect 380066 221252 380072 221264
rect 347924 221224 380072 221252
rect 347924 221212 347930 221224
rect 380066 221212 380072 221224
rect 380124 221212 380130 221264
rect 383746 221212 383752 221264
rect 383804 221252 383810 221264
rect 386782 221252 386788 221264
rect 383804 221224 386788 221252
rect 383804 221212 383810 221224
rect 386782 221212 386788 221224
rect 386840 221212 386846 221264
rect 388990 221212 388996 221264
rect 389048 221252 389054 221264
rect 392670 221252 392676 221264
rect 389048 221224 392676 221252
rect 389048 221212 389054 221224
rect 392670 221212 392676 221224
rect 392728 221212 392734 221264
rect 402146 221212 402152 221264
rect 402204 221252 402210 221264
rect 403618 221252 403624 221264
rect 402204 221224 403624 221252
rect 402204 221212 402210 221224
rect 403618 221212 403624 221224
rect 403676 221212 403682 221264
rect 476850 221252 476856 221264
rect 410444 221224 476856 221252
rect 353294 221184 353300 221196
rect 346780 221156 353300 221184
rect 353294 221144 353300 221156
rect 353352 221144 353358 221196
rect 369578 221144 369584 221196
rect 369636 221184 369642 221196
rect 410334 221184 410340 221196
rect 369636 221156 410340 221184
rect 369636 221144 369642 221156
rect 410334 221144 410340 221156
rect 410392 221144 410398 221196
rect 179690 221076 179696 221128
rect 179748 221116 179754 221128
rect 217962 221116 217968 221128
rect 179748 221088 217968 221116
rect 179748 221076 179754 221088
rect 217962 221076 217968 221088
rect 218020 221076 218026 221128
rect 237282 221116 237288 221128
rect 226306 221088 237288 221116
rect 206646 221008 206652 221060
rect 206704 221048 206710 221060
rect 226306 221048 226334 221088
rect 237282 221076 237288 221088
rect 237340 221076 237346 221128
rect 252922 221076 252928 221128
rect 252980 221116 252986 221128
rect 257246 221116 257252 221128
rect 252980 221088 257252 221116
rect 252980 221076 252986 221088
rect 257246 221076 257252 221088
rect 257304 221076 257310 221128
rect 265526 221076 265532 221128
rect 265584 221116 265590 221128
rect 282086 221116 282092 221128
rect 265584 221088 282092 221116
rect 265584 221076 265590 221088
rect 282086 221076 282092 221088
rect 282144 221076 282150 221128
rect 282362 221076 282368 221128
rect 282420 221116 282426 221128
rect 287146 221116 287152 221128
rect 282420 221088 287152 221116
rect 282420 221076 282426 221088
rect 287146 221076 287152 221088
rect 287204 221076 287210 221128
rect 288250 221076 288256 221128
rect 288308 221116 288314 221128
rect 292758 221116 292764 221128
rect 288308 221088 292764 221116
rect 288308 221076 288314 221088
rect 292758 221076 292764 221088
rect 292816 221076 292822 221128
rect 329834 221076 329840 221128
rect 329892 221116 329898 221128
rect 343726 221116 343732 221128
rect 329892 221088 343732 221116
rect 329892 221076 329898 221088
rect 343726 221076 343732 221088
rect 343784 221076 343790 221128
rect 368106 221076 368112 221128
rect 368164 221116 368170 221128
rect 407022 221116 407028 221128
rect 368164 221088 407028 221116
rect 368164 221076 368170 221088
rect 407022 221076 407028 221088
rect 407080 221076 407086 221128
rect 206704 221020 226334 221048
rect 206704 221008 206710 221020
rect 226794 221008 226800 221060
rect 226852 221048 226858 221060
rect 239950 221048 239956 221060
rect 226852 221020 239956 221048
rect 226852 221008 226858 221020
rect 239950 221008 239956 221020
rect 240008 221008 240014 221060
rect 278130 221008 278136 221060
rect 278188 221048 278194 221060
rect 287054 221048 287060 221060
rect 278188 221020 287060 221048
rect 278188 221008 278194 221020
rect 287054 221008 287060 221020
rect 287112 221008 287118 221060
rect 287330 221008 287336 221060
rect 287388 221048 287394 221060
rect 291010 221048 291016 221060
rect 287388 221020 291016 221048
rect 287388 221008 287394 221020
rect 291010 221008 291016 221020
rect 291068 221008 291074 221060
rect 329190 221008 329196 221060
rect 329248 221048 329254 221060
rect 343542 221048 343548 221060
rect 329248 221020 343548 221048
rect 329248 221008 329254 221020
rect 343542 221008 343548 221020
rect 343600 221008 343606 221060
rect 409506 221048 409512 221060
rect 394712 221020 409512 221048
rect 196526 220940 196532 220992
rect 196584 220980 196590 220992
rect 204254 220980 204260 220992
rect 196584 220952 204260 220980
rect 196584 220940 196590 220952
rect 204254 220940 204260 220952
rect 204312 220940 204318 220992
rect 213362 220940 213368 220992
rect 213420 220980 213426 220992
rect 237098 220980 237104 220992
rect 213420 220952 237104 220980
rect 213420 220940 213426 220952
rect 237098 220940 237104 220952
rect 237156 220940 237162 220992
rect 268010 220940 268016 220992
rect 268068 220980 268074 220992
rect 284202 220980 284208 220992
rect 268068 220952 284208 220980
rect 268068 220940 268074 220952
rect 284202 220940 284208 220952
rect 284260 220940 284266 220992
rect 285674 220940 285680 220992
rect 285732 220980 285738 220992
rect 290642 220980 290648 220992
rect 285732 220952 290648 220980
rect 285732 220940 285738 220952
rect 290642 220940 290648 220952
rect 290700 220940 290706 220992
rect 291562 220940 291568 220992
rect 291620 220980 291626 220992
rect 294230 220980 294236 220992
rect 291620 220952 294236 220980
rect 291620 220940 291626 220952
rect 294230 220940 294236 220952
rect 294288 220940 294294 220992
rect 334158 220940 334164 220992
rect 334216 220980 334222 220992
rect 349890 220980 349896 220992
rect 334216 220952 349896 220980
rect 334216 220940 334222 220952
rect 349890 220940 349896 220952
rect 349948 220940 349954 220992
rect 381170 220940 381176 220992
rect 381228 220980 381234 220992
rect 394712 220980 394740 221020
rect 409506 221008 409512 221020
rect 409564 221008 409570 221060
rect 381228 220952 394740 220980
rect 381228 220940 381234 220952
rect 394786 220940 394792 220992
rect 394844 220980 394850 220992
rect 401134 220980 401140 220992
rect 394844 220952 401140 220980
rect 394844 220940 394850 220952
rect 401134 220940 401140 220952
rect 401192 220940 401198 220992
rect 162026 220872 162032 220924
rect 162084 220912 162090 220924
rect 238938 220912 238944 220924
rect 162084 220884 238944 220912
rect 162084 220872 162090 220884
rect 238938 220872 238944 220884
rect 238996 220872 239002 220924
rect 276474 220872 276480 220924
rect 276532 220912 276538 220924
rect 287422 220912 287428 220924
rect 276532 220884 287428 220912
rect 276532 220872 276538 220884
rect 287422 220872 287428 220884
rect 287480 220872 287486 220924
rect 369670 220872 369676 220924
rect 369728 220912 369734 220924
rect 382642 220912 382648 220924
rect 369728 220884 382648 220912
rect 369728 220872 369734 220884
rect 382642 220872 382648 220884
rect 382700 220872 382706 220924
rect 391842 220872 391848 220924
rect 391900 220912 391906 220924
rect 399478 220912 399484 220924
rect 391900 220884 399484 220912
rect 391900 220872 391906 220884
rect 399478 220872 399484 220884
rect 399536 220872 399542 220924
rect 400490 220872 400496 220924
rect 400548 220912 400554 220924
rect 410444 220912 410472 221224
rect 476850 221212 476856 221224
rect 476908 221212 476914 221264
rect 527542 221212 527548 221264
rect 527600 221252 527606 221264
rect 628006 221252 628012 221264
rect 527600 221224 628012 221252
rect 527600 221212 527606 221224
rect 628006 221212 628012 221224
rect 628064 221212 628070 221264
rect 411898 221144 411904 221196
rect 411956 221184 411962 221196
rect 485222 221184 485228 221196
rect 411956 221156 485228 221184
rect 411956 221144 411962 221156
rect 485222 221144 485228 221156
rect 485280 221144 485286 221196
rect 505738 221144 505744 221196
rect 505796 221184 505802 221196
rect 609422 221184 609428 221196
rect 505796 221156 609428 221184
rect 505796 221144 505802 221156
rect 609422 221144 609428 221156
rect 609480 221144 609486 221196
rect 670050 221144 670056 221196
rect 670108 221184 670114 221196
rect 675938 221184 675944 221196
rect 670108 221156 675944 221184
rect 670108 221144 670114 221156
rect 675938 221144 675944 221156
rect 675996 221144 676002 221196
rect 503530 221076 503536 221128
rect 503588 221116 503594 221128
rect 608962 221116 608968 221128
rect 503588 221088 608968 221116
rect 503588 221076 503594 221088
rect 608962 221076 608968 221088
rect 609020 221076 609026 221128
rect 517238 221008 517244 221060
rect 517296 221048 517302 221060
rect 517882 221048 517888 221060
rect 517296 221020 517888 221048
rect 517296 221008 517302 221020
rect 517882 221008 517888 221020
rect 517940 221048 517946 221060
rect 626166 221048 626172 221060
rect 517940 221020 626172 221048
rect 517940 221008 517946 221020
rect 626166 221008 626172 221020
rect 626224 221008 626230 221060
rect 669038 221008 669044 221060
rect 669096 221048 669102 221060
rect 676030 221048 676036 221060
rect 669096 221020 676036 221048
rect 669096 221008 669102 221020
rect 676030 221008 676036 221020
rect 676088 221008 676094 221060
rect 500678 220940 500684 220992
rect 500736 220980 500742 220992
rect 608502 220980 608508 220992
rect 500736 220952 608508 220980
rect 500736 220940 500742 220952
rect 608502 220940 608508 220952
rect 608560 220940 608566 220992
rect 400548 220884 410472 220912
rect 400548 220872 400554 220884
rect 499022 220872 499028 220924
rect 499080 220912 499086 220924
rect 608042 220912 608048 220924
rect 499080 220884 608048 220912
rect 499080 220872 499086 220884
rect 608042 220872 608048 220884
rect 608100 220872 608106 220924
rect 194042 220804 194048 220856
rect 194100 220844 194106 220856
rect 252830 220844 252836 220856
rect 194100 220816 252836 220844
rect 194100 220804 194106 220816
rect 252830 220804 252836 220816
rect 252888 220804 252894 220856
rect 385402 220804 385408 220856
rect 385460 220844 385466 220856
rect 507946 220844 507952 220856
rect 385460 220816 507952 220844
rect 385460 220804 385466 220816
rect 507946 220804 507952 220816
rect 508004 220804 508010 220856
rect 548334 220804 548340 220856
rect 548392 220844 548398 220856
rect 617334 220844 617340 220856
rect 548392 220816 617340 220844
rect 548392 220804 548398 220816
rect 617334 220804 617340 220816
rect 617392 220804 617398 220856
rect 666462 220804 666468 220856
rect 666520 220844 666526 220856
rect 675662 220844 675668 220856
rect 666520 220816 675668 220844
rect 666520 220804 666526 220816
rect 675662 220804 675668 220816
rect 675720 220804 675726 220856
rect 347682 220736 347688 220788
rect 347740 220776 347746 220788
rect 419718 220776 419724 220788
rect 347740 220748 419724 220776
rect 347740 220736 347746 220748
rect 419718 220736 419724 220748
rect 419776 220736 419782 220788
rect 571702 220736 571708 220788
rect 571760 220776 571766 220788
rect 572714 220776 572720 220788
rect 571760 220748 572720 220776
rect 571760 220736 571766 220748
rect 572714 220736 572720 220748
rect 572772 220736 572778 220788
rect 574094 220736 574100 220788
rect 574152 220776 574158 220788
rect 575198 220776 575204 220788
rect 574152 220748 575204 220776
rect 574152 220736 574158 220748
rect 575198 220736 575204 220748
rect 575256 220736 575262 220788
rect 351270 220668 351276 220720
rect 351328 220708 351334 220720
rect 425514 220708 425520 220720
rect 351328 220680 425520 220708
rect 351328 220668 351334 220680
rect 425514 220668 425520 220680
rect 425572 220668 425578 220720
rect 571610 220668 571616 220720
rect 571668 220708 571674 220720
rect 573542 220708 573548 220720
rect 571668 220680 573548 220708
rect 571668 220668 571674 220680
rect 573542 220668 573548 220680
rect 573600 220668 573606 220720
rect 352006 220600 352012 220652
rect 352064 220640 352070 220652
rect 429746 220640 429752 220652
rect 352064 220612 429752 220640
rect 352064 220600 352070 220612
rect 429746 220600 429752 220612
rect 429804 220600 429810 220652
rect 353386 220532 353392 220584
rect 353444 220572 353450 220584
rect 433334 220572 433340 220584
rect 353444 220544 433340 220572
rect 353444 220532 353450 220544
rect 433334 220532 433340 220544
rect 433392 220532 433398 220584
rect 356238 220464 356244 220516
rect 356296 220504 356302 220516
rect 439774 220504 439780 220516
rect 356296 220476 439780 220504
rect 356296 220464 356302 220476
rect 439774 220464 439780 220476
rect 439832 220464 439838 220516
rect 355042 220396 355048 220448
rect 355100 220436 355106 220448
rect 436462 220436 436468 220448
rect 355100 220408 436468 220436
rect 355100 220396 355106 220408
rect 436462 220396 436468 220408
rect 436520 220396 436526 220448
rect 359366 220328 359372 220380
rect 359424 220368 359430 220380
rect 446582 220368 446588 220380
rect 359424 220340 446588 220368
rect 359424 220328 359430 220340
rect 446582 220328 446588 220340
rect 446640 220328 446646 220380
rect 139302 220260 139308 220312
rect 139360 220300 139366 220312
rect 228266 220300 228272 220312
rect 139360 220272 228272 220300
rect 139360 220260 139366 220272
rect 228266 220260 228272 220272
rect 228324 220260 228330 220312
rect 357710 220260 357716 220312
rect 357768 220300 357774 220312
rect 443178 220300 443184 220312
rect 357768 220272 443184 220300
rect 357768 220260 357774 220272
rect 443178 220260 443184 220272
rect 443236 220260 443242 220312
rect 142706 220192 142712 220244
rect 142764 220232 142770 220244
rect 229646 220232 229652 220244
rect 142764 220204 229652 220232
rect 142764 220192 142770 220204
rect 229646 220192 229652 220204
rect 229704 220192 229710 220244
rect 361942 220192 361948 220244
rect 362000 220232 362006 220244
rect 453298 220232 453304 220244
rect 362000 220204 453304 220232
rect 362000 220192 362006 220204
rect 453298 220192 453304 220204
rect 453356 220192 453362 220244
rect 135990 220124 135996 220176
rect 136048 220164 136054 220176
rect 226610 220164 226616 220176
rect 136048 220136 226616 220164
rect 136048 220124 136054 220136
rect 226610 220124 226616 220136
rect 226668 220124 226674 220176
rect 360562 220124 360568 220176
rect 360620 220164 360626 220176
rect 449894 220164 449900 220176
rect 360620 220136 449900 220164
rect 360620 220124 360626 220136
rect 449894 220124 449900 220136
rect 449952 220124 449958 220176
rect 132402 220056 132408 220108
rect 132460 220096 132466 220108
rect 225414 220096 225420 220108
rect 132460 220068 225420 220096
rect 132460 220056 132466 220068
rect 225414 220056 225420 220068
rect 225472 220056 225478 220108
rect 364794 220056 364800 220108
rect 364852 220096 364858 220108
rect 460014 220096 460020 220108
rect 364852 220068 460020 220096
rect 364852 220056 364858 220068
rect 460014 220056 460020 220068
rect 460072 220056 460078 220108
rect 129274 219988 129280 220040
rect 129332 220028 129338 220040
rect 223942 220028 223948 220040
rect 129332 220000 223948 220028
rect 129332 219988 129338 220000
rect 223942 219988 223948 220000
rect 224000 219988 224006 220040
rect 363414 219988 363420 220040
rect 363472 220028 363478 220040
rect 456610 220028 456616 220040
rect 363472 220000 456616 220028
rect 363472 219988 363478 220000
rect 456610 219988 456616 220000
rect 456668 219988 456674 220040
rect 125870 219920 125876 219972
rect 125928 219960 125934 219972
rect 222286 219960 222292 219972
rect 125928 219932 222292 219960
rect 125928 219920 125934 219932
rect 222286 219920 222292 219932
rect 222344 219920 222350 219972
rect 367646 219920 367652 219972
rect 367704 219960 367710 219972
rect 466730 219960 466736 219972
rect 367704 219932 466736 219960
rect 367704 219920 367710 219932
rect 466730 219920 466736 219932
rect 466788 219920 466794 219972
rect 122466 219852 122472 219904
rect 122524 219892 122530 219904
rect 221090 219892 221096 219904
rect 122524 219864 221096 219892
rect 122524 219852 122530 219864
rect 221090 219852 221096 219864
rect 221148 219852 221154 219904
rect 366266 219852 366272 219904
rect 366324 219892 366330 219904
rect 463694 219892 463700 219904
rect 366324 219864 463700 219892
rect 366324 219852 366330 219864
rect 463694 219852 463700 219864
rect 463752 219852 463758 219904
rect 58618 219784 58624 219836
rect 58676 219824 58682 219836
rect 193766 219824 193772 219836
rect 58676 219796 193772 219824
rect 58676 219784 58682 219796
rect 193766 219784 193772 219796
rect 193824 219784 193830 219836
rect 369302 219784 369308 219836
rect 369360 219824 369366 219836
rect 470134 219824 470140 219836
rect 369360 219796 470140 219824
rect 369360 219784 369366 219796
rect 470134 219784 470140 219796
rect 470192 219784 470198 219836
rect 48498 219716 48504 219768
rect 48556 219756 48562 219768
rect 648522 219756 648528 219768
rect 48556 219728 648528 219756
rect 48556 219716 48562 219728
rect 648522 219716 648528 219728
rect 648580 219716 648586 219768
rect 46014 219648 46020 219700
rect 46072 219688 46078 219700
rect 647142 219688 647148 219700
rect 46072 219660 647148 219688
rect 46072 219648 46078 219660
rect 647142 219648 647148 219660
rect 647200 219648 647206 219700
rect 48590 219580 48596 219632
rect 48648 219620 48654 219632
rect 651282 219620 651288 219632
rect 48648 219592 651288 219620
rect 48648 219580 48654 219592
rect 651282 219580 651288 219592
rect 651340 219580 651346 219632
rect 652754 219580 652760 219632
rect 652812 219580 652818 219632
rect 46290 219512 46296 219564
rect 46348 219552 46354 219564
rect 649902 219552 649908 219564
rect 46348 219524 649908 219552
rect 46348 219512 46354 219524
rect 649902 219512 649908 219524
rect 649960 219512 649966 219564
rect 652772 219552 652800 219580
rect 675570 219552 675576 219564
rect 652772 219524 675576 219552
rect 675570 219512 675576 219524
rect 675628 219552 675634 219564
rect 676030 219552 676036 219564
rect 675628 219524 676036 219552
rect 675628 219512 675634 219524
rect 676030 219512 676036 219524
rect 676088 219512 676094 219564
rect 48682 219444 48688 219496
rect 48740 219484 48746 219496
rect 652754 219484 652760 219496
rect 48740 219456 652760 219484
rect 48740 219444 48746 219456
rect 652754 219444 652760 219456
rect 652812 219444 652818 219496
rect 48774 219376 48780 219428
rect 48832 219416 48838 219428
rect 654134 219416 654140 219428
rect 48832 219388 654140 219416
rect 48832 219376 48838 219388
rect 654134 219376 654140 219388
rect 654192 219376 654198 219428
rect 349154 219308 349160 219360
rect 349212 219348 349218 219360
rect 423030 219348 423036 219360
rect 349212 219320 423036 219348
rect 349212 219308 349218 219320
rect 423030 219308 423036 219320
rect 423088 219308 423094 219360
rect 652662 219308 652668 219360
rect 652720 219348 652726 219360
rect 674834 219348 674840 219360
rect 652720 219320 674840 219348
rect 652720 219308 652726 219320
rect 674834 219308 674840 219320
rect 674892 219348 674898 219360
rect 676030 219348 676036 219360
rect 674892 219320 676036 219348
rect 674892 219308 674898 219320
rect 676030 219308 676036 219320
rect 676088 219308 676094 219360
rect 350534 219240 350540 219292
rect 350592 219280 350598 219292
rect 426342 219280 426348 219292
rect 350592 219252 426348 219280
rect 350592 219240 350598 219252
rect 426342 219240 426348 219252
rect 426400 219240 426406 219292
rect 344830 219172 344836 219224
rect 344888 219212 344894 219224
rect 412910 219212 412916 219224
rect 344888 219184 412916 219212
rect 344888 219172 344894 219184
rect 412910 219172 412916 219184
rect 412968 219172 412974 219224
rect 346302 219104 346308 219156
rect 346360 219144 346366 219156
rect 416222 219144 416228 219156
rect 346360 219116 416228 219144
rect 346360 219104 346366 219116
rect 416222 219104 416228 219116
rect 416280 219104 416286 219156
rect 523402 218492 523408 218544
rect 523460 218532 523466 218544
rect 612642 218532 612648 218544
rect 523460 218504 612648 218532
rect 523460 218492 523466 218504
rect 612642 218492 612648 218504
rect 612700 218492 612706 218544
rect 525794 218424 525800 218476
rect 525852 218464 525858 218476
rect 613102 218464 613108 218476
rect 525852 218436 613108 218464
rect 525852 218424 525858 218436
rect 613102 218424 613108 218436
rect 613160 218424 613166 218476
rect 520826 218356 520832 218408
rect 520884 218396 520890 218408
rect 612182 218396 612188 218408
rect 520884 218368 612188 218396
rect 520884 218356 520890 218368
rect 612182 218356 612188 218368
rect 612240 218356 612246 218408
rect 518710 218288 518716 218340
rect 518768 218328 518774 218340
rect 611722 218328 611728 218340
rect 518768 218300 611728 218328
rect 518768 218288 518774 218300
rect 611722 218288 611728 218300
rect 611780 218288 611786 218340
rect 674098 218288 674104 218340
rect 674156 218328 674162 218340
rect 676030 218328 676036 218340
rect 674156 218300 676036 218328
rect 674156 218288 674162 218300
rect 676030 218288 676036 218300
rect 676088 218288 676094 218340
rect 513466 218220 513472 218272
rect 513524 218260 513530 218272
rect 515766 218260 515772 218272
rect 513524 218232 515772 218260
rect 513524 218220 513530 218232
rect 515766 218220 515772 218232
rect 515824 218260 515830 218272
rect 611262 218260 611268 218272
rect 515824 218232 611268 218260
rect 515824 218220 515830 218232
rect 611262 218220 611268 218232
rect 611320 218220 611326 218272
rect 662598 218220 662604 218272
rect 662656 218260 662662 218272
rect 663978 218260 663984 218272
rect 662656 218232 663984 218260
rect 662656 218220 662662 218232
rect 663978 218220 663984 218232
rect 664036 218220 664042 218272
rect 490282 218152 490288 218204
rect 490340 218192 490346 218204
rect 607122 218192 607128 218204
rect 490340 218164 607128 218192
rect 490340 218152 490346 218164
rect 607122 218152 607128 218164
rect 607180 218152 607186 218204
rect 487154 218084 487160 218136
rect 487212 218124 487218 218136
rect 606662 218124 606668 218136
rect 487212 218096 606668 218124
rect 487212 218084 487218 218096
rect 606662 218084 606668 218096
rect 606720 218084 606726 218136
rect 662598 218084 662604 218136
rect 662656 218124 662662 218136
rect 662874 218124 662880 218136
rect 662656 218096 662880 218124
rect 662656 218084 662662 218096
rect 662874 218084 662880 218096
rect 662932 218084 662938 218136
rect 673454 218084 673460 218136
rect 673512 218124 673518 218136
rect 675938 218124 675944 218136
rect 673512 218096 675944 218124
rect 673512 218084 673518 218096
rect 675938 218084 675944 218096
rect 675996 218084 676002 218136
rect 46934 218016 46940 218068
rect 46992 218056 46998 218068
rect 671154 218056 671160 218068
rect 46992 218028 671160 218056
rect 46992 218016 46998 218028
rect 671154 218016 671160 218028
rect 671212 218016 671218 218068
rect 674374 218016 674380 218068
rect 674432 218056 674438 218068
rect 676030 218056 676036 218068
rect 674432 218028 676036 218056
rect 674432 218016 674438 218028
rect 676030 218016 676036 218028
rect 676088 218016 676094 218068
rect 418154 217948 418160 218000
rect 418212 217988 418218 218000
rect 418614 217988 418620 218000
rect 418212 217960 418620 217988
rect 418212 217948 418218 217960
rect 418614 217948 418620 217960
rect 418672 217948 418678 218000
rect 646958 217948 646964 218000
rect 647016 217988 647022 218000
rect 651650 217988 651656 218000
rect 647016 217960 651656 217988
rect 647016 217948 647022 217960
rect 651650 217948 651656 217960
rect 651708 217948 651714 218000
rect 642726 217880 642732 217932
rect 642784 217920 642790 217932
rect 651374 217920 651380 217932
rect 642784 217892 651380 217920
rect 642784 217880 642790 217892
rect 651374 217880 651380 217892
rect 651432 217880 651438 217932
rect 662506 217880 662512 217932
rect 662564 217920 662570 217932
rect 664438 217920 664444 217932
rect 662564 217892 664444 217920
rect 662564 217880 662570 217892
rect 664438 217880 664444 217892
rect 664496 217880 664502 217932
rect 644106 217812 644112 217864
rect 644164 217852 644170 217864
rect 651466 217852 651472 217864
rect 644164 217824 651472 217852
rect 644164 217812 644170 217824
rect 651466 217812 651472 217824
rect 651524 217812 651530 217864
rect 570690 217404 570696 217456
rect 570748 217444 570754 217456
rect 635918 217444 635924 217456
rect 570748 217416 635924 217444
rect 570748 217404 570754 217416
rect 635918 217404 635924 217416
rect 635976 217404 635982 217456
rect 563054 217336 563060 217388
rect 563112 217376 563118 217388
rect 634538 217376 634544 217388
rect 563112 217348 634544 217376
rect 563112 217336 563118 217348
rect 634538 217336 634544 217348
rect 634596 217336 634602 217388
rect 558178 217268 558184 217320
rect 558236 217308 558242 217320
rect 633618 217308 633624 217320
rect 558236 217280 633624 217308
rect 558236 217268 558242 217280
rect 633618 217268 633624 217280
rect 633676 217268 633682 217320
rect 550634 217200 550640 217252
rect 550692 217240 550698 217252
rect 632238 217240 632244 217252
rect 550692 217212 632244 217240
rect 550692 217200 550698 217212
rect 632238 217200 632244 217212
rect 632296 217200 632302 217252
rect 540514 217132 540520 217184
rect 540572 217172 540578 217184
rect 630398 217172 630404 217184
rect 540572 217144 630404 217172
rect 540572 217132 540578 217144
rect 630398 217132 630404 217144
rect 630456 217132 630462 217184
rect 535362 217064 535368 217116
rect 535420 217104 535426 217116
rect 629478 217104 629484 217116
rect 535420 217076 629484 217104
rect 535420 217064 535426 217076
rect 629478 217064 629484 217076
rect 629536 217064 629542 217116
rect 673638 217064 673644 217116
rect 673696 217104 673702 217116
rect 675938 217104 675944 217116
rect 673696 217076 675944 217104
rect 673696 217064 673702 217076
rect 675938 217064 675944 217076
rect 675996 217064 676002 217116
rect 530302 216996 530308 217048
rect 530360 217036 530366 217048
rect 628466 217036 628472 217048
rect 530360 217008 628472 217036
rect 530360 216996 530366 217008
rect 628466 216996 628472 217008
rect 628524 216996 628530 217048
rect 513466 216928 513472 216980
rect 513524 216968 513530 216980
rect 610802 216968 610808 216980
rect 513524 216940 610808 216968
rect 513524 216928 513530 216940
rect 610802 216928 610808 216940
rect 610860 216928 610866 216980
rect 525426 216860 525432 216912
rect 525484 216900 525490 216912
rect 627546 216900 627552 216912
rect 525484 216872 627552 216900
rect 525484 216860 525490 216872
rect 627546 216860 627552 216872
rect 627604 216860 627610 216912
rect 418522 216792 418528 216844
rect 418580 216832 418586 216844
rect 639690 216832 639696 216844
rect 418580 216804 639696 216832
rect 418580 216792 418586 216804
rect 639690 216792 639696 216804
rect 639748 216792 639754 216844
rect 41414 216724 41420 216776
rect 41472 216764 41478 216776
rect 59262 216764 59268 216776
rect 41472 216736 59268 216764
rect 41472 216724 41478 216736
rect 59262 216724 59268 216736
rect 59320 216724 59326 216776
rect 418430 216724 418436 216776
rect 418488 216764 418494 216776
rect 640610 216764 640616 216776
rect 418488 216736 640616 216764
rect 418488 216724 418494 216736
rect 640610 216724 640616 216736
rect 640668 216724 640674 216776
rect 41598 216656 41604 216708
rect 41656 216696 41662 216708
rect 59446 216696 59452 216708
rect 41656 216668 59452 216696
rect 41656 216656 41662 216668
rect 59446 216656 59452 216668
rect 59504 216656 59510 216708
rect 418614 216656 418620 216708
rect 418672 216696 418678 216708
rect 640150 216696 640156 216708
rect 418672 216668 640156 216696
rect 418672 216656 418678 216668
rect 640150 216656 640156 216668
rect 640208 216656 640214 216708
rect 645578 216656 645584 216708
rect 645636 216696 645642 216708
rect 651558 216696 651564 216708
rect 645636 216668 651564 216696
rect 645636 216656 645642 216668
rect 651558 216656 651564 216668
rect 651616 216656 651622 216708
rect 674190 216656 674196 216708
rect 674248 216696 674254 216708
rect 676030 216696 676036 216708
rect 674248 216668 676036 216696
rect 674248 216656 674254 216668
rect 676030 216656 676036 216668
rect 676088 216656 676094 216708
rect 41506 216588 41512 216640
rect 41564 216628 41570 216640
rect 59354 216628 59360 216640
rect 41564 216600 59360 216628
rect 41564 216588 41570 216600
rect 59354 216588 59360 216600
rect 59412 216588 59418 216640
rect 417878 216588 417884 216640
rect 417936 216628 417942 216640
rect 641070 216628 641076 216640
rect 417936 216600 641076 216628
rect 417936 216588 417942 216600
rect 641070 216588 641076 216600
rect 641128 216588 641134 216640
rect 492490 216520 492496 216572
rect 492548 216560 492554 216572
rect 504450 216560 504456 216572
rect 492548 216532 504456 216560
rect 492548 216520 492554 216532
rect 504450 216520 504456 216532
rect 504508 216520 504514 216572
rect 505002 216520 505008 216572
rect 505060 216560 505066 216572
rect 505060 216532 508544 216560
rect 505060 216520 505066 216532
rect 495986 216452 495992 216504
rect 496044 216492 496050 216504
rect 496044 216464 504864 216492
rect 496044 216452 496050 216464
rect 484210 216384 484216 216436
rect 484268 216424 484274 216436
rect 484268 216396 486096 216424
rect 484268 216384 484274 216396
rect 486068 215948 486096 216396
rect 486694 216384 486700 216436
rect 486752 216424 486758 216436
rect 486752 216396 488534 216424
rect 486752 216384 486758 216396
rect 488506 216016 488534 216396
rect 490098 216384 490104 216436
rect 490156 216424 490162 216436
rect 490156 216396 495710 216424
rect 490156 216384 490162 216396
rect 495682 216084 495710 216396
rect 500218 216384 500224 216436
rect 500276 216424 500282 216436
rect 500276 216396 502472 216424
rect 500276 216384 500282 216396
rect 502444 216152 502472 216396
rect 504450 216384 504456 216436
rect 504508 216384 504514 216436
rect 504836 216424 504864 216464
rect 504836 216396 505140 216424
rect 504468 216220 504496 216384
rect 505112 216288 505140 216396
rect 508516 216356 508544 216532
rect 520366 216520 520372 216572
rect 520424 216560 520430 216572
rect 626626 216560 626632 216572
rect 520424 216532 626632 216560
rect 520424 216520 520430 216532
rect 626626 216520 626632 216532
rect 626684 216520 626690 216572
rect 515214 216452 515220 216504
rect 515272 216492 515278 216504
rect 625706 216492 625712 216504
rect 515272 216464 625712 216492
rect 515272 216452 515278 216464
rect 625706 216452 625712 216464
rect 625764 216452 625770 216504
rect 510246 216384 510252 216436
rect 510304 216424 510310 216436
rect 624786 216424 624792 216436
rect 510304 216396 624792 216424
rect 510304 216384 510310 216396
rect 624786 216384 624792 216396
rect 624844 216384 624850 216436
rect 623866 216356 623872 216368
rect 508516 216328 623872 216356
rect 623866 216316 623872 216328
rect 623924 216316 623930 216368
rect 622486 216288 622492 216300
rect 505112 216260 622492 216288
rect 622486 216248 622492 216260
rect 622544 216248 622550 216300
rect 673546 216248 673552 216300
rect 673604 216288 673610 216300
rect 675938 216288 675944 216300
rect 673604 216260 675944 216288
rect 673604 216248 673610 216260
rect 675938 216248 675944 216260
rect 675996 216248 676002 216300
rect 622026 216220 622032 216232
rect 504468 216192 622032 216220
rect 622026 216180 622032 216192
rect 622084 216180 622090 216232
rect 637850 216152 637856 216164
rect 502444 216124 637856 216152
rect 637850 216112 637856 216124
rect 637908 216112 637914 216164
rect 636378 216084 636384 216096
rect 495682 216056 636384 216084
rect 636378 216044 636384 216056
rect 636436 216044 636442 216096
rect 638310 216016 638316 216028
rect 488506 215988 638316 216016
rect 638310 215976 638316 215988
rect 638368 215976 638374 216028
rect 638770 215948 638776 215960
rect 486068 215920 638776 215948
rect 638770 215908 638776 215920
rect 638828 215908 638834 215960
rect 48222 215840 48228 215892
rect 48280 215880 48286 215892
rect 666186 215880 666192 215892
rect 48280 215852 666192 215880
rect 48280 215840 48286 215852
rect 666186 215840 666192 215852
rect 666244 215840 666250 215892
rect 31662 215772 31668 215824
rect 31720 215812 31726 215824
rect 665266 215812 665272 215824
rect 31720 215784 665272 215812
rect 31720 215772 31726 215784
rect 665266 215772 665272 215784
rect 665324 215772 665330 215824
rect 29178 215704 29184 215756
rect 29236 215744 29242 215756
rect 665726 215744 665732 215756
rect 29236 215716 665732 215744
rect 29236 215704 29242 215716
rect 665726 215704 665732 215716
rect 665784 215704 665790 215756
rect 580166 215568 580172 215620
rect 580224 215608 580230 215620
rect 599762 215608 599768 215620
rect 580224 215580 599768 215608
rect 580224 215568 580230 215580
rect 599762 215568 599768 215580
rect 599820 215568 599826 215620
rect 673914 215432 673920 215484
rect 673972 215472 673978 215484
rect 675846 215472 675852 215484
rect 673972 215444 675852 215472
rect 673972 215432 673978 215444
rect 675846 215432 675852 215444
rect 675904 215432 675910 215484
rect 674282 215364 674288 215416
rect 674340 215404 674346 215416
rect 675938 215404 675944 215416
rect 674340 215376 675944 215404
rect 674340 215364 674346 215376
rect 675938 215364 675944 215376
rect 675996 215364 676002 215416
rect 674466 215296 674472 215348
rect 674524 215336 674530 215348
rect 676030 215336 676036 215348
rect 674524 215308 676036 215336
rect 674524 215296 674530 215308
rect 676030 215296 676036 215308
rect 676088 215296 676094 215348
rect 656894 215092 656900 215144
rect 656952 215132 656958 215144
rect 657906 215132 657912 215144
rect 656952 215104 657912 215132
rect 656952 215092 656958 215104
rect 657906 215092 657912 215104
rect 657964 215092 657970 215144
rect 659654 215092 659660 215144
rect 659712 215132 659718 215144
rect 660758 215132 660764 215144
rect 659712 215104 660764 215132
rect 659712 215092 659718 215104
rect 660758 215092 660764 215104
rect 660816 215092 660822 215144
rect 673822 214616 673828 214668
rect 673880 214656 673886 214668
rect 676030 214656 676036 214668
rect 673880 214628 676036 214656
rect 673880 214616 673886 214628
rect 676030 214616 676036 214628
rect 676088 214616 676094 214668
rect 41506 214208 41512 214260
rect 41564 214248 41570 214260
rect 43438 214248 43444 214260
rect 41564 214220 43444 214248
rect 41564 214208 41570 214220
rect 43438 214208 43444 214220
rect 43496 214208 43502 214260
rect 41414 213868 41420 213920
rect 41472 213908 41478 213920
rect 45554 213908 45560 213920
rect 41472 213880 45560 213908
rect 41472 213868 41478 213880
rect 45554 213868 45560 213880
rect 45612 213868 45618 213920
rect 674006 213800 674012 213852
rect 674064 213840 674070 213852
rect 676030 213840 676036 213852
rect 674064 213812 676036 213840
rect 674064 213800 674070 213812
rect 676030 213800 676036 213812
rect 676088 213800 676094 213852
rect 582282 212576 582288 212628
rect 582340 212616 582346 212628
rect 599946 212616 599952 212628
rect 582340 212588 599952 212616
rect 582340 212576 582346 212588
rect 599946 212576 599952 212588
rect 600004 212576 600010 212628
rect 673730 212576 673736 212628
rect 673788 212616 673794 212628
rect 675938 212616 675944 212628
rect 673788 212588 675944 212616
rect 673788 212576 673794 212588
rect 675938 212576 675944 212588
rect 675996 212576 676002 212628
rect 580258 212508 580264 212560
rect 580316 212548 580322 212560
rect 599854 212548 599860 212560
rect 580316 212520 599860 212548
rect 580316 212508 580322 212520
rect 599854 212508 599860 212520
rect 599912 212508 599918 212560
rect 675202 212508 675208 212560
rect 675260 212548 675266 212560
rect 676030 212548 676036 212560
rect 675260 212520 676036 212548
rect 675260 212508 675266 212520
rect 676030 212508 676036 212520
rect 676088 212508 676094 212560
rect 651282 212440 651288 212492
rect 651340 212480 651346 212492
rect 651374 212480 651380 212492
rect 651340 212452 651380 212480
rect 651340 212440 651346 212452
rect 651374 212440 651380 212452
rect 651432 212440 651438 212492
rect 673178 212032 673184 212084
rect 673236 212072 673242 212084
rect 676030 212072 676036 212084
rect 673236 212044 676036 212072
rect 673236 212032 673242 212044
rect 676030 212032 676036 212044
rect 676088 212032 676094 212084
rect 662414 210876 662420 210928
rect 662472 210916 662478 210928
rect 662690 210916 662696 210928
rect 662472 210888 662696 210916
rect 662472 210876 662478 210888
rect 662690 210876 662696 210888
rect 662748 210876 662754 210928
rect 581638 209856 581644 209908
rect 581696 209896 581702 209908
rect 600038 209896 600044 209908
rect 581696 209868 600044 209896
rect 581696 209856 581702 209868
rect 600038 209856 600044 209868
rect 600096 209856 600102 209908
rect 580534 209788 580540 209840
rect 580592 209828 580598 209840
rect 599118 209828 599124 209840
rect 580592 209800 599124 209828
rect 580592 209788 580598 209800
rect 599118 209788 599124 209800
rect 599176 209788 599182 209840
rect 579706 207068 579712 207120
rect 579764 207108 579770 207120
rect 601510 207108 601516 207120
rect 579764 207080 601516 207108
rect 579764 207068 579770 207080
rect 601510 207068 601516 207080
rect 601568 207068 601574 207120
rect 582282 207000 582288 207052
rect 582340 207040 582346 207052
rect 601418 207040 601424 207052
rect 582340 207012 601424 207040
rect 582340 207000 582346 207012
rect 601418 207000 601424 207012
rect 601476 207000 601482 207052
rect 674558 206116 674564 206168
rect 674616 206156 674622 206168
rect 674834 206156 674840 206168
rect 674616 206128 674840 206156
rect 674616 206116 674622 206128
rect 674834 206116 674840 206128
rect 674892 206116 674898 206168
rect 674834 205980 674840 206032
rect 674892 206020 674898 206032
rect 675386 206020 675392 206032
rect 674892 205992 675392 206020
rect 674892 205980 674898 205992
rect 675386 205980 675392 205992
rect 675444 205980 675450 206032
rect 675754 205980 675760 206032
rect 675812 205980 675818 206032
rect 674650 205708 674656 205760
rect 674708 205748 674714 205760
rect 675202 205748 675208 205760
rect 674708 205720 675208 205748
rect 674708 205708 674714 205720
rect 675202 205708 675208 205720
rect 675260 205708 675266 205760
rect 674374 205504 674380 205556
rect 674432 205544 674438 205556
rect 675294 205544 675300 205556
rect 674432 205516 675300 205544
rect 674432 205504 674438 205516
rect 675294 205504 675300 205516
rect 675352 205504 675358 205556
rect 675772 205476 675800 205980
rect 674392 205448 675800 205476
rect 674392 205420 674420 205448
rect 674374 205368 674380 205420
rect 674432 205368 674438 205420
rect 674466 205164 674472 205216
rect 674524 205204 674530 205216
rect 675294 205204 675300 205216
rect 674524 205176 675300 205204
rect 674524 205164 674530 205176
rect 675294 205164 675300 205176
rect 675352 205164 675358 205216
rect 674098 204552 674104 204604
rect 674156 204592 674162 204604
rect 675294 204592 675300 204604
rect 674156 204564 675300 204592
rect 674156 204552 674162 204564
rect 675294 204552 675300 204564
rect 675352 204552 675358 204604
rect 582282 204280 582288 204332
rect 582340 204320 582346 204332
rect 599946 204320 599952 204332
rect 582340 204292 599952 204320
rect 582340 204280 582346 204292
rect 599946 204280 599952 204292
rect 600004 204280 600010 204332
rect 674190 202716 674196 202768
rect 674248 202756 674254 202768
rect 675478 202756 675484 202768
rect 674248 202728 675484 202756
rect 674248 202716 674254 202728
rect 675478 202716 675484 202728
rect 675536 202716 675542 202768
rect 674282 201832 674288 201884
rect 674340 201872 674346 201884
rect 675386 201872 675392 201884
rect 674340 201844 675392 201872
rect 674340 201832 674346 201844
rect 675386 201832 675392 201844
rect 675444 201832 675450 201884
rect 581086 201560 581092 201612
rect 581144 201600 581150 201612
rect 599946 201600 599952 201612
rect 581144 201572 599952 201600
rect 581144 201560 581150 201572
rect 599946 201560 599952 201572
rect 600004 201560 600010 201612
rect 580718 201492 580724 201544
rect 580776 201532 580782 201544
rect 598934 201532 598940 201544
rect 580776 201504 598940 201532
rect 580776 201492 580782 201504
rect 598934 201492 598940 201504
rect 598992 201492 598998 201544
rect 673914 201492 673920 201544
rect 673972 201532 673978 201544
rect 675386 201532 675392 201544
rect 673972 201504 675392 201532
rect 673972 201492 673978 201504
rect 675386 201492 675392 201504
rect 675444 201492 675450 201544
rect 674006 200676 674012 200728
rect 674064 200716 674070 200728
rect 675386 200716 675392 200728
rect 674064 200688 675392 200716
rect 674064 200676 674070 200688
rect 675386 200676 675392 200688
rect 675444 200676 675450 200728
rect 33042 200200 33048 200252
rect 33100 200240 33106 200252
rect 41874 200240 41880 200252
rect 33100 200212 41880 200240
rect 33100 200200 33106 200212
rect 41874 200200 41880 200212
rect 41932 200200 41938 200252
rect 581086 200064 581092 200116
rect 581144 200104 581150 200116
rect 599946 200104 599952 200116
rect 581144 200076 599952 200104
rect 581144 200064 581150 200076
rect 599946 200064 599952 200076
rect 600004 200064 600010 200116
rect 32950 199996 32956 200048
rect 33008 200036 33014 200048
rect 42518 200036 42524 200048
rect 33008 200008 42524 200036
rect 33008 199996 33014 200008
rect 42518 199996 42524 200008
rect 42576 199996 42582 200048
rect 582282 198704 582288 198756
rect 582340 198744 582346 198756
rect 599118 198744 599124 198756
rect 582340 198716 599124 198744
rect 582340 198704 582346 198716
rect 599118 198704 599124 198716
rect 599176 198704 599182 198756
rect 673638 198364 673644 198416
rect 673696 198404 673702 198416
rect 675386 198404 675392 198416
rect 673696 198376 675392 198404
rect 673696 198364 673702 198376
rect 675386 198364 675392 198376
rect 675444 198364 675450 198416
rect 673730 197548 673736 197600
rect 673788 197588 673794 197600
rect 675478 197588 675484 197600
rect 673788 197560 675484 197588
rect 673788 197548 673794 197560
rect 675478 197548 675484 197560
rect 675536 197548 675542 197600
rect 41874 197412 41880 197464
rect 41932 197412 41938 197464
rect 41892 197192 41920 197412
rect 582282 197344 582288 197396
rect 582340 197384 582346 197396
rect 599854 197384 599860 197396
rect 582340 197356 599860 197384
rect 582340 197344 582346 197356
rect 599854 197344 599860 197356
rect 599912 197344 599918 197396
rect 580718 197276 580724 197328
rect 580776 197316 580782 197328
rect 599946 197316 599952 197328
rect 580776 197288 599952 197316
rect 580776 197276 580782 197288
rect 599946 197276 599952 197288
rect 600004 197276 600010 197328
rect 41874 197140 41880 197192
rect 41932 197140 41938 197192
rect 673822 197004 673828 197056
rect 673880 197044 673886 197056
rect 675386 197044 675392 197056
rect 673880 197016 675392 197044
rect 673880 197004 673886 197016
rect 675386 197004 675392 197016
rect 675444 197004 675450 197056
rect 674650 196528 674656 196580
rect 674708 196568 674714 196580
rect 675386 196568 675392 196580
rect 674708 196540 675392 196568
rect 674708 196528 674714 196540
rect 675386 196528 675392 196540
rect 675444 196528 675450 196580
rect 674466 196392 674472 196444
rect 674524 196432 674530 196444
rect 674650 196432 674656 196444
rect 674524 196404 674656 196432
rect 674524 196392 674530 196404
rect 674650 196392 674656 196404
rect 674708 196392 674714 196444
rect 674834 195304 674840 195356
rect 674892 195344 674898 195356
rect 675386 195344 675392 195356
rect 674892 195316 675392 195344
rect 674892 195304 674898 195316
rect 675386 195304 675392 195316
rect 675444 195304 675450 195356
rect 42150 195236 42156 195288
rect 42208 195276 42214 195288
rect 42518 195276 42524 195288
rect 42208 195248 42524 195276
rect 42208 195236 42214 195248
rect 42518 195236 42524 195248
rect 42576 195236 42582 195288
rect 674374 195168 674380 195220
rect 674432 195208 674438 195220
rect 674834 195208 674840 195220
rect 674432 195180 674840 195208
rect 674432 195168 674438 195180
rect 674834 195168 674840 195180
rect 674892 195168 674898 195220
rect 582190 194624 582196 194676
rect 582248 194664 582254 194676
rect 599118 194664 599124 194676
rect 582248 194636 599124 194664
rect 582248 194624 582254 194636
rect 599118 194624 599124 194636
rect 599176 194624 599182 194676
rect 582282 194556 582288 194608
rect 582340 194596 582346 194608
rect 599946 194596 599952 194608
rect 582340 194568 599952 194596
rect 582340 194556 582346 194568
rect 599946 194556 599952 194568
rect 600004 194556 600010 194608
rect 42058 193468 42064 193520
rect 42116 193508 42122 193520
rect 42886 193508 42892 193520
rect 42116 193480 42892 193508
rect 42116 193468 42122 193480
rect 42886 193468 42892 193480
rect 42944 193468 42950 193520
rect 673454 193468 673460 193520
rect 673512 193508 673518 193520
rect 675386 193508 675392 193520
rect 673512 193480 675392 193508
rect 673512 193468 673518 193480
rect 675386 193468 675392 193480
rect 675444 193468 675450 193520
rect 42150 192176 42156 192228
rect 42208 192216 42214 192228
rect 42794 192216 42800 192228
rect 42208 192188 42800 192216
rect 42208 192176 42214 192188
rect 42794 192176 42800 192188
rect 42852 192176 42858 192228
rect 582190 191836 582196 191888
rect 582248 191876 582254 191888
rect 599118 191876 599124 191888
rect 582248 191848 599124 191876
rect 582248 191836 582254 191848
rect 599118 191836 599124 191848
rect 599176 191836 599182 191888
rect 582282 191768 582288 191820
rect 582340 191808 582346 191820
rect 599946 191808 599952 191820
rect 582340 191780 599952 191808
rect 582340 191768 582346 191780
rect 599946 191768 599952 191780
rect 600004 191768 600010 191820
rect 673546 191632 673552 191684
rect 673604 191672 673610 191684
rect 675386 191672 675392 191684
rect 673604 191644 675392 191672
rect 673604 191632 673610 191644
rect 675386 191632 675392 191644
rect 675444 191632 675450 191684
rect 42058 191428 42064 191480
rect 42116 191468 42122 191480
rect 43070 191468 43076 191480
rect 42116 191440 43076 191468
rect 42116 191428 42122 191440
rect 43070 191428 43076 191440
rect 43128 191428 43134 191480
rect 42150 190952 42156 191004
rect 42208 190992 42214 191004
rect 42978 190992 42984 191004
rect 42208 190964 42984 190992
rect 42208 190952 42214 190964
rect 42978 190952 42984 190964
rect 43036 190952 43042 191004
rect 579798 190408 579804 190460
rect 579856 190448 579862 190460
rect 599854 190448 599860 190460
rect 579856 190420 599860 190448
rect 579856 190408 579862 190420
rect 599854 190408 599860 190420
rect 599912 190408 599918 190460
rect 582190 187620 582196 187672
rect 582248 187660 582254 187672
rect 601602 187660 601608 187672
rect 582248 187632 601608 187660
rect 582248 187620 582254 187632
rect 601602 187620 601608 187632
rect 601660 187620 601666 187672
rect 582282 187552 582288 187604
rect 582340 187592 582346 187604
rect 600958 187592 600964 187604
rect 582340 187564 600964 187592
rect 582340 187552 582346 187564
rect 600958 187552 600964 187564
rect 601016 187552 601022 187604
rect 580258 184832 580264 184884
rect 580316 184872 580322 184884
rect 599946 184872 599952 184884
rect 580316 184844 599952 184872
rect 580316 184832 580322 184844
rect 599946 184832 599952 184844
rect 600004 184832 600010 184884
rect 580902 184764 580908 184816
rect 580960 184804 580966 184816
rect 601418 184804 601424 184816
rect 580960 184776 601424 184804
rect 580960 184764 580966 184776
rect 601418 184764 601424 184776
rect 601476 184764 601482 184816
rect 666646 183880 666652 183932
rect 666704 183920 666710 183932
rect 667014 183920 667020 183932
rect 666704 183892 667020 183920
rect 666704 183880 666710 183892
rect 667014 183880 667020 183892
rect 667072 183880 667078 183932
rect 580626 182112 580632 182164
rect 580684 182152 580690 182164
rect 600038 182152 600044 182164
rect 580684 182124 600044 182152
rect 580684 182112 580690 182124
rect 600038 182112 600044 182124
rect 600096 182112 600102 182164
rect 580534 182044 580540 182096
rect 580592 182084 580598 182096
rect 599854 182084 599860 182096
rect 580592 182056 599860 182084
rect 580592 182044 580598 182056
rect 599854 182044 599860 182056
rect 599912 182044 599918 182096
rect 580718 179324 580724 179376
rect 580776 179364 580782 179376
rect 599946 179364 599952 179376
rect 580776 179336 599952 179364
rect 580776 179324 580782 179336
rect 599946 179324 599952 179336
rect 600004 179324 600010 179376
rect 666830 179324 666836 179376
rect 666888 179364 666894 179376
rect 671430 179364 671436 179376
rect 666888 179336 671436 179364
rect 666888 179324 666894 179336
rect 671430 179324 671436 179336
rect 671488 179324 671494 179376
rect 674742 179324 674748 179376
rect 674800 179364 674806 179376
rect 675846 179364 675852 179376
rect 674800 179336 675852 179364
rect 674800 179324 674806 179336
rect 675846 179324 675852 179336
rect 675904 179324 675910 179376
rect 581086 179256 581092 179308
rect 581144 179296 581150 179308
rect 599762 179296 599768 179308
rect 581144 179268 599768 179296
rect 581144 179256 581150 179268
rect 599762 179256 599768 179268
rect 599820 179256 599826 179308
rect 669498 177080 669504 177132
rect 669556 177120 669562 177132
rect 675938 177120 675944 177132
rect 669556 177092 675944 177120
rect 669556 177080 669562 177092
rect 675938 177080 675944 177092
rect 675996 177080 676002 177132
rect 669130 176944 669136 176996
rect 669188 176984 669194 176996
rect 676030 176984 676036 176996
rect 669188 176956 676036 176984
rect 669188 176944 669194 176956
rect 676030 176944 676036 176956
rect 676088 176944 676094 176996
rect 671430 176876 671436 176928
rect 671488 176916 671494 176928
rect 673270 176916 673276 176928
rect 671488 176888 673276 176916
rect 671488 176876 671494 176888
rect 673270 176876 673276 176888
rect 673328 176916 673334 176928
rect 675938 176916 675944 176928
rect 673328 176888 675944 176916
rect 673328 176876 673334 176888
rect 675938 176876 675944 176888
rect 675996 176876 676002 176928
rect 666922 176808 666928 176860
rect 666980 176848 666986 176860
rect 675754 176848 675760 176860
rect 666980 176820 675760 176848
rect 666980 176808 666986 176820
rect 675754 176808 675760 176820
rect 675812 176808 675818 176860
rect 580994 176672 581000 176724
rect 581052 176712 581058 176724
rect 598934 176712 598940 176724
rect 581052 176684 598940 176712
rect 581052 176672 581058 176684
rect 598934 176672 598940 176684
rect 598992 176672 598998 176724
rect 581454 176604 581460 176656
rect 581512 176644 581518 176656
rect 600038 176644 600044 176656
rect 581512 176616 600044 176644
rect 581512 176604 581518 176616
rect 600038 176604 600044 176616
rect 600096 176604 600102 176656
rect 666738 176604 666744 176656
rect 666796 176644 666802 176656
rect 671338 176644 671344 176656
rect 666796 176616 671344 176644
rect 666796 176604 666802 176616
rect 671338 176604 671344 176616
rect 671396 176604 671402 176656
rect 674834 176604 674840 176656
rect 674892 176644 674898 176656
rect 676030 176644 676036 176656
rect 674892 176616 676036 176644
rect 674892 176604 674898 176616
rect 676030 176604 676036 176616
rect 676088 176604 676094 176656
rect 667014 176536 667020 176588
rect 667072 176576 667078 176588
rect 672166 176576 672172 176588
rect 667072 176548 672172 176576
rect 667072 176536 667078 176548
rect 672166 176536 672172 176548
rect 672224 176536 672230 176588
rect 674650 176332 674656 176384
rect 674708 176372 674714 176384
rect 676030 176372 676036 176384
rect 674708 176344 676036 176372
rect 674708 176332 674714 176344
rect 676030 176332 676036 176344
rect 676088 176332 676094 176384
rect 673362 175992 673368 176044
rect 673420 176032 673426 176044
rect 675938 176032 675944 176044
rect 673420 176004 675944 176032
rect 673420 175992 673426 176004
rect 675938 175992 675944 176004
rect 675996 175992 676002 176044
rect 674558 175516 674564 175568
rect 674616 175556 674622 175568
rect 676030 175556 676036 175568
rect 674616 175528 676036 175556
rect 674616 175516 674622 175528
rect 676030 175516 676036 175528
rect 676088 175516 676094 175568
rect 671338 175244 671344 175296
rect 671396 175284 671402 175296
rect 672258 175284 672264 175296
rect 671396 175256 672264 175284
rect 671396 175244 671402 175256
rect 672258 175244 672264 175256
rect 672316 175284 672322 175296
rect 675938 175284 675944 175296
rect 672316 175256 675944 175284
rect 672316 175244 672322 175256
rect 675938 175244 675944 175256
rect 675996 175244 676002 175296
rect 671890 174428 671896 174480
rect 671948 174468 671954 174480
rect 672166 174468 672172 174480
rect 671948 174440 672172 174468
rect 671948 174428 671954 174440
rect 672166 174428 672172 174440
rect 672224 174468 672230 174480
rect 676030 174468 676036 174480
rect 672224 174440 676036 174468
rect 672224 174428 672230 174440
rect 676030 174428 676036 174440
rect 676088 174428 676094 174480
rect 580810 173884 580816 173936
rect 580868 173924 580874 173936
rect 599946 173924 599952 173936
rect 580868 173896 599952 173924
rect 580868 173884 580874 173896
rect 599946 173884 599952 173896
rect 600004 173884 600010 173936
rect 674098 173884 674104 173936
rect 674156 173924 674162 173936
rect 676030 173924 676036 173936
rect 674156 173896 676036 173924
rect 674156 173884 674162 173896
rect 676030 173884 676036 173896
rect 676088 173884 676094 173936
rect 579706 173816 579712 173868
rect 579764 173856 579770 173868
rect 599854 173856 599860 173868
rect 579764 173828 599860 173856
rect 579764 173816 579770 173828
rect 599854 173816 599860 173828
rect 599912 173816 599918 173868
rect 582282 173748 582288 173800
rect 582340 173788 582346 173800
rect 600130 173788 600136 173800
rect 582340 173760 600136 173788
rect 582340 173748 582346 173760
rect 600130 173748 600136 173760
rect 600188 173748 600194 173800
rect 674650 171640 674656 171692
rect 674708 171680 674714 171692
rect 676030 171680 676036 171692
rect 674708 171652 676036 171680
rect 674708 171640 674714 171652
rect 676030 171640 676036 171652
rect 676088 171640 676094 171692
rect 673730 171300 673736 171352
rect 673788 171340 673794 171352
rect 675938 171340 675944 171352
rect 673788 171312 675944 171340
rect 673788 171300 673794 171312
rect 675938 171300 675944 171312
rect 675996 171300 676002 171352
rect 582190 171164 582196 171216
rect 582248 171204 582254 171216
rect 599946 171204 599952 171216
rect 582248 171176 599952 171204
rect 582248 171164 582254 171176
rect 599946 171164 599952 171176
rect 600004 171164 600010 171216
rect 674558 171164 674564 171216
rect 674616 171204 674622 171216
rect 675938 171204 675944 171216
rect 674616 171176 675944 171204
rect 674616 171164 674622 171176
rect 675938 171164 675944 171176
rect 675996 171164 676002 171216
rect 579890 171096 579896 171148
rect 579948 171136 579954 171148
rect 599854 171136 599860 171148
rect 579948 171108 599860 171136
rect 579948 171096 579954 171108
rect 599854 171096 599860 171108
rect 599912 171096 599918 171148
rect 674834 171096 674840 171148
rect 674892 171136 674898 171148
rect 676030 171136 676036 171148
rect 674892 171108 676036 171136
rect 674892 171096 674898 171108
rect 676030 171096 676036 171108
rect 676088 171096 676094 171148
rect 582006 171028 582012 171080
rect 582064 171068 582070 171080
rect 599762 171068 599768 171080
rect 582064 171040 599768 171068
rect 582064 171028 582070 171040
rect 599762 171028 599768 171040
rect 599820 171028 599826 171080
rect 580534 170960 580540 171012
rect 580592 171000 580598 171012
rect 599670 171000 599676 171012
rect 580592 170972 599676 171000
rect 580592 170960 580598 170972
rect 599670 170960 599676 170972
rect 599728 170960 599734 171012
rect 673454 170008 673460 170060
rect 673512 170048 673518 170060
rect 675938 170048 675944 170060
rect 673512 170020 675944 170048
rect 673512 170008 673518 170020
rect 675938 170008 675944 170020
rect 675996 170008 676002 170060
rect 673638 169192 673644 169244
rect 673696 169232 673702 169244
rect 675938 169232 675944 169244
rect 673696 169204 675944 169232
rect 673696 169192 673702 169204
rect 675938 169192 675944 169204
rect 675996 169192 676002 169244
rect 673822 168716 673828 168768
rect 673880 168756 673886 168768
rect 675938 168756 675944 168768
rect 673880 168728 675944 168756
rect 673880 168716 673886 168728
rect 675938 168716 675944 168728
rect 675996 168716 676002 168768
rect 674742 168648 674748 168700
rect 674800 168688 674806 168700
rect 676030 168688 676036 168700
rect 674800 168660 676036 168688
rect 674800 168648 674806 168660
rect 676030 168648 676036 168660
rect 676088 168648 676094 168700
rect 579706 168512 579712 168564
rect 579764 168552 579770 168564
rect 599946 168552 599952 168564
rect 579764 168524 599952 168552
rect 579764 168512 579770 168524
rect 599946 168512 599952 168524
rect 600004 168512 600010 168564
rect 673546 168512 673552 168564
rect 673604 168552 673610 168564
rect 675846 168552 675852 168564
rect 673604 168524 675852 168552
rect 673604 168512 673610 168524
rect 675846 168512 675852 168524
rect 675904 168512 675910 168564
rect 582098 168444 582104 168496
rect 582156 168484 582162 168496
rect 599026 168484 599032 168496
rect 582156 168456 599032 168484
rect 582156 168444 582162 168456
rect 599026 168444 599032 168456
rect 599084 168444 599090 168496
rect 580166 168376 580172 168428
rect 580224 168416 580230 168428
rect 599762 168416 599768 168428
rect 580224 168388 599768 168416
rect 580224 168376 580230 168388
rect 599762 168376 599768 168388
rect 599820 168376 599826 168428
rect 582282 168308 582288 168360
rect 582340 168348 582346 168360
rect 600314 168348 600320 168360
rect 582340 168320 600320 168348
rect 582340 168308 582346 168320
rect 600314 168308 600320 168320
rect 600372 168308 600378 168360
rect 672166 168240 672172 168292
rect 672224 168280 672230 168292
rect 676030 168280 676036 168292
rect 672224 168252 676036 168280
rect 672224 168240 672230 168252
rect 676030 168240 676036 168252
rect 676088 168240 676094 168292
rect 672350 167832 672356 167884
rect 672408 167872 672414 167884
rect 676030 167872 676036 167884
rect 672408 167844 676036 167872
rect 672408 167832 672414 167844
rect 676030 167832 676036 167844
rect 676088 167832 676094 167884
rect 672074 167016 672080 167068
rect 672132 167056 672138 167068
rect 676030 167056 676036 167068
rect 672132 167028 676036 167056
rect 672132 167016 672138 167028
rect 676030 167016 676036 167028
rect 676088 167016 676094 167068
rect 581270 165724 581276 165776
rect 581328 165764 581334 165776
rect 599854 165764 599860 165776
rect 581328 165736 599860 165764
rect 581328 165724 581334 165736
rect 599854 165724 599860 165736
rect 599912 165724 599918 165776
rect 580350 165656 580356 165708
rect 580408 165696 580414 165708
rect 600038 165696 600044 165708
rect 580408 165668 600044 165696
rect 580408 165656 580414 165668
rect 600038 165656 600044 165668
rect 600096 165656 600102 165708
rect 581914 165588 581920 165640
rect 581972 165628 581978 165640
rect 599946 165628 599952 165640
rect 581972 165600 599952 165628
rect 581972 165588 581978 165600
rect 599946 165588 599952 165600
rect 600004 165588 600010 165640
rect 581822 165520 581828 165572
rect 581880 165560 581886 165572
rect 601142 165560 601148 165572
rect 581880 165532 601148 165560
rect 581880 165520 581886 165532
rect 601142 165520 601148 165532
rect 601200 165520 601206 165572
rect 581454 162936 581460 162988
rect 581512 162976 581518 162988
rect 599854 162976 599860 162988
rect 581512 162948 599860 162976
rect 581512 162936 581518 162948
rect 599854 162936 599860 162948
rect 599912 162936 599918 162988
rect 580994 162868 581000 162920
rect 581052 162908 581058 162920
rect 599946 162908 599952 162920
rect 581052 162880 599952 162908
rect 581052 162868 581058 162880
rect 599946 162868 599952 162880
rect 600004 162868 600010 162920
rect 675754 160964 675760 161016
rect 675812 160964 675818 161016
rect 675772 160812 675800 160964
rect 675754 160760 675760 160812
rect 675812 160760 675818 160812
rect 581178 160216 581184 160268
rect 581236 160256 581242 160268
rect 600038 160256 600044 160268
rect 581236 160228 600044 160256
rect 581236 160216 581242 160228
rect 600038 160216 600044 160228
rect 600096 160216 600102 160268
rect 580902 160148 580908 160200
rect 580960 160188 580966 160200
rect 599946 160188 599952 160200
rect 580960 160160 599952 160188
rect 580960 160148 580966 160160
rect 599946 160148 599952 160160
rect 600004 160148 600010 160200
rect 580534 160080 580540 160132
rect 580592 160120 580598 160132
rect 599854 160120 599860 160132
rect 580592 160092 599860 160120
rect 580592 160080 580598 160092
rect 599854 160080 599860 160092
rect 599912 160080 599918 160132
rect 674834 159876 674840 159928
rect 674892 159916 674898 159928
rect 675386 159916 675392 159928
rect 674892 159888 675392 159916
rect 674892 159876 674898 159888
rect 675386 159876 675392 159888
rect 675444 159876 675450 159928
rect 674098 159332 674104 159384
rect 674156 159372 674162 159384
rect 675478 159372 675484 159384
rect 674156 159344 675484 159372
rect 674156 159332 674162 159344
rect 675478 159332 675484 159344
rect 675536 159332 675542 159384
rect 674650 157700 674656 157752
rect 674708 157740 674714 157752
rect 675478 157740 675484 157752
rect 674708 157712 675484 157740
rect 674708 157700 674714 157712
rect 675478 157700 675484 157712
rect 675536 157700 675542 157752
rect 582006 157496 582012 157548
rect 582064 157536 582070 157548
rect 599946 157536 599952 157548
rect 582064 157508 599952 157536
rect 582064 157496 582070 157508
rect 599946 157496 599952 157508
rect 600004 157496 600010 157548
rect 581086 157428 581092 157480
rect 581144 157468 581150 157480
rect 599854 157468 599860 157480
rect 581144 157440 599860 157468
rect 581144 157428 581150 157440
rect 599854 157428 599860 157440
rect 599912 157428 599918 157480
rect 580810 157360 580816 157412
rect 580868 157400 580874 157412
rect 598934 157400 598940 157412
rect 580868 157372 598940 157400
rect 580868 157360 580874 157372
rect 598934 157360 598940 157372
rect 598992 157360 598998 157412
rect 674558 156884 674564 156936
rect 674616 156924 674622 156936
rect 675386 156924 675392 156936
rect 674616 156896 675392 156924
rect 674616 156884 674622 156896
rect 675386 156884 675392 156896
rect 675444 156884 675450 156936
rect 674742 155660 674748 155712
rect 674800 155700 674806 155712
rect 675478 155700 675484 155712
rect 674800 155672 675484 155700
rect 674800 155660 674806 155672
rect 675478 155660 675484 155672
rect 675536 155660 675542 155712
rect 582190 154640 582196 154692
rect 582248 154680 582254 154692
rect 599946 154680 599952 154692
rect 582248 154652 599952 154680
rect 582248 154640 582254 154652
rect 599946 154640 599952 154652
rect 600004 154640 600010 154692
rect 580718 154572 580724 154624
rect 580776 154612 580782 154624
rect 599854 154612 599860 154624
rect 580776 154584 599860 154612
rect 580776 154572 580782 154584
rect 599854 154572 599860 154584
rect 599912 154572 599918 154624
rect 673730 153348 673736 153400
rect 673788 153388 673794 153400
rect 675386 153388 675392 153400
rect 673788 153360 675392 153388
rect 673788 153348 673794 153360
rect 675386 153348 675392 153360
rect 675444 153348 675450 153400
rect 673822 152532 673828 152584
rect 673880 152572 673886 152584
rect 675386 152572 675392 152584
rect 673880 152544 675392 152572
rect 673880 152532 673886 152544
rect 675386 152532 675392 152544
rect 675444 152532 675450 152584
rect 673638 151988 673644 152040
rect 673696 152028 673702 152040
rect 675386 152028 675392 152040
rect 673696 152000 675392 152028
rect 673696 151988 673702 152000
rect 675386 151988 675392 152000
rect 675444 151988 675450 152040
rect 582282 151920 582288 151972
rect 582340 151960 582346 151972
rect 599854 151960 599860 151972
rect 582340 151932 599860 151960
rect 582340 151920 582346 151932
rect 599854 151920 599860 151932
rect 599912 151920 599918 151972
rect 581822 151852 581828 151904
rect 581880 151892 581886 151904
rect 599946 151892 599952 151904
rect 581880 151864 599952 151892
rect 581880 151852 581886 151864
rect 599946 151852 599952 151864
rect 600004 151852 600010 151904
rect 582098 151784 582104 151836
rect 582156 151824 582162 151836
rect 600038 151824 600044 151836
rect 582156 151796 600044 151824
rect 582156 151784 582162 151796
rect 600038 151784 600044 151796
rect 600096 151784 600102 151836
rect 673546 151376 673552 151428
rect 673604 151416 673610 151428
rect 675386 151416 675392 151428
rect 673604 151388 675392 151416
rect 673604 151376 673610 151388
rect 675386 151376 675392 151388
rect 675444 151376 675450 151428
rect 673454 150356 673460 150408
rect 673512 150396 673518 150408
rect 675386 150396 675392 150408
rect 673512 150368 675392 150396
rect 673512 150356 673518 150368
rect 675386 150356 675392 150368
rect 675444 150356 675450 150408
rect 581914 149200 581920 149252
rect 581972 149240 581978 149252
rect 598934 149240 598940 149252
rect 581972 149212 598940 149240
rect 581972 149200 581978 149212
rect 598934 149200 598940 149212
rect 598992 149200 598998 149252
rect 581546 149132 581552 149184
rect 581604 149172 581610 149184
rect 599854 149172 599860 149184
rect 581604 149144 599860 149172
rect 581604 149132 581610 149144
rect 599854 149132 599860 149144
rect 599912 149132 599918 149184
rect 581362 149064 581368 149116
rect 581420 149104 581426 149116
rect 599946 149104 599952 149116
rect 581420 149076 599952 149104
rect 581420 149064 581426 149076
rect 599946 149064 599952 149076
rect 600004 149064 600010 149116
rect 581454 146344 581460 146396
rect 581512 146384 581518 146396
rect 599946 146384 599952 146396
rect 581512 146356 599952 146384
rect 581512 146344 581518 146356
rect 599946 146344 599952 146356
rect 600004 146344 600010 146396
rect 580626 146276 580632 146328
rect 580684 146316 580690 146328
rect 599854 146316 599860 146328
rect 580684 146288 599860 146316
rect 580684 146276 580690 146288
rect 599854 146276 599860 146288
rect 599912 146276 599918 146328
rect 581730 143692 581736 143744
rect 581788 143732 581794 143744
rect 599946 143732 599952 143744
rect 581788 143704 599952 143732
rect 581788 143692 581794 143704
rect 599946 143692 599952 143704
rect 600004 143692 600010 143744
rect 581270 143624 581276 143676
rect 581328 143664 581334 143676
rect 599854 143664 599860 143676
rect 581328 143636 599860 143664
rect 581328 143624 581334 143636
rect 599854 143624 599860 143636
rect 599912 143624 599918 143676
rect 579706 143556 579712 143608
rect 579764 143596 579770 143608
rect 600038 143596 600044 143608
rect 579764 143568 600044 143596
rect 579764 143556 579770 143568
rect 600038 143556 600044 143568
rect 600096 143556 600102 143608
rect 581638 140904 581644 140956
rect 581696 140944 581702 140956
rect 599854 140944 599860 140956
rect 581696 140916 599860 140944
rect 581696 140904 581702 140916
rect 599854 140904 599860 140916
rect 599912 140904 599918 140956
rect 580994 140836 581000 140888
rect 581052 140876 581058 140888
rect 599946 140876 599952 140888
rect 581052 140848 599952 140876
rect 581052 140836 581058 140848
rect 599946 140836 599952 140848
rect 600004 140836 600010 140888
rect 581178 140768 581184 140820
rect 581236 140808 581242 140820
rect 599302 140808 599308 140820
rect 581236 140780 599308 140808
rect 581236 140768 581242 140780
rect 599302 140768 599308 140780
rect 599360 140768 599366 140820
rect 581086 138116 581092 138168
rect 581144 138156 581150 138168
rect 599946 138156 599952 138168
rect 581144 138128 599952 138156
rect 581144 138116 581150 138128
rect 599946 138116 599952 138128
rect 600004 138116 600010 138168
rect 579798 138048 579804 138100
rect 579856 138088 579862 138100
rect 599854 138088 599860 138100
rect 579856 138060 599860 138088
rect 579856 138048 579862 138060
rect 599854 138048 599860 138060
rect 599912 138048 599918 138100
rect 580074 137980 580080 138032
rect 580132 138020 580138 138032
rect 599762 138020 599768 138032
rect 580132 137992 599768 138020
rect 580132 137980 580138 137992
rect 599762 137980 599768 137992
rect 599820 137980 599826 138032
rect 580166 135328 580172 135380
rect 580224 135368 580230 135380
rect 599946 135368 599952 135380
rect 580224 135340 599952 135368
rect 580224 135328 580230 135340
rect 599946 135328 599952 135340
rect 600004 135328 600010 135380
rect 579890 135260 579896 135312
rect 579948 135300 579954 135312
rect 599854 135300 599860 135312
rect 579948 135272 599860 135300
rect 579948 135260 579954 135272
rect 599854 135260 599860 135272
rect 599912 135260 599918 135312
rect 670510 132880 670516 132932
rect 670568 132920 670574 132932
rect 676214 132920 676220 132932
rect 670568 132892 676220 132920
rect 670568 132880 670574 132892
rect 676214 132880 676220 132892
rect 676272 132880 676278 132932
rect 669590 132744 669596 132796
rect 669648 132784 669654 132796
rect 676122 132784 676128 132796
rect 669648 132756 676128 132784
rect 669648 132744 669654 132756
rect 676122 132744 676128 132756
rect 676180 132744 676186 132796
rect 580902 132608 580908 132660
rect 580960 132648 580966 132660
rect 599854 132648 599860 132660
rect 580960 132620 599860 132648
rect 580960 132608 580966 132620
rect 599854 132608 599860 132620
rect 599912 132608 599918 132660
rect 669406 132608 669412 132660
rect 669464 132648 669470 132660
rect 676030 132648 676036 132660
rect 669464 132620 676036 132648
rect 669464 132608 669470 132620
rect 676030 132608 676036 132620
rect 676088 132608 676094 132660
rect 580258 132540 580264 132592
rect 580316 132580 580322 132592
rect 599946 132580 599952 132592
rect 580316 132552 599952 132580
rect 580316 132540 580322 132552
rect 599946 132540 599952 132552
rect 600004 132540 600010 132592
rect 579982 132472 579988 132524
rect 580040 132512 580046 132524
rect 600038 132512 600044 132524
rect 580040 132484 600044 132512
rect 580040 132472 580046 132484
rect 600038 132472 600044 132484
rect 600096 132472 600102 132524
rect 673270 132268 673276 132320
rect 673328 132308 673334 132320
rect 676214 132308 676220 132320
rect 673328 132280 676220 132308
rect 673328 132268 673334 132280
rect 676214 132268 676220 132280
rect 676272 132268 676278 132320
rect 670786 131656 670792 131708
rect 670844 131696 670850 131708
rect 676030 131696 676036 131708
rect 670844 131668 676036 131696
rect 670844 131656 670850 131668
rect 676030 131656 676036 131668
rect 676088 131656 676094 131708
rect 673362 131452 673368 131504
rect 673420 131492 673426 131504
rect 676214 131492 676220 131504
rect 673420 131464 676220 131492
rect 673420 131452 673426 131464
rect 676214 131452 676220 131464
rect 676272 131452 676278 131504
rect 672442 130840 672448 130892
rect 672500 130880 672506 130892
rect 676030 130880 676036 130892
rect 672500 130852 676036 130880
rect 672500 130840 672506 130852
rect 676030 130840 676036 130852
rect 676088 130840 676094 130892
rect 672258 130636 672264 130688
rect 672316 130676 672322 130688
rect 676214 130676 676220 130688
rect 672316 130648 676220 130676
rect 672316 130636 672322 130648
rect 676214 130636 676220 130648
rect 676272 130636 676278 130688
rect 670878 130024 670884 130076
rect 670936 130064 670942 130076
rect 676030 130064 676036 130076
rect 670936 130036 676036 130064
rect 670936 130024 670942 130036
rect 676030 130024 676036 130036
rect 676088 130024 676094 130076
rect 580718 129888 580724 129940
rect 580776 129928 580782 129940
rect 599762 129928 599768 129940
rect 580776 129900 599768 129928
rect 580776 129888 580782 129900
rect 599762 129888 599768 129900
rect 599820 129888 599826 129940
rect 580350 129820 580356 129872
rect 580408 129860 580414 129872
rect 599854 129860 599860 129872
rect 580408 129832 599860 129860
rect 580408 129820 580414 129832
rect 599854 129820 599860 129832
rect 599912 129820 599918 129872
rect 669314 129820 669320 129872
rect 669372 129860 669378 129872
rect 670786 129860 670792 129872
rect 669372 129832 670792 129860
rect 669372 129820 669378 129832
rect 670786 129820 670792 129832
rect 670844 129820 670850 129872
rect 580534 129752 580540 129804
rect 580592 129792 580598 129804
rect 599946 129792 599952 129804
rect 580592 129764 599952 129792
rect 580592 129752 580598 129764
rect 599946 129752 599952 129764
rect 600004 129752 600010 129804
rect 669222 129752 669228 129804
rect 669280 129792 669286 129804
rect 670878 129792 670884 129804
rect 669280 129764 670884 129792
rect 669280 129752 669286 129764
rect 670878 129752 670884 129764
rect 670936 129752 670942 129804
rect 671890 129684 671896 129736
rect 671948 129724 671954 129736
rect 676030 129724 676036 129736
rect 671948 129696 676036 129724
rect 671948 129684 671954 129696
rect 676030 129684 676036 129696
rect 676088 129684 676094 129736
rect 671982 129412 671988 129464
rect 672040 129452 672046 129464
rect 676214 129452 676220 129464
rect 672040 129424 676220 129452
rect 672040 129412 672046 129424
rect 676214 129412 676220 129424
rect 676272 129412 676278 129464
rect 674374 127712 674380 127764
rect 674432 127752 674438 127764
rect 676030 127752 676036 127764
rect 674432 127724 676036 127752
rect 674432 127712 674438 127724
rect 676030 127712 676036 127724
rect 676088 127712 676094 127764
rect 580810 127032 580816 127084
rect 580868 127072 580874 127084
rect 599946 127072 599952 127084
rect 580868 127044 599952 127072
rect 580868 127032 580874 127044
rect 599946 127032 599952 127044
rect 600004 127032 600010 127084
rect 673638 127032 673644 127084
rect 673696 127072 673702 127084
rect 675938 127072 675944 127084
rect 673696 127044 675944 127072
rect 673696 127032 673702 127044
rect 675938 127032 675944 127044
rect 675996 127032 676002 127084
rect 580442 126964 580448 127016
rect 580500 127004 580506 127016
rect 599854 127004 599860 127016
rect 580500 126976 599860 127004
rect 580500 126964 580506 126976
rect 599854 126964 599860 126976
rect 599912 126964 599918 127016
rect 674558 126964 674564 127016
rect 674616 127004 674622 127016
rect 676030 127004 676036 127016
rect 674616 126976 676036 127004
rect 674616 126964 674622 126976
rect 676030 126964 676036 126976
rect 676088 126964 676094 127016
rect 673546 124516 673552 124568
rect 673604 124556 673610 124568
rect 675662 124556 675668 124568
rect 673604 124528 675668 124556
rect 673604 124516 673610 124528
rect 675662 124516 675668 124528
rect 675720 124516 675726 124568
rect 674742 124448 674748 124500
rect 674800 124488 674806 124500
rect 675938 124488 675944 124500
rect 674800 124460 675944 124488
rect 674800 124448 674806 124460
rect 675938 124448 675944 124460
rect 675996 124448 676002 124500
rect 674466 124380 674472 124432
rect 674524 124420 674530 124432
rect 675846 124420 675852 124432
rect 674524 124392 675852 124420
rect 674524 124380 674530 124392
rect 675846 124380 675852 124392
rect 675904 124380 675910 124432
rect 582282 124312 582288 124364
rect 582340 124352 582346 124364
rect 600038 124352 600044 124364
rect 582340 124324 600044 124352
rect 582340 124312 582346 124324
rect 600038 124312 600044 124324
rect 600096 124312 600102 124364
rect 674650 124312 674656 124364
rect 674708 124352 674714 124364
rect 676122 124352 676128 124364
rect 674708 124324 676128 124352
rect 674708 124312 674714 124324
rect 676122 124312 676128 124324
rect 676180 124312 676186 124364
rect 582006 124244 582012 124296
rect 582064 124284 582070 124296
rect 599946 124284 599952 124296
rect 582064 124256 599952 124284
rect 582064 124244 582070 124256
rect 599946 124244 599952 124256
rect 600004 124244 600010 124296
rect 675110 124244 675116 124296
rect 675168 124284 675174 124296
rect 675938 124284 675944 124296
rect 675168 124256 675944 124284
rect 675168 124244 675174 124256
rect 675938 124244 675944 124256
rect 675996 124244 676002 124296
rect 580626 124176 580632 124228
rect 580684 124216 580690 124228
rect 599762 124216 599768 124228
rect 580684 124188 599768 124216
rect 580684 124176 580690 124188
rect 599762 124176 599768 124188
rect 599820 124176 599826 124228
rect 675202 124176 675208 124228
rect 675260 124216 675266 124228
rect 676030 124216 676036 124228
rect 675260 124188 676036 124216
rect 675260 124176 675266 124188
rect 676030 124176 676036 124188
rect 676088 124176 676094 124228
rect 673822 123224 673828 123276
rect 673880 123264 673886 123276
rect 676030 123264 676036 123276
rect 673880 123236 676036 123264
rect 673880 123224 673886 123236
rect 676030 123224 676036 123236
rect 676088 123224 676094 123276
rect 672902 123088 672908 123140
rect 672960 123128 672966 123140
rect 676030 123128 676036 123140
rect 672960 123100 676036 123128
rect 672960 123088 672966 123100
rect 676030 123088 676036 123100
rect 676088 123088 676094 123140
rect 671614 122680 671620 122732
rect 671672 122720 671678 122732
rect 676030 122720 676036 122732
rect 671672 122692 676036 122720
rect 671672 122680 671678 122692
rect 676030 122680 676036 122692
rect 676088 122680 676094 122732
rect 672258 121864 672264 121916
rect 672316 121904 672322 121916
rect 676030 121904 676036 121916
rect 672316 121876 676036 121904
rect 672316 121864 672322 121876
rect 676030 121864 676036 121876
rect 676088 121864 676094 121916
rect 582098 121592 582104 121644
rect 582156 121632 582162 121644
rect 599854 121632 599860 121644
rect 582156 121604 599860 121632
rect 582156 121592 582162 121604
rect 599854 121592 599860 121604
rect 599912 121592 599918 121644
rect 581914 121524 581920 121576
rect 581972 121564 581978 121576
rect 599946 121564 599952 121576
rect 581972 121536 599952 121564
rect 581972 121524 581978 121536
rect 599946 121524 599952 121536
rect 600004 121524 600010 121576
rect 582190 121456 582196 121508
rect 582248 121496 582254 121508
rect 600038 121496 600044 121508
rect 582248 121468 600044 121496
rect 582248 121456 582254 121468
rect 600038 121456 600044 121468
rect 600096 121456 600102 121508
rect 673730 121456 673736 121508
rect 673788 121496 673794 121508
rect 675938 121496 675944 121508
rect 673788 121468 675944 121496
rect 673788 121456 673794 121468
rect 675938 121456 675944 121468
rect 675996 121456 676002 121508
rect 583662 118804 583668 118856
rect 583720 118844 583726 118856
rect 599946 118844 599952 118856
rect 583720 118816 599952 118844
rect 583720 118804 583726 118816
rect 599946 118804 599952 118816
rect 600004 118804 600010 118856
rect 581822 118736 581828 118788
rect 581880 118776 581886 118788
rect 600038 118776 600044 118788
rect 581880 118748 600044 118776
rect 581880 118736 581886 118748
rect 600038 118736 600044 118748
rect 600096 118736 600102 118788
rect 581546 118668 581552 118720
rect 581604 118708 581610 118720
rect 599854 118708 599860 118720
rect 581604 118680 599860 118708
rect 581604 118668 581610 118680
rect 599854 118668 599860 118680
rect 599912 118668 599918 118720
rect 581730 116016 581736 116068
rect 581788 116056 581794 116068
rect 599854 116056 599860 116068
rect 581788 116028 599860 116056
rect 581788 116016 581794 116028
rect 599854 116016 599860 116028
rect 599912 116016 599918 116068
rect 581270 115948 581276 116000
rect 581328 115988 581334 116000
rect 599946 115988 599952 116000
rect 581328 115960 599952 115988
rect 581328 115948 581334 115960
rect 599946 115948 599952 115960
rect 600004 115948 600010 116000
rect 675754 115744 675760 115796
rect 675812 115744 675818 115796
rect 675772 115592 675800 115744
rect 675754 115540 675760 115592
rect 675812 115540 675818 115592
rect 675202 114996 675208 115048
rect 675260 115036 675266 115048
rect 675386 115036 675392 115048
rect 675260 115008 675392 115036
rect 675260 114996 675266 115008
rect 675386 114996 675392 115008
rect 675444 114996 675450 115048
rect 674374 114180 674380 114232
rect 674432 114220 674438 114232
rect 675386 114220 675392 114232
rect 674432 114192 675392 114220
rect 674432 114180 674438 114192
rect 675386 114180 675392 114192
rect 675444 114180 675450 114232
rect 581638 113228 581644 113280
rect 581696 113268 581702 113280
rect 599946 113268 599952 113280
rect 581696 113240 599952 113268
rect 581696 113228 581702 113240
rect 599946 113228 599952 113240
rect 600004 113228 600010 113280
rect 581454 113160 581460 113212
rect 581512 113200 581518 113212
rect 599854 113200 599860 113212
rect 581512 113172 599860 113200
rect 581512 113160 581518 113172
rect 599854 113160 599860 113172
rect 599912 113160 599918 113212
rect 674558 112344 674564 112396
rect 674616 112384 674622 112396
rect 675386 112384 675392 112396
rect 674616 112356 675392 112384
rect 674616 112344 674622 112356
rect 675386 112344 675392 112356
rect 675444 112344 675450 112396
rect 674742 111868 674748 111920
rect 674800 111908 674806 111920
rect 675386 111908 675392 111920
rect 674800 111880 675392 111908
rect 674800 111868 674806 111880
rect 675386 111868 675392 111880
rect 675444 111868 675450 111920
rect 674650 111120 674656 111172
rect 674708 111160 674714 111172
rect 675386 111160 675392 111172
rect 674708 111132 675392 111160
rect 674708 111120 674714 111132
rect 675386 111120 675392 111132
rect 675444 111120 675450 111172
rect 675110 110644 675116 110696
rect 675168 110684 675174 110696
rect 675386 110684 675392 110696
rect 675168 110656 675392 110684
rect 675168 110644 675174 110656
rect 675386 110644 675392 110656
rect 675444 110644 675450 110696
rect 581362 110508 581368 110560
rect 581420 110548 581426 110560
rect 599946 110548 599952 110560
rect 581420 110520 599952 110548
rect 581420 110508 581426 110520
rect 599946 110508 599952 110520
rect 600004 110508 600010 110560
rect 580994 110440 581000 110492
rect 581052 110480 581058 110492
rect 599762 110480 599768 110492
rect 581052 110452 599768 110480
rect 581052 110440 581058 110452
rect 599762 110440 599768 110452
rect 599820 110440 599826 110492
rect 673638 108196 673644 108248
rect 673696 108236 673702 108248
rect 675478 108236 675484 108248
rect 673696 108208 675484 108236
rect 673696 108196 673702 108208
rect 675478 108196 675484 108208
rect 675536 108196 675542 108248
rect 581178 107652 581184 107704
rect 581236 107692 581242 107704
rect 599946 107692 599952 107704
rect 581236 107664 599952 107692
rect 581236 107652 581242 107664
rect 599946 107652 599952 107664
rect 600004 107652 600010 107704
rect 673822 107516 673828 107568
rect 673880 107556 673886 107568
rect 675386 107556 675392 107568
rect 673880 107528 675392 107556
rect 673880 107516 673886 107528
rect 675386 107516 675392 107528
rect 675444 107516 675450 107568
rect 673546 106972 673552 107024
rect 673604 107012 673610 107024
rect 675386 107012 675392 107024
rect 673604 106984 675392 107012
rect 673604 106972 673610 106984
rect 675386 106972 675392 106984
rect 675444 106972 675450 107024
rect 673730 106360 673736 106412
rect 673788 106400 673794 106412
rect 675386 106400 675392 106412
rect 673788 106372 675392 106400
rect 673788 106360 673794 106372
rect 675386 106360 675392 106372
rect 675444 106360 675450 106412
rect 674466 105136 674472 105188
rect 674524 105176 674530 105188
rect 675478 105176 675484 105188
rect 674524 105148 675484 105176
rect 674524 105136 674530 105148
rect 675478 105136 675484 105148
rect 675536 105136 675542 105188
rect 581086 104864 581092 104916
rect 581144 104904 581150 104916
rect 599946 104904 599952 104916
rect 581144 104876 599952 104904
rect 581144 104864 581150 104876
rect 599946 104864 599952 104876
rect 600004 104864 600010 104916
rect 657722 99764 657728 99816
rect 657780 99804 657786 99816
rect 660896 99804 660902 99816
rect 657780 99776 660902 99804
rect 657780 99764 657786 99776
rect 660896 99764 660902 99776
rect 660954 99764 660960 99816
rect 580902 99356 580908 99408
rect 580960 99396 580966 99408
rect 599946 99396 599952 99408
rect 580960 99368 599952 99396
rect 580960 99356 580966 99368
rect 599946 99356 599952 99368
rect 600004 99356 600010 99408
rect 633066 96568 633072 96620
rect 633124 96608 633130 96620
rect 635274 96608 635280 96620
rect 633124 96580 635280 96608
rect 633124 96568 633130 96580
rect 635274 96568 635280 96580
rect 635332 96568 635338 96620
rect 636286 96568 636292 96620
rect 636344 96608 636350 96620
rect 640978 96608 640984 96620
rect 636344 96580 640984 96608
rect 636344 96568 636350 96580
rect 640978 96568 640984 96580
rect 641036 96568 641042 96620
rect 655974 96568 655980 96620
rect 656032 96608 656038 96620
rect 659562 96608 659568 96620
rect 656032 96580 659568 96608
rect 656032 96568 656038 96580
rect 659562 96568 659568 96580
rect 659620 96568 659626 96620
rect 661862 96568 661868 96620
rect 661920 96608 661926 96620
rect 663058 96608 663064 96620
rect 661920 96580 663064 96608
rect 661920 96568 661926 96580
rect 663058 96568 663064 96580
rect 663116 96568 663122 96620
rect 633802 96500 633808 96552
rect 633860 96540 633866 96552
rect 636378 96540 636384 96552
rect 633860 96512 636384 96540
rect 633860 96500 633866 96512
rect 636378 96500 636384 96512
rect 636436 96500 636442 96552
rect 637022 96500 637028 96552
rect 637080 96540 637086 96552
rect 642358 96540 642364 96552
rect 637080 96512 642364 96540
rect 637080 96500 637086 96512
rect 642358 96500 642364 96512
rect 642416 96500 642422 96552
rect 654686 96500 654692 96552
rect 654744 96540 654750 96552
rect 658274 96540 658280 96552
rect 654744 96512 658280 96540
rect 654744 96500 654750 96512
rect 658274 96500 658280 96512
rect 658332 96500 658338 96552
rect 659102 96500 659108 96552
rect 659160 96540 659166 96552
rect 662506 96540 662512 96552
rect 659160 96512 662512 96540
rect 659160 96500 659166 96512
rect 662506 96500 662512 96512
rect 662564 96500 662570 96552
rect 634446 96432 634452 96484
rect 634504 96472 634510 96484
rect 637574 96472 637580 96484
rect 634504 96444 637580 96472
rect 634504 96432 634510 96444
rect 637574 96432 637580 96444
rect 637632 96432 637638 96484
rect 652018 96432 652024 96484
rect 652076 96472 652082 96484
rect 661954 96472 661960 96484
rect 652076 96444 661960 96472
rect 652076 96432 652082 96444
rect 661954 96432 661960 96444
rect 662012 96432 662018 96484
rect 635734 96364 635740 96416
rect 635792 96404 635798 96416
rect 639874 96404 639880 96416
rect 635792 96376 639880 96404
rect 635792 96364 635798 96376
rect 639874 96364 639880 96376
rect 639932 96364 639938 96416
rect 631134 96024 631140 96076
rect 631192 96064 631198 96076
rect 632100 96064 632106 96076
rect 631192 96036 632106 96064
rect 631192 96024 631198 96036
rect 632100 96024 632106 96036
rect 632158 96024 632164 96076
rect 632422 96024 632428 96076
rect 632480 96064 632486 96076
rect 634400 96064 634406 96076
rect 632480 96036 634406 96064
rect 632480 96024 632486 96036
rect 634400 96024 634406 96036
rect 634458 96024 634464 96076
rect 635090 96024 635096 96076
rect 635148 96064 635154 96076
rect 639000 96064 639006 96076
rect 635148 96036 639006 96064
rect 635148 96024 635154 96036
rect 639000 96024 639006 96036
rect 639058 96024 639064 96076
rect 647510 96024 647516 96076
rect 647568 96064 647574 96076
rect 652754 96064 652760 96076
rect 647568 96036 652760 96064
rect 647568 96024 647574 96036
rect 652754 96024 652760 96036
rect 652812 96024 652818 96076
rect 631778 95888 631784 95940
rect 631836 95928 631842 95940
rect 632974 95928 632980 95940
rect 631836 95900 632980 95928
rect 631836 95888 631842 95900
rect 632974 95888 632980 95900
rect 633032 95888 633038 95940
rect 640058 95888 640064 95940
rect 640116 95928 640122 95940
rect 646038 95928 646044 95940
rect 640116 95900 646044 95928
rect 640116 95888 640122 95900
rect 646038 95888 646044 95900
rect 646096 95888 646102 95940
rect 646774 95888 646780 95940
rect 646832 95928 646838 95940
rect 663334 95928 663340 95940
rect 646832 95900 663340 95928
rect 646832 95888 646838 95900
rect 663334 95888 663340 95900
rect 663392 95888 663398 95940
rect 638862 95820 638868 95872
rect 638920 95860 638926 95872
rect 646222 95860 646228 95872
rect 638920 95832 646228 95860
rect 638920 95820 638926 95832
rect 646222 95820 646228 95832
rect 646280 95820 646286 95872
rect 614758 95752 614764 95804
rect 614816 95792 614822 95804
rect 614816 95764 632054 95792
rect 614816 95752 614822 95764
rect 620002 95616 620008 95668
rect 620060 95656 620066 95668
rect 623498 95656 623504 95668
rect 620060 95628 623504 95656
rect 620060 95616 620066 95628
rect 623498 95616 623504 95628
rect 623556 95616 623562 95668
rect 607214 95548 607220 95600
rect 607272 95588 607278 95600
rect 608962 95588 608968 95600
rect 607272 95560 608968 95588
rect 607272 95548 607278 95560
rect 608962 95548 608968 95560
rect 609020 95548 609026 95600
rect 610250 95548 610256 95600
rect 610308 95588 610314 95600
rect 611538 95588 611544 95600
rect 610308 95560 611544 95588
rect 610308 95548 610314 95560
rect 611538 95548 611544 95560
rect 611596 95548 611602 95600
rect 613010 95548 613016 95600
rect 613068 95588 613074 95600
rect 614850 95588 614856 95600
rect 613068 95560 614856 95588
rect 613068 95548 613074 95560
rect 614850 95548 614856 95560
rect 614908 95548 614914 95600
rect 618254 95548 618260 95600
rect 618312 95588 618318 95600
rect 620094 95588 620100 95600
rect 618312 95560 620100 95588
rect 618312 95548 618318 95560
rect 620094 95548 620100 95560
rect 620152 95548 620158 95600
rect 621198 95548 621204 95600
rect 621256 95588 621262 95600
rect 622670 95588 622676 95600
rect 621256 95560 622676 95588
rect 621256 95548 621262 95560
rect 622670 95548 622676 95560
rect 622728 95548 622734 95600
rect 623774 95548 623780 95600
rect 623832 95588 623838 95600
rect 624602 95588 624608 95600
rect 623832 95560 624608 95588
rect 623832 95548 623838 95560
rect 624602 95548 624608 95560
rect 624660 95548 624666 95600
rect 621290 95480 621296 95532
rect 621348 95520 621354 95532
rect 623314 95520 623320 95532
rect 621348 95492 623320 95520
rect 621348 95480 621354 95492
rect 623314 95480 623320 95492
rect 623372 95480 623378 95532
rect 616138 95412 616144 95464
rect 616196 95452 616202 95464
rect 623222 95452 623228 95464
rect 616196 95424 623228 95452
rect 616196 95412 616202 95424
rect 623222 95412 623228 95424
rect 623280 95412 623286 95464
rect 596174 95344 596180 95396
rect 596232 95384 596238 95396
rect 612918 95384 612924 95396
rect 596232 95356 612924 95384
rect 596232 95344 596238 95356
rect 612918 95344 612924 95356
rect 612976 95344 612982 95396
rect 619358 95344 619364 95396
rect 619416 95384 619422 95396
rect 622118 95384 622124 95396
rect 619416 95356 622124 95384
rect 619416 95344 619422 95356
rect 622118 95344 622124 95356
rect 622176 95344 622182 95396
rect 578142 95276 578148 95328
rect 578200 95316 578206 95328
rect 606386 95316 606392 95328
rect 578200 95288 606392 95316
rect 578200 95276 578206 95288
rect 606386 95276 606392 95288
rect 606444 95276 606450 95328
rect 575658 95208 575664 95260
rect 575716 95248 575722 95260
rect 610342 95248 610348 95260
rect 575716 95220 610348 95248
rect 575716 95208 575722 95220
rect 610342 95208 610348 95220
rect 610400 95208 610406 95260
rect 618714 95208 618720 95260
rect 618772 95248 618778 95260
rect 622670 95248 622676 95260
rect 618772 95220 622676 95248
rect 618772 95208 618778 95220
rect 622670 95208 622676 95220
rect 622728 95208 622734 95260
rect 632026 95180 632054 95764
rect 639598 95752 639604 95804
rect 639656 95792 639662 95804
rect 645946 95792 645952 95804
rect 639656 95764 645952 95792
rect 639656 95752 639662 95764
rect 645946 95752 645952 95764
rect 646004 95752 646010 95804
rect 637482 95684 637488 95736
rect 637540 95724 637546 95736
rect 640518 95724 640524 95736
rect 637540 95696 640524 95724
rect 637540 95684 637546 95696
rect 640518 95684 640524 95696
rect 640576 95684 640582 95736
rect 640886 95684 640892 95736
rect 640944 95724 640950 95736
rect 645854 95724 645860 95736
rect 640944 95696 645860 95724
rect 640944 95684 640950 95696
rect 645854 95684 645860 95696
rect 645912 95684 645918 95736
rect 641622 95616 641628 95668
rect 641680 95656 641686 95668
rect 642818 95656 642824 95668
rect 641680 95628 642824 95656
rect 641680 95616 641686 95628
rect 642818 95616 642824 95628
rect 642876 95616 642882 95668
rect 652662 95616 652668 95668
rect 652720 95656 652726 95668
rect 663794 95656 663800 95668
rect 652720 95628 663800 95656
rect 652720 95616 652726 95628
rect 663794 95616 663800 95628
rect 663852 95616 663858 95668
rect 638310 95548 638316 95600
rect 638368 95548 638374 95600
rect 642266 95548 642272 95600
rect 642324 95588 642330 95600
rect 642910 95588 642916 95600
rect 642324 95560 642916 95588
rect 642324 95548 642330 95560
rect 642910 95548 642916 95560
rect 642968 95548 642974 95600
rect 646406 95548 646412 95600
rect 646464 95588 646470 95600
rect 648154 95588 648160 95600
rect 646464 95560 648160 95588
rect 646464 95548 646470 95560
rect 648154 95548 648160 95560
rect 648212 95548 648218 95600
rect 656986 95548 656992 95600
rect 657044 95588 657050 95600
rect 659194 95588 659200 95600
rect 657044 95560 659200 95588
rect 657044 95548 657050 95560
rect 659194 95548 659200 95560
rect 659252 95548 659258 95600
rect 638328 95520 638356 95548
rect 642726 95520 642732 95532
rect 638328 95492 642732 95520
rect 642726 95480 642732 95492
rect 642784 95480 642790 95532
rect 660574 95480 660580 95532
rect 660632 95520 660638 95532
rect 661402 95520 661408 95532
rect 660632 95492 661408 95520
rect 660632 95480 660638 95492
rect 661402 95480 661408 95492
rect 661460 95480 661466 95532
rect 648614 95344 648620 95396
rect 648672 95384 648678 95396
rect 650730 95384 650736 95396
rect 648672 95356 650736 95384
rect 648672 95344 648678 95356
rect 650730 95344 650736 95356
rect 650788 95344 650794 95396
rect 656618 95344 656624 95396
rect 656676 95384 656682 95396
rect 663150 95384 663156 95396
rect 656676 95356 663156 95384
rect 656676 95344 656682 95356
rect 663150 95344 663156 95356
rect 663208 95344 663214 95396
rect 646130 95276 646136 95328
rect 646188 95316 646194 95328
rect 663426 95316 663432 95328
rect 646188 95288 663432 95316
rect 646188 95276 646194 95288
rect 663426 95276 663432 95288
rect 663484 95276 663490 95328
rect 657078 95208 657084 95260
rect 657136 95248 657142 95260
rect 657906 95248 657912 95260
rect 657136 95220 657912 95248
rect 657136 95208 657142 95220
rect 657906 95208 657912 95220
rect 657964 95208 657970 95260
rect 665174 95180 665180 95192
rect 632026 95152 665180 95180
rect 665174 95140 665180 95152
rect 665232 95140 665238 95192
rect 617426 94936 617432 94988
rect 617484 94976 617490 94988
rect 623314 94976 623320 94988
rect 617484 94948 623320 94976
rect 617484 94936 617490 94948
rect 623314 94936 623320 94948
rect 623372 94936 623378 94988
rect 643094 94936 643100 94988
rect 643152 94976 643158 94988
rect 644842 94976 644848 94988
rect 643152 94948 644848 94976
rect 643152 94936 643158 94948
rect 644842 94936 644848 94948
rect 644900 94936 644906 94988
rect 645946 94868 645952 94920
rect 646004 94908 646010 94920
rect 646222 94908 646228 94920
rect 646004 94880 646228 94908
rect 646004 94868 646010 94880
rect 646222 94868 646228 94880
rect 646280 94868 646286 94920
rect 618070 94800 618076 94852
rect 618128 94840 618134 94852
rect 621934 94840 621940 94852
rect 618128 94812 621940 94840
rect 618128 94800 618134 94812
rect 621934 94800 621940 94812
rect 621992 94800 621998 94852
rect 651834 94800 651840 94852
rect 651892 94840 651898 94852
rect 653398 94840 653404 94852
rect 651892 94812 653404 94840
rect 651892 94800 651898 94812
rect 653398 94800 653404 94812
rect 653456 94800 653462 94852
rect 648706 94664 648712 94716
rect 648764 94704 648770 94716
rect 649442 94704 649448 94716
rect 648764 94676 649448 94704
rect 648764 94664 648770 94676
rect 649442 94664 649448 94676
rect 649500 94664 649506 94716
rect 653306 94664 653312 94716
rect 653364 94704 653370 94716
rect 663702 94704 663708 94716
rect 653364 94676 663708 94704
rect 653364 94664 653370 94676
rect 663702 94664 663708 94676
rect 663760 94664 663766 94716
rect 657262 94596 657268 94648
rect 657320 94636 657326 94648
rect 663518 94636 663524 94648
rect 657320 94608 663524 94636
rect 657320 94596 657326 94608
rect 663518 94596 663524 94608
rect 663576 94596 663582 94648
rect 616782 94528 616788 94580
rect 616840 94568 616846 94580
rect 623130 94568 623136 94580
rect 616840 94540 623136 94568
rect 616840 94528 616846 94540
rect 623130 94528 623136 94540
rect 623188 94528 623194 94580
rect 648890 94528 648896 94580
rect 648948 94568 648954 94580
rect 650086 94568 650092 94580
rect 648948 94540 650092 94568
rect 648948 94528 648954 94540
rect 650086 94528 650092 94540
rect 650144 94528 650150 94580
rect 656894 94528 656900 94580
rect 656952 94568 656958 94580
rect 658550 94568 658556 94580
rect 656952 94540 658556 94568
rect 656952 94528 656958 94540
rect 658550 94528 658556 94540
rect 658608 94528 658614 94580
rect 648062 94460 648068 94512
rect 648120 94500 648126 94512
rect 659838 94500 659844 94512
rect 648120 94472 659844 94500
rect 648120 94460 648126 94472
rect 659838 94460 659844 94472
rect 659896 94460 659902 94512
rect 660390 94460 660396 94512
rect 660448 94460 660454 94512
rect 643554 94188 643560 94240
rect 643612 94228 643618 94240
rect 660408 94228 660436 94460
rect 643612 94200 660436 94228
rect 643612 94188 643618 94200
rect 644198 94052 644204 94104
rect 644256 94092 644262 94104
rect 654042 94092 654048 94104
rect 644256 94064 654048 94092
rect 644256 94052 644262 94064
rect 654042 94052 654048 94064
rect 654100 94052 654106 94104
rect 649350 93984 649356 94036
rect 649408 94024 649414 94036
rect 656894 94024 656900 94036
rect 649408 93996 656900 94024
rect 649408 93984 649414 93996
rect 656894 93984 656900 93996
rect 656952 93984 656958 94036
rect 605742 93848 605748 93900
rect 605800 93888 605806 93900
rect 613562 93888 613568 93900
rect 605800 93860 613568 93888
rect 605800 93848 605806 93860
rect 613562 93848 613568 93860
rect 613620 93848 613626 93900
rect 644750 93848 644756 93900
rect 644808 93888 644814 93900
rect 652938 93888 652944 93900
rect 644808 93860 652944 93888
rect 644808 93848 644814 93860
rect 652938 93848 652944 93860
rect 652996 93848 653002 93900
rect 607306 93780 607312 93832
rect 607364 93820 607370 93832
rect 612182 93820 612188 93832
rect 607364 93792 612188 93820
rect 607364 93780 607370 93792
rect 612182 93780 612188 93792
rect 612240 93780 612246 93832
rect 609974 91100 609980 91112
rect 607232 91072 609980 91100
rect 601694 90992 601700 91044
rect 601752 91032 601758 91044
rect 607232 91032 607260 91072
rect 609974 91060 609980 91072
rect 610032 91060 610038 91112
rect 601752 91004 607260 91032
rect 601752 90992 601758 91004
rect 657078 88816 657084 88868
rect 657136 88856 657142 88868
rect 657998 88856 658004 88868
rect 657136 88828 658004 88856
rect 657136 88816 657142 88828
rect 657998 88816 658004 88828
rect 658056 88816 658062 88868
rect 659470 88816 659476 88868
rect 659528 88856 659534 88868
rect 663610 88856 663616 88868
rect 659528 88828 663616 88856
rect 659528 88816 659534 88828
rect 663610 88816 663616 88828
rect 663668 88816 663674 88868
rect 648890 85484 648896 85536
rect 648948 85524 648954 85536
rect 657722 85524 657728 85536
rect 648948 85496 657728 85524
rect 648948 85484 648954 85496
rect 657722 85484 657728 85496
rect 657780 85484 657786 85536
rect 651834 85416 651840 85468
rect 651892 85456 651898 85468
rect 658826 85456 658832 85468
rect 651892 85428 658832 85456
rect 651892 85416 651898 85428
rect 658826 85416 658832 85428
rect 658884 85416 658890 85468
rect 648706 85348 648712 85400
rect 648764 85388 648770 85400
rect 660666 85388 660672 85400
rect 648764 85360 660672 85388
rect 648764 85348 648770 85360
rect 660666 85348 660672 85360
rect 660724 85348 660730 85400
rect 648614 85280 648620 85332
rect 648672 85320 648678 85332
rect 657170 85320 657176 85332
rect 648672 85292 657176 85320
rect 648672 85280 648678 85292
rect 657170 85280 657176 85292
rect 657228 85280 657234 85332
rect 643094 85212 643100 85264
rect 643152 85252 643158 85264
rect 660114 85252 660120 85264
rect 643152 85224 660120 85252
rect 643152 85212 643158 85224
rect 660114 85212 660120 85224
rect 660172 85212 660178 85264
rect 646406 85144 646412 85196
rect 646464 85184 646470 85196
rect 661402 85184 661408 85196
rect 646464 85156 661408 85184
rect 646464 85144 646470 85156
rect 661402 85144 661408 85156
rect 661460 85144 661466 85196
rect 586422 84600 586428 84652
rect 586480 84640 586486 84652
rect 600314 84640 600320 84652
rect 586480 84612 600320 84640
rect 586480 84600 586486 84612
rect 600314 84600 600320 84612
rect 600372 84600 600378 84652
rect 583846 84532 583852 84584
rect 583904 84572 583910 84584
rect 600498 84572 600504 84584
rect 583904 84544 600504 84572
rect 583904 84532 583910 84544
rect 600498 84532 600504 84544
rect 600556 84532 600562 84584
rect 583754 84464 583760 84516
rect 583812 84504 583818 84516
rect 600682 84504 600688 84516
rect 583812 84476 600688 84504
rect 583812 84464 583818 84476
rect 600682 84464 600688 84476
rect 600740 84464 600746 84516
rect 582282 84396 582288 84448
rect 582340 84436 582346 84448
rect 600222 84436 600228 84448
rect 582340 84408 600228 84436
rect 582340 84396 582346 84408
rect 600222 84396 600228 84408
rect 600280 84396 600286 84448
rect 582190 84328 582196 84380
rect 582248 84368 582254 84380
rect 600406 84368 600412 84380
rect 582248 84340 600412 84368
rect 582248 84328 582254 84340
rect 600406 84328 600412 84340
rect 600464 84328 600470 84380
rect 582006 84260 582012 84312
rect 582064 84300 582070 84312
rect 600590 84300 600596 84312
rect 582064 84272 600596 84300
rect 582064 84260 582070 84272
rect 600590 84260 600596 84272
rect 600648 84260 600654 84312
rect 582098 84192 582104 84244
rect 582156 84232 582162 84244
rect 600774 84232 600780 84244
rect 582156 84204 600780 84232
rect 582156 84192 582162 84204
rect 600774 84192 600780 84204
rect 600832 84192 600838 84244
rect 581914 84124 581920 84176
rect 581972 84164 581978 84176
rect 600866 84164 600872 84176
rect 581972 84136 600872 84164
rect 581972 84124 581978 84136
rect 600866 84124 600872 84136
rect 600924 84124 600930 84176
rect 579614 82628 579620 82680
rect 579672 82668 579678 82680
rect 583662 82668 583668 82680
rect 579672 82640 583668 82668
rect 579672 82628 579678 82640
rect 583662 82628 583668 82640
rect 583720 82628 583726 82680
rect 591942 80792 591948 80844
rect 592000 80832 592006 80844
rect 596174 80832 596180 80844
rect 592000 80804 596180 80832
rect 592000 80792 592006 80804
rect 596174 80792 596180 80804
rect 596232 80792 596238 80844
rect 600222 78480 600228 78532
rect 600280 78520 600286 78532
rect 610342 78520 610348 78532
rect 600280 78492 610348 78520
rect 600280 78480 600286 78492
rect 610342 78480 610348 78492
rect 610400 78480 610406 78532
rect 605834 77800 605840 77852
rect 605892 77840 605898 77852
rect 607306 77840 607312 77852
rect 605892 77812 607312 77840
rect 605892 77800 605898 77812
rect 607306 77800 607312 77812
rect 607364 77800 607370 77852
rect 600038 74468 600044 74520
rect 600096 74508 600102 74520
rect 605742 74508 605748 74520
rect 600096 74480 605748 74508
rect 600096 74468 600102 74480
rect 605742 74468 605748 74480
rect 605800 74468 605806 74520
rect 590654 73108 590660 73160
rect 590712 73148 590718 73160
rect 601602 73148 601608 73160
rect 590712 73120 601608 73148
rect 590712 73108 590718 73120
rect 601602 73108 601608 73120
rect 601660 73108 601666 73160
rect 598934 69028 598940 69080
rect 598992 69068 598998 69080
rect 605834 69068 605840 69080
rect 598992 69040 605840 69068
rect 598992 69028 598998 69040
rect 605834 69028 605840 69040
rect 605892 69028 605898 69080
rect 583662 66240 583668 66292
rect 583720 66280 583726 66292
rect 590654 66280 590660 66292
rect 583720 66252 590660 66280
rect 583720 66240 583726 66252
rect 590654 66240 590660 66252
rect 590712 66240 590718 66292
rect 580534 66172 580540 66224
rect 580592 66212 580598 66224
rect 586422 66212 586428 66224
rect 580592 66184 586428 66212
rect 580592 66172 580598 66184
rect 586422 66172 586428 66184
rect 586480 66172 586486 66224
rect 590654 64812 590660 64864
rect 590712 64852 590718 64864
rect 600038 64852 600044 64864
rect 590712 64824 600044 64852
rect 590712 64812 590718 64824
rect 600038 64812 600044 64824
rect 600096 64812 600102 64864
rect 600314 63520 600320 63572
rect 600372 63560 600378 63572
rect 607490 63560 607496 63572
rect 600372 63532 607496 63560
rect 600372 63520 600378 63532
rect 607490 63520 607496 63532
rect 607548 63520 607554 63572
rect 590746 62092 590752 62144
rect 590804 62132 590810 62144
rect 598934 62132 598940 62144
rect 590804 62104 598940 62132
rect 590804 62092 590810 62104
rect 598934 62092 598940 62104
rect 598992 62092 598998 62144
rect 595070 60800 595076 60852
rect 595128 60840 595134 60852
rect 600222 60840 600228 60852
rect 595128 60812 600228 60840
rect 595128 60800 595134 60812
rect 600222 60800 600228 60812
rect 600280 60800 600286 60852
rect 583662 60772 583668 60784
rect 579632 60744 583668 60772
rect 578234 60664 578240 60716
rect 578292 60704 578298 60716
rect 579632 60704 579660 60744
rect 583662 60732 583668 60744
rect 583720 60732 583726 60784
rect 578292 60676 579660 60704
rect 578292 60664 578298 60676
rect 579614 60460 579620 60512
rect 579672 60500 579678 60512
rect 583754 60500 583760 60512
rect 579672 60472 583760 60500
rect 579672 60460 579678 60472
rect 583754 60460 583760 60472
rect 583812 60460 583818 60512
rect 579614 58624 579620 58676
rect 579672 58664 579678 58676
rect 583846 58664 583852 58676
rect 579672 58636 583852 58664
rect 579672 58624 579678 58636
rect 583846 58624 583852 58636
rect 583904 58624 583910 58676
rect 582558 58080 582564 58132
rect 582616 58120 582622 58132
rect 591942 58120 591948 58132
rect 582616 58092 591948 58120
rect 582616 58080 582622 58092
rect 591942 58080 591948 58092
rect 592000 58080 592006 58132
rect 586422 57944 586428 57996
rect 586480 57984 586486 57996
rect 590654 57984 590660 57996
rect 586480 57956 590660 57984
rect 586480 57944 586486 57956
rect 590654 57944 590660 57956
rect 590712 57944 590718 57996
rect 590746 57944 590752 57996
rect 590804 57944 590810 57996
rect 585134 57876 585140 57928
rect 585192 57916 585198 57928
rect 590764 57916 590792 57944
rect 585192 57888 590792 57916
rect 585192 57876 585198 57888
rect 587894 55224 587900 55276
rect 587952 55264 587958 55276
rect 595070 55264 595076 55276
rect 587952 55236 595076 55264
rect 587952 55224 587958 55236
rect 595070 55224 595076 55236
rect 595128 55224 595134 55276
rect 582558 53632 582564 53644
rect 571352 53604 582564 53632
rect 571352 53576 571380 53604
rect 582558 53592 582564 53604
rect 582616 53592 582622 53644
rect 571334 53524 571340 53576
rect 571392 53524 571398 53576
rect 346854 52368 346860 52420
rect 346912 52408 346918 52420
rect 642910 52408 642916 52420
rect 346912 52380 642916 52408
rect 346912 52368 346918 52380
rect 642910 52368 642916 52380
rect 642968 52368 642974 52420
rect 52086 51008 52092 51060
rect 52144 51048 52150 51060
rect 213822 51048 213828 51060
rect 52144 51020 213828 51048
rect 52144 51008 52150 51020
rect 213822 51008 213828 51020
rect 213880 51048 213886 51060
rect 346486 51048 346492 51060
rect 213880 51020 346492 51048
rect 213880 51008 213886 51020
rect 346486 51008 346492 51020
rect 346544 51008 346550 51060
rect 587986 51008 587992 51060
rect 588044 51048 588050 51060
rect 600314 51048 600320 51060
rect 588044 51020 600320 51048
rect 588044 51008 588050 51020
rect 600314 51008 600320 51020
rect 600372 51008 600378 51060
rect 579614 49784 579620 49836
rect 579672 49824 579678 49836
rect 585134 49824 585140 49836
rect 579672 49796 585140 49824
rect 579672 49784 579678 49796
rect 585134 49784 585140 49796
rect 585192 49784 585198 49836
rect 578602 49716 578608 49768
rect 578660 49756 578666 49768
rect 587894 49756 587900 49768
rect 578660 49728 587900 49756
rect 578660 49716 578666 49728
rect 587894 49716 587900 49728
rect 587952 49716 587958 49768
rect 478138 48424 478144 48476
rect 478196 48464 478202 48476
rect 518802 48464 518808 48476
rect 478196 48436 518808 48464
rect 478196 48424 478202 48436
rect 518802 48424 518808 48436
rect 518860 48424 518866 48476
rect 149238 48356 149244 48408
rect 149296 48396 149302 48408
rect 150250 48396 150256 48408
rect 149296 48368 150256 48396
rect 149296 48356 149302 48368
rect 150250 48356 150256 48368
rect 150308 48396 150314 48408
rect 218054 48396 218060 48408
rect 150308 48368 218060 48396
rect 150308 48356 150314 48368
rect 218054 48356 218060 48368
rect 218112 48356 218118 48408
rect 412634 48356 412640 48408
rect 412692 48396 412698 48408
rect 494054 48396 494060 48408
rect 412692 48368 494060 48396
rect 412692 48356 412698 48368
rect 494054 48356 494060 48368
rect 494112 48356 494118 48408
rect 216122 48288 216128 48340
rect 216180 48328 216186 48340
rect 521838 48328 521844 48340
rect 216180 48300 521844 48328
rect 216180 48288 216186 48300
rect 521838 48288 521844 48300
rect 521896 48288 521902 48340
rect 552014 48288 552020 48340
rect 552072 48328 552078 48340
rect 575658 48328 575664 48340
rect 552072 48300 575664 48328
rect 552072 48288 552078 48300
rect 575658 48288 575664 48300
rect 575716 48288 575722 48340
rect 52270 47064 52276 47116
rect 52328 47104 52334 47116
rect 149238 47104 149244 47116
rect 52328 47076 149244 47104
rect 52328 47064 52334 47076
rect 149238 47064 149244 47076
rect 149296 47064 149302 47116
rect 574830 46928 574836 46980
rect 574888 46968 574894 46980
rect 578234 46968 578240 46980
rect 574888 46940 578240 46968
rect 574888 46928 574894 46940
rect 578234 46928 578240 46940
rect 578292 46928 578298 46980
rect 218054 46860 218060 46912
rect 218112 46900 218118 46912
rect 642634 46900 642640 46912
rect 218112 46872 642640 46900
rect 218112 46860 218118 46872
rect 642634 46860 642640 46872
rect 642692 46860 642698 46912
rect 494054 46792 494060 46844
rect 494112 46832 494118 46844
rect 502242 46832 502248 46844
rect 494112 46804 502248 46832
rect 494112 46792 494118 46804
rect 502242 46792 502248 46804
rect 502300 46792 502306 46844
rect 460658 45840 460664 45892
rect 460716 45880 460722 45892
rect 610250 45880 610256 45892
rect 460716 45852 610256 45880
rect 460716 45840 460722 45852
rect 610250 45840 610256 45852
rect 610308 45840 610314 45892
rect 367094 45772 367100 45824
rect 367152 45812 367158 45824
rect 607398 45812 607404 45824
rect 367152 45784 607404 45812
rect 367152 45772 367158 45784
rect 607398 45772 607404 45784
rect 607456 45772 607462 45824
rect 311894 45704 311900 45756
rect 311952 45744 311958 45756
rect 607582 45744 607588 45756
rect 311952 45716 607588 45744
rect 311952 45704 311958 45716
rect 607582 45704 607588 45716
rect 607640 45704 607646 45756
rect 85114 45636 85120 45688
rect 85172 45676 85178 45688
rect 475654 45676 475660 45688
rect 85172 45648 475660 45676
rect 85172 45636 85178 45648
rect 475654 45636 475660 45648
rect 475712 45636 475718 45688
rect 540882 45636 540888 45688
rect 540940 45676 540946 45688
rect 578602 45676 578608 45688
rect 540940 45648 578608 45676
rect 540940 45636 540946 45648
rect 578602 45636 578608 45648
rect 578660 45636 578666 45688
rect 233142 45568 233148 45620
rect 233200 45608 233206 45620
rect 642818 45608 642824 45620
rect 233200 45580 642824 45608
rect 233200 45568 233206 45580
rect 642818 45568 642824 45580
rect 642876 45568 642882 45620
rect 212442 45500 212448 45552
rect 212500 45540 212506 45552
rect 639322 45540 639328 45552
rect 212500 45512 639328 45540
rect 212500 45500 212506 45512
rect 639322 45500 639328 45512
rect 639380 45500 639386 45552
rect 311894 44180 311900 44192
rect 310440 44152 311900 44180
rect 310440 44124 310468 44152
rect 311894 44140 311900 44152
rect 311952 44140 311958 44192
rect 367094 44180 367100 44192
rect 365180 44152 367100 44180
rect 365180 44124 365208 44152
rect 367094 44140 367100 44152
rect 367152 44140 367158 44192
rect 563606 44140 563612 44192
rect 563664 44180 563670 44192
rect 578142 44180 578148 44192
rect 563664 44152 578148 44180
rect 563664 44140 563670 44152
rect 578142 44140 578148 44152
rect 578200 44140 578206 44192
rect 310422 44072 310428 44124
rect 310480 44072 310486 44124
rect 365162 44072 365168 44124
rect 365220 44072 365226 44124
rect 474458 44072 474464 44124
rect 474516 44112 474522 44124
rect 586422 44112 586428 44124
rect 474516 44084 586428 44112
rect 474516 44072 474522 44084
rect 586422 44072 586428 44084
rect 586480 44072 586486 44124
rect 419718 44004 419724 44056
rect 419776 44044 419782 44056
rect 540882 44044 540888 44056
rect 419776 44016 540888 44044
rect 419776 44004 419782 44016
rect 540882 44004 540888 44016
rect 540940 44004 540946 44056
rect 405550 43936 405556 43988
rect 405608 43976 405614 43988
rect 607214 43976 607220 43988
rect 405608 43948 607220 43976
rect 405608 43936 405614 43948
rect 607214 43936 607220 43948
rect 607272 43936 607278 43988
rect 230934 43868 230940 43920
rect 230992 43908 230998 43920
rect 613010 43908 613016 43920
rect 230992 43880 613016 43908
rect 230992 43868 230998 43880
rect 613010 43868 613016 43880
rect 613068 43868 613074 43920
rect 230382 43800 230388 43852
rect 230440 43840 230446 43852
rect 618254 43840 618260 43852
rect 230440 43812 618260 43840
rect 230440 43800 230446 43812
rect 618254 43800 618260 43812
rect 618312 43800 618318 43852
rect 230750 43732 230756 43784
rect 230808 43772 230814 43784
rect 621198 43772 621204 43784
rect 230808 43744 621204 43772
rect 230808 43732 230814 43744
rect 621198 43732 621204 43744
rect 621256 43732 621262 43784
rect 230842 43664 230848 43716
rect 230900 43704 230906 43716
rect 621290 43704 621296 43716
rect 230900 43676 621296 43704
rect 230900 43664 230906 43676
rect 621290 43664 621296 43676
rect 621348 43664 621354 43716
rect 230566 43596 230572 43648
rect 230624 43636 230630 43648
rect 621474 43636 621480 43648
rect 230624 43608 621480 43636
rect 230624 43596 230630 43608
rect 621474 43596 621480 43608
rect 621532 43596 621538 43648
rect 230474 43528 230480 43580
rect 230532 43568 230538 43580
rect 621106 43568 621112 43580
rect 230532 43540 621112 43568
rect 230532 43528 230538 43540
rect 621106 43528 621112 43540
rect 621164 43528 621170 43580
rect 230658 43460 230664 43512
rect 230716 43500 230722 43512
rect 621382 43500 621388 43512
rect 230716 43472 621388 43500
rect 230716 43460 230722 43472
rect 621382 43460 621388 43472
rect 621440 43460 621446 43512
rect 226242 43392 226248 43444
rect 226300 43432 226306 43444
rect 622486 43432 622492 43444
rect 226300 43404 622492 43432
rect 226300 43392 226306 43404
rect 622486 43392 622492 43404
rect 622544 43392 622550 43444
rect 223482 43324 223488 43376
rect 223540 43364 223546 43376
rect 622302 43364 622308 43376
rect 223540 43336 622308 43364
rect 223540 43324 223546 43336
rect 622302 43324 622308 43336
rect 622360 43324 622366 43376
rect 209682 43256 209688 43308
rect 209740 43296 209746 43308
rect 631870 43296 631876 43308
rect 209740 43268 631876 43296
rect 209740 43256 209746 43268
rect 631870 43256 631876 43268
rect 631928 43256 631934 43308
rect 52178 42848 52184 42900
rect 52236 42888 52242 42900
rect 215294 42888 215300 42900
rect 52236 42860 215300 42888
rect 52236 42848 52242 42860
rect 215294 42848 215300 42860
rect 215352 42848 215358 42900
rect 530670 42344 530676 42356
rect 525720 42316 530676 42344
rect 455414 42236 455420 42288
rect 455472 42276 455478 42288
rect 525720 42276 525748 42316
rect 530670 42304 530676 42316
rect 530728 42304 530734 42356
rect 531038 42304 531044 42356
rect 531096 42304 531102 42356
rect 455472 42248 525748 42276
rect 531056 42276 531084 42304
rect 574830 42276 574836 42288
rect 531056 42248 574836 42276
rect 455472 42236 455478 42248
rect 574830 42236 574836 42248
rect 574888 42236 574894 42288
rect 510614 42168 510620 42220
rect 510672 42208 510678 42220
rect 530670 42208 530676 42220
rect 510672 42180 530676 42208
rect 510672 42168 510678 42180
rect 530670 42168 530676 42180
rect 530728 42168 530734 42220
rect 531038 42168 531044 42220
rect 531096 42208 531102 42220
rect 579522 42208 579528 42220
rect 531096 42180 579528 42208
rect 531096 42168 531102 42180
rect 579522 42168 579528 42180
rect 579580 42168 579586 42220
rect 502242 41828 502248 41880
rect 502300 41868 502306 41880
rect 518526 41868 518532 41880
rect 502300 41840 518532 41868
rect 502300 41828 502306 41840
rect 518526 41828 518532 41840
rect 518584 41828 518590 41880
rect 416682 41760 416688 41812
rect 416740 41800 416746 41812
rect 420730 41800 420736 41812
rect 416740 41772 420736 41800
rect 416740 41760 416746 41772
rect 420730 41760 420736 41772
rect 420788 41760 420794 41812
rect 471698 41760 471704 41812
rect 471756 41800 471762 41812
rect 475562 41800 475568 41812
rect 471756 41772 475568 41800
rect 471756 41760 471762 41772
rect 475562 41760 475568 41772
rect 475620 41760 475626 41812
rect 514018 41760 514024 41812
rect 514076 41800 514082 41812
rect 514846 41800 514852 41812
rect 514076 41772 514852 41800
rect 514076 41760 514082 41772
rect 514846 41760 514852 41772
rect 514904 41760 514910 41812
rect 529658 41760 529664 41812
rect 529716 41800 529722 41812
rect 530210 41800 530216 41812
rect 529716 41772 530216 41800
rect 529716 41760 529722 41772
rect 530210 41760 530216 41772
rect 530268 41760 530274 41812
rect 141786 41488 141792 41540
rect 141844 41528 141850 41540
rect 207014 41528 207020 41540
rect 141844 41500 207020 41528
rect 141844 41488 141850 41500
rect 207014 41488 207020 41500
rect 207072 41528 207078 41540
rect 209682 41528 209688 41540
rect 207072 41500 209688 41528
rect 207072 41488 207078 41500
rect 209682 41488 209688 41500
rect 209740 41488 209746 41540
rect 505646 38632 505652 38684
rect 505704 38672 505710 38684
rect 510614 38672 510620 38684
rect 505704 38644 510620 38672
rect 505704 38632 505710 38644
rect 510614 38632 510620 38644
rect 510672 38632 510678 38684
rect 420730 38564 420736 38616
rect 420788 38604 420794 38616
rect 455414 38604 455420 38616
rect 420788 38576 455420 38604
rect 420788 38564 420794 38576
rect 455414 38564 455420 38576
rect 455472 38564 455478 38616
rect 475654 38564 475660 38616
rect 475712 38604 475718 38616
rect 514018 38604 514024 38616
rect 475712 38576 514024 38604
rect 475712 38564 475718 38576
rect 514018 38564 514024 38576
rect 514076 38564 514082 38616
rect 475562 38496 475568 38548
rect 475620 38536 475626 38548
rect 505646 38536 505652 38548
rect 475620 38508 505652 38536
rect 475620 38496 475626 38508
rect 505646 38496 505652 38508
rect 505704 38496 505710 38548
rect 213178 24760 213184 24812
rect 213236 24800 213242 24812
rect 213822 24800 213828 24812
rect 213236 24772 213828 24800
rect 213236 24760 213242 24772
rect 213822 24760 213828 24772
rect 213880 24760 213886 24812
rect 224586 22992 224592 23044
rect 224644 23032 224650 23044
rect 226242 23032 226248 23044
rect 224644 23004 226248 23032
rect 224644 22992 224650 23004
rect 226242 22992 226248 23004
rect 226300 22992 226306 23044
rect 221734 22516 221740 22568
rect 221792 22556 221798 22568
rect 223482 22556 223488 22568
rect 221792 22528 223488 22556
rect 221792 22516 221798 22528
rect 223482 22516 223488 22528
rect 223540 22516 223546 22568
rect 229370 6468 229376 6520
rect 229428 6508 229434 6520
rect 233142 6508 233148 6520
rect 229428 6480 233148 6508
rect 229428 6468 229434 6480
rect 233142 6468 233148 6480
rect 233200 6468 233206 6520
<< via1 >>
rect 145196 1007428 145248 1007480
rect 154580 1007428 154632 1007480
rect 501328 1007360 501380 1007412
rect 517336 1007360 517388 1007412
rect 424692 1006000 424744 1006052
rect 466460 1006000 466512 1006052
rect 423864 1005864 423916 1005916
rect 440148 1005864 440200 1005916
rect 424324 1005796 424376 1005848
rect 440424 1005796 440476 1005848
rect 503352 1005796 503404 1005848
rect 520188 1005796 520240 1005848
rect 502984 1005728 503036 1005780
rect 520004 1005728 520056 1005780
rect 356060 1005660 356112 1005712
rect 374276 1005660 374328 1005712
rect 502524 1005660 502576 1005712
rect 519176 1005660 519228 1005712
rect 356520 1005592 356572 1005644
rect 377312 1005592 377364 1005644
rect 504548 1005592 504600 1005644
rect 517244 1005592 517296 1005644
rect 200028 1005524 200080 1005576
rect 207204 1005524 207256 1005576
rect 505836 1005524 505888 1005576
rect 517612 1005524 517664 1005576
rect 144828 1005456 144880 1005508
rect 160284 1005456 160336 1005508
rect 195336 1005456 195388 1005508
rect 209596 1005456 209648 1005508
rect 361028 1005456 361080 1005508
rect 377956 1005456 378008 1005508
rect 505376 1005456 505428 1005508
rect 517428 1005456 517480 1005508
rect 145104 1005388 145156 1005440
rect 154948 1005388 155000 1005440
rect 92500 1005320 92552 1005372
rect 109316 1005320 109368 1005372
rect 145012 1005320 145064 1005372
rect 153752 1005320 153804 1005372
rect 360200 1005320 360252 1005372
rect 380808 1005320 380860 1005372
rect 423496 1005320 423548 1005372
rect 467840 1005320 467892 1005372
rect 144920 1005252 144972 1005304
rect 153292 1005252 153344 1005304
rect 259828 1005252 259880 1005304
rect 280344 1005252 280396 1005304
rect 428372 1005252 428424 1005304
rect 453948 1005252 454000 1005304
rect 148876 1005184 148928 1005236
rect 151268 1005184 151320 1005236
rect 260196 1005184 260248 1005236
rect 265256 1005184 265308 1005236
rect 359740 1005184 359792 1005236
rect 370412 1005184 370464 1005236
rect 106464 1005116 106516 1005168
rect 125600 1005116 125652 1005168
rect 201868 1005116 201920 1005168
rect 227628 1005116 227680 1005168
rect 261852 1005116 261904 1005168
rect 149704 1005048 149756 1005100
rect 150440 1005048 150492 1005100
rect 175188 1005048 175240 1005100
rect 208400 1005048 208452 1005100
rect 227812 1005048 227864 1005100
rect 263048 1005048 263100 1005100
rect 265536 1005048 265588 1005100
rect 504180 1005116 504232 1005168
rect 520372 1005116 520424 1005168
rect 270468 1005048 270520 1005100
rect 358176 1005048 358228 1005100
rect 366732 1005048 366784 1005100
rect 428832 1005048 428884 1005100
rect 464252 1005048 464304 1005100
rect 551928 1005048 551980 1005100
rect 568580 1005048 568632 1005100
rect 148876 1004980 148928 1005032
rect 150900 1004980 150952 1005032
rect 148140 1004912 148192 1004964
rect 154120 1004912 154172 1004964
rect 159456 1004912 159508 1004964
rect 173900 1004912 173952 1004964
rect 204168 1004912 204220 1004964
rect 211620 1004980 211672 1005032
rect 260656 1004980 260708 1005032
rect 209228 1004912 209280 1004964
rect 227720 1004912 227772 1004964
rect 262680 1004912 262732 1004964
rect 265536 1004912 265588 1004964
rect 356888 1004980 356940 1005032
rect 378048 1004980 378100 1005032
rect 425520 1004980 425572 1005032
rect 455604 1004980 455656 1005032
rect 280160 1004912 280212 1004964
rect 358544 1004912 358596 1004964
rect 383098 1004912 383150 1004964
rect 426808 1004912 426860 1004964
rect 455512 1004912 455564 1004964
rect 505008 1004912 505060 1004964
rect 522948 1004912 523000 1004964
rect 551652 1004912 551704 1004964
rect 554780 1004912 554832 1004964
rect 108028 1004844 108080 1004896
rect 92960 1004708 93012 1004760
rect 108856 1004776 108908 1004828
rect 148876 1004844 148928 1004896
rect 152096 1004844 152148 1004896
rect 210884 1004844 210936 1004896
rect 125692 1004776 125744 1004828
rect 148784 1004776 148836 1004828
rect 152924 1004776 152976 1004828
rect 156972 1004776 157024 1004828
rect 174084 1004776 174136 1004828
rect 195704 1004776 195756 1004828
rect 206376 1004776 206428 1004828
rect 261024 1004844 261076 1004896
rect 265072 1004844 265124 1004896
rect 357348 1004844 357400 1004896
rect 362500 1004844 362552 1004896
rect 427176 1004844 427228 1004896
rect 455420 1004844 455472 1004896
rect 553124 1004844 553176 1004896
rect 555516 1004844 555568 1004896
rect 227904 1004776 227956 1004828
rect 262220 1004776 262272 1004828
rect 280252 1004776 280304 1004828
rect 357716 1004776 357768 1004828
rect 364248 1004776 364300 1004828
rect 427544 1004776 427596 1004828
rect 466552 1004776 466604 1004828
rect 500500 1004776 500552 1004828
rect 509332 1004776 509384 1004828
rect 553952 1004776 554004 1004828
rect 555700 1004776 555752 1004828
rect 105636 1004708 105688 1004760
rect 125784 1004708 125836 1004760
rect 148876 1004708 148928 1004760
rect 151728 1004708 151780 1004760
rect 157800 1004708 157852 1004760
rect 173992 1004708 174044 1004760
rect 201040 1004708 201092 1004760
rect 201868 1004708 201920 1004760
rect 261484 1004708 261536 1004760
rect 265164 1004708 265216 1004760
rect 360568 1004708 360620 1004760
rect 366364 1004708 366416 1004760
rect 419080 1004708 419132 1004760
rect 421840 1004708 421892 1004760
rect 422668 1004708 422720 1004760
rect 425152 1004708 425204 1004760
rect 467748 1004708 467800 1004760
rect 496636 1004708 496688 1004760
rect 498844 1004708 498896 1004760
rect 499672 1004708 499724 1004760
rect 501696 1004708 501748 1004760
rect 509240 1004708 509292 1004760
rect 549444 1004708 549496 1004760
rect 550272 1004708 550324 1004760
rect 551100 1004708 551152 1004760
rect 552756 1004708 552808 1004760
rect 571248 1004844 571300 1004896
rect 98276 1004640 98328 1004692
rect 99104 1004640 99156 1004692
rect 125508 1004640 125560 1004692
rect 148968 1004640 149020 1004692
rect 152556 1004640 152608 1004692
rect 154488 1004640 154540 1004692
rect 160652 1004640 160704 1004692
rect 195152 1004640 195204 1004692
rect 205916 1004640 205968 1004692
rect 252468 1004640 252520 1004692
rect 253296 1004640 253348 1004692
rect 280068 1004640 280120 1004692
rect 315120 1004640 315172 1004692
rect 331220 1004640 331272 1004692
rect 361396 1004640 361448 1004692
rect 365444 1004640 365496 1004692
rect 366732 1004640 366784 1004692
rect 383282 1004640 383334 1004692
rect 466460 1004640 466512 1004692
rect 472256 1004640 472308 1004692
rect 502156 1004640 502208 1004692
rect 509148 1004640 509200 1004692
rect 517336 1004640 517388 1004692
rect 523592 1004640 523644 1004692
rect 555700 1004164 555752 1004216
rect 569868 1004164 569920 1004216
rect 555516 1003892 555568 1003944
rect 569960 1003892 570012 1003944
rect 553492 1003484 553544 1003536
rect 556160 1003484 556212 1003536
rect 455420 1003280 455472 1003332
rect 469036 1003280 469088 1003332
rect 554688 1003280 554740 1003332
rect 571616 1003280 571668 1003332
rect 455512 1003212 455564 1003264
rect 469128 1003212 469180 1003264
rect 554320 1003212 554372 1003264
rect 571432 1003212 571484 1003264
rect 568580 1002056 568632 1002108
rect 571524 1002056 571576 1002108
rect 440148 1001988 440200 1002040
rect 440424 1001920 440476 1001972
rect 143908 1001852 143960 1001904
rect 148784 1001852 148836 1001904
rect 362500 1001852 362552 1001904
rect 364432 1001852 364484 1001904
rect 447140 1001852 447192 1001904
rect 466552 1001920 466604 1001972
rect 472624 1001920 472676 1001972
rect 519176 1001920 519228 1001972
rect 523776 1001920 523828 1001972
rect 590660 1001920 590712 1001972
rect 625804 1001920 625856 1001972
rect 447324 1001852 447376 1001904
rect 377312 1001716 377364 1001768
rect 378324 1001716 378376 1001768
rect 556160 1001240 556212 1001292
rect 571248 1001240 571300 1001292
rect 366364 1000764 366416 1000816
rect 383558 1000764 383610 1000816
rect 455604 1000696 455656 1000748
rect 472164 1000696 472216 1000748
rect 365444 1000628 365496 1000680
rect 383374 1000628 383426 1000680
rect 428004 1000628 428056 1000680
rect 472624 1000628 472676 1000680
rect 370412 1000560 370464 1000612
rect 383466 1000560 383518 1000612
rect 426348 1000560 426400 1000612
rect 472532 1000560 472584 1000612
rect 358912 1000492 358964 1000544
rect 383558 1000492 383610 1000544
rect 425980 1000492 426032 1000544
rect 472348 1000492 472400 1000544
rect 374276 1000424 374328 1000476
rect 380992 1000424 381044 1000476
rect 380900 1000356 380952 1000408
rect 383558 1000356 383610 1000408
rect 555976 1000016 556028 1000068
rect 567016 1000016 567068 1000068
rect 92408 999880 92460 999932
rect 118700 999880 118752 999932
rect 246764 999880 246816 999932
rect 258632 999880 258684 999932
rect 92592 999812 92644 999864
rect 104348 999812 104400 999864
rect 246672 999812 246724 999864
rect 257344 999812 257396 999864
rect 312176 999812 312228 999864
rect 318892 999812 318944 999864
rect 430856 999812 430908 999864
rect 439824 999812 439876 999864
rect 93052 999744 93104 999796
rect 102784 999744 102836 999796
rect 246580 999744 246632 999796
rect 256976 999744 257028 999796
rect 310152 999744 310204 999796
rect 314936 999744 314988 999796
rect 431684 999744 431736 999796
rect 437940 999744 437992 999796
rect 508688 999744 508740 999796
rect 515220 999744 515272 999796
rect 92316 999676 92368 999728
rect 100668 999676 100720 999728
rect 195428 999676 195480 999728
rect 205548 999676 205600 999728
rect 246856 999676 246908 999728
rect 257804 999676 257856 999728
rect 311440 999676 311492 999728
rect 315948 999676 316000 999728
rect 361856 999676 361908 999728
rect 368756 999676 368808 999728
rect 429200 999676 429252 999728
rect 434628 999676 434680 999728
rect 506204 999676 506256 999728
rect 512092 999676 512144 999728
rect 92868 999608 92920 999660
rect 102324 999608 102376 999660
rect 195520 999608 195572 999660
rect 203892 999608 203944 999660
rect 249708 999608 249760 999660
rect 254860 999608 254912 999660
rect 313832 999608 313884 999660
rect 318708 999608 318760 999660
rect 362592 999608 362644 999660
rect 368572 999608 368624 999660
rect 430028 999608 430080 999660
rect 434812 999608 434864 999660
rect 508228 999608 508280 999660
rect 513472 999608 513524 999660
rect 92776 999540 92828 999592
rect 101956 999540 102008 999592
rect 155776 999540 155828 999592
rect 160284 999540 160336 999592
rect 195612 999540 195664 999592
rect 203524 999540 203576 999592
rect 250444 999540 250496 999592
rect 256148 999540 256200 999592
rect 312636 999540 312688 999592
rect 315120 999540 315172 999592
rect 363420 999540 363472 999592
rect 368940 999540 368992 999592
rect 431224 999540 431276 999592
rect 436192 999540 436244 999592
rect 507032 999540 507084 999592
rect 511908 999540 511960 999592
rect 95148 999472 95200 999524
rect 101496 999472 101548 999524
rect 159088 999472 159140 999524
rect 162860 999472 162912 999524
rect 198464 999472 198516 999524
rect 204352 999472 204404 999524
rect 250260 999472 250312 999524
rect 255688 999472 255740 999524
rect 314844 999472 314896 999524
rect 319076 999472 319128 999524
rect 365076 999472 365128 999524
rect 371516 999472 371568 999524
rect 432420 999472 432472 999524
rect 437572 999472 437624 999524
rect 507860 999472 507912 999524
rect 512276 999472 512328 999524
rect 97908 999404 97960 999456
rect 103152 999404 103204 999456
rect 198372 999404 198424 999456
rect 204720 999404 204772 999456
rect 208860 999404 208912 999456
rect 212724 999404 212776 999456
rect 250076 999404 250128 999456
rect 255320 999404 255372 999456
rect 362224 999404 362276 999456
rect 367192 999404 367244 999456
rect 432880 999404 432932 999456
rect 437756 999404 437808 999456
rect 506664 999404 506716 999456
rect 510712 999404 510764 999456
rect 92684 999336 92736 999388
rect 99472 999336 99524 999388
rect 195244 999336 195296 999388
rect 202236 999336 202288 999388
rect 210424 999336 210476 999388
rect 218972 999336 219024 999388
rect 246948 999336 247000 999388
rect 253664 999336 253716 999388
rect 364708 999336 364760 999388
rect 369860 999336 369912 999388
rect 429660 999336 429712 999388
rect 433340 999336 433392 999388
rect 509056 999336 509108 999388
rect 513380 999336 513432 999388
rect 95700 999268 95752 999320
rect 101128 999268 101180 999320
rect 200120 999268 200172 999320
rect 205180 999268 205232 999320
rect 209596 999268 209648 999320
rect 212632 999268 212684 999320
rect 249892 999268 249944 999320
rect 254492 999268 254544 999320
rect 365444 999268 365496 999320
rect 371148 999268 371200 999320
rect 430396 999268 430448 999320
rect 433432 999268 433484 999320
rect 507400 999268 507452 999320
rect 510620 999268 510672 999320
rect 540336 999268 540388 999320
rect 564256 999948 564308 1000000
rect 558460 999880 558512 999932
rect 564532 999880 564584 999932
rect 560852 999812 560904 999864
rect 567292 999812 567344 999864
rect 556344 999744 556396 999796
rect 562140 999744 562192 999796
rect 560484 999676 560536 999728
rect 565820 999676 565872 999728
rect 559196 999608 559248 999660
rect 564348 999608 564400 999660
rect 560024 999540 560076 999592
rect 564716 999540 564768 999592
rect 558000 999472 558052 999524
rect 563060 999472 563112 999524
rect 556804 999404 556856 999456
rect 561772 999404 561824 999456
rect 590752 999404 590804 999456
rect 625436 999404 625488 999456
rect 557172 999336 557224 999388
rect 561956 999336 562008 999388
rect 558828 999268 558880 999320
rect 563152 999268 563204 999320
rect 607128 999268 607180 999320
rect 625620 999268 625672 999320
rect 95332 999200 95384 999252
rect 100300 999200 100352 999252
rect 198648 999200 198700 999252
rect 202696 999200 202748 999252
rect 211712 999200 211764 999252
rect 216588 999200 216640 999252
rect 252468 999200 252520 999252
rect 256516 999200 256568 999252
rect 364248 999200 364300 999252
rect 368388 999200 368440 999252
rect 432052 999200 432104 999252
rect 436100 999200 436152 999252
rect 500868 999200 500920 999252
rect 507860 999200 507912 999252
rect 509516 999200 509568 999252
rect 514668 999200 514720 999252
rect 548892 999200 548944 999252
rect 554320 999200 554372 999252
rect 559656 999200 559708 999252
rect 563244 999200 563296 999252
rect 602252 999200 602304 999252
rect 625712 999200 625764 999252
rect 92316 999132 92368 999184
rect 93052 999132 93104 999184
rect 95516 999132 95568 999184
rect 99932 999132 99984 999184
rect 143816 999132 143868 999184
rect 148968 999132 149020 999184
rect 154120 999132 154172 999184
rect 155776 999132 155828 999184
rect 198556 999132 198608 999184
rect 203064 999132 203116 999184
rect 211252 999132 211304 999184
rect 215300 999132 215352 999184
rect 250628 999132 250680 999184
rect 254124 999132 254176 999184
rect 258540 999132 258592 999184
rect 262220 999132 262272 999184
rect 355968 999132 356020 999184
rect 358912 999132 358964 999184
rect 363052 999132 363104 999184
rect 367100 999132 367152 999184
rect 378048 999132 378100 999184
rect 383190 999132 383242 999184
rect 400036 999132 400088 999184
rect 444380 999132 444432 999184
rect 464252 999132 464304 999184
rect 472440 999132 472492 999184
rect 499488 999132 499540 999184
rect 503352 999132 503404 999184
rect 509884 999132 509936 999184
rect 514852 999132 514904 999184
rect 549076 999132 549128 999184
rect 551928 999132 551980 999184
rect 557632 999132 557684 999184
rect 561588 999132 561640 999184
rect 561680 999132 561732 999184
rect 567108 999132 567160 999184
rect 612740 999132 612792 999184
rect 625804 999132 625856 999184
rect 118700 999064 118752 999116
rect 122104 999064 122156 999116
rect 144000 999064 144052 999116
rect 158260 999064 158312 999116
rect 247960 999064 248012 999116
rect 265164 999064 265216 999116
rect 298744 999064 298796 999116
rect 312636 999064 312688 999116
rect 399944 999064 399996 999116
rect 436192 999064 436244 999116
rect 453948 999064 454000 999116
rect 462780 999064 462832 999116
rect 488908 999064 488960 999116
rect 513472 999064 513524 999116
rect 509332 998996 509384 999048
rect 521292 998996 521344 999048
rect 509240 998928 509292 998980
rect 521476 998928 521528 998980
rect 509148 998860 509200 998912
rect 521384 998860 521436 998912
rect 507860 998792 507912 998844
rect 521568 998792 521620 998844
rect 467748 998316 467800 998368
rect 470876 998316 470928 998368
rect 364340 998180 364392 998232
rect 375196 998180 375248 998232
rect 467840 998112 467892 998164
rect 469404 998112 469456 998164
rect 364432 997908 364484 997960
rect 374460 997908 374512 997960
rect 549076 997772 549128 997824
rect 575572 997772 575624 997824
rect 144092 997704 144144 997756
rect 156144 997704 156196 997756
rect 571524 997704 571576 997756
rect 623780 997704 623832 997756
rect 561956 997636 562008 997688
rect 590660 997636 590712 997688
rect 548892 997568 548944 997620
rect 612740 997568 612792 997620
rect 571340 997500 571392 997552
rect 590752 997500 590804 997552
rect 569868 997432 569920 997484
rect 607128 997432 607180 997484
rect 571432 997364 571484 997416
rect 602252 997364 602304 997416
rect 562140 997296 562192 997348
rect 623688 997296 623740 997348
rect 107660 997160 107712 997212
rect 115940 997160 115992 997212
rect 144000 997092 144052 997144
rect 147772 997092 147824 997144
rect 301780 996276 301832 996328
rect 308128 996276 308180 996328
rect 300216 996208 300268 996260
rect 305736 996208 305788 996260
rect 125600 996135 125652 996187
rect 157800 996135 157852 996187
rect 173900 996135 173952 996187
rect 215300 996135 215352 996187
rect 227904 996135 227956 996187
rect 267832 996135 267884 996187
rect 270408 996135 270460 996187
rect 280252 996130 280304 996182
rect 314292 996140 314344 996192
rect 512276 996130 512328 996182
rect 563244 996130 563296 996182
rect 108488 996072 108540 996124
rect 113364 996072 113416 996124
rect 125692 996067 125744 996119
rect 159456 996067 159508 996119
rect 173992 996067 174044 996119
rect 212632 996067 212684 996119
rect 227812 996067 227864 996119
rect 265256 996067 265308 996119
rect 267648 996067 267700 996119
rect 280160 996062 280212 996114
rect 315120 996072 315172 996124
rect 317512 996072 317564 996124
rect 125784 995999 125836 996051
rect 156972 995999 157024 996051
rect 160468 995999 160520 996051
rect 174084 995999 174136 996051
rect 212724 995999 212776 996051
rect 227720 995999 227772 996051
rect 265072 995999 265124 996051
rect 267556 995999 267608 996051
rect 280344 995994 280396 996046
rect 311808 995994 311860 996046
rect 92684 995936 92736 995988
rect 86592 995800 86644 995852
rect 88984 995800 89036 995852
rect 92408 995868 92460 995920
rect 86040 995732 86092 995784
rect 92234 995800 92286 995852
rect 136272 995800 136324 995852
rect 145196 995931 145248 995983
rect 143724 995862 143776 995914
rect 136824 995800 136876 995852
rect 137928 995800 137980 995852
rect 143632 995800 143684 995852
rect 91560 995732 91612 995784
rect 92326 995732 92378 995784
rect 139216 995732 139268 995784
rect 143816 995732 143868 995784
rect 183284 995732 183336 995784
rect 195704 995931 195756 995983
rect 195612 995863 195664 995915
rect 246948 995868 247000 995920
rect 307760 995926 307812 995978
rect 383466 995936 383518 995988
rect 188804 995786 188856 995838
rect 189448 995790 189500 995842
rect 195244 995795 195296 995847
rect 240876 995800 240928 995852
rect 245568 995800 245620 995852
rect 246488 995800 246540 995852
rect 286784 995800 286836 995852
rect 306932 995858 306984 995910
rect 383374 995868 383426 995920
rect 472164 995936 472216 995988
rect 472716 995868 472768 995920
rect 293592 995790 293644 995842
rect 295064 995790 295116 995842
rect 310152 995800 310204 995852
rect 383742 995800 383794 995852
rect 384396 995800 384448 995852
rect 385684 995800 385736 995852
rect 391940 995800 391992 995852
rect 396632 995800 396684 995852
rect 400036 995800 400088 995852
rect 472532 995800 472584 995852
rect 474004 995800 474056 995852
rect 476396 995800 476448 995852
rect 625620 995936 625672 995988
rect 523592 995868 523644 995920
rect 625896 995868 625948 995920
rect 477684 995800 477736 995852
rect 522948 995800 523000 995852
rect 524788 995800 524840 995852
rect 530124 995800 530176 995852
rect 537024 995800 537076 995852
rect 540336 995800 540388 995852
rect 623688 995800 623740 995852
rect 626540 995800 626592 995852
rect 627828 995800 627880 995852
rect 630864 995800 630916 995852
rect 194324 995732 194376 995784
rect 195428 995732 195480 995784
rect 239036 995732 239088 995784
rect 246672 995732 246724 995784
rect 383650 995732 383702 995784
rect 384948 995732 385000 995784
rect 472624 995732 472676 995784
rect 473268 995732 473320 995784
rect 523776 995732 523828 995784
rect 529020 995732 529072 995784
rect 625804 995732 625856 995784
rect 627184 995732 627236 995784
rect 89720 995664 89772 995716
rect 92592 995664 92644 995716
rect 141056 995664 141108 995716
rect 154120 995664 154172 995716
rect 188160 995664 188212 995716
rect 198648 995664 198700 995716
rect 243912 995664 243964 995716
rect 246764 995664 246816 995716
rect 291752 995664 291804 995716
rect 306472 995664 306524 995716
rect 383282 995664 383334 995716
rect 388628 995664 388680 995716
rect 472440 995664 472492 995716
rect 474740 995664 474792 995716
rect 521568 995664 521620 995716
rect 532700 995664 532752 995716
rect 625712 995664 625764 995716
rect 630220 995664 630272 995716
rect 77944 995596 77996 995648
rect 92868 995596 92920 995648
rect 133144 995596 133196 995648
rect 143908 995596 143960 995648
rect 184664 995596 184716 995648
rect 198556 995596 198608 995648
rect 239588 995596 239640 995648
rect 250628 995596 250680 995648
rect 287520 995596 287572 995648
rect 307300 995596 307352 995648
rect 383558 995596 383610 995648
rect 387524 995596 387576 995648
rect 472256 995596 472308 995648
rect 481916 995596 481968 995648
rect 521476 995596 521528 995648
rect 533436 995596 533488 995648
rect 625436 995596 625488 995648
rect 631508 995596 631560 995648
rect 132408 995528 132460 995580
rect 144920 995528 144972 995580
rect 190644 995528 190696 995580
rect 195520 995528 195572 995580
rect 383190 995528 383242 995580
rect 389364 995528 389416 995580
rect 472348 995528 472400 995580
rect 476948 995528 477000 995580
rect 130016 995460 130068 995512
rect 144092 995460 144144 995512
rect 184480 995460 184532 995512
rect 198464 995460 198516 995512
rect 380992 995460 381044 995512
rect 393596 995460 393648 995512
rect 131856 995392 131908 995444
rect 145104 995392 145156 995444
rect 183836 995392 183888 995444
rect 198372 995392 198424 995444
rect 469404 995392 469456 995444
rect 482652 995528 482704 995580
rect 521292 995528 521344 995580
rect 533988 995528 534040 995580
rect 623780 995528 623832 995580
rect 635832 995528 635884 995580
rect 469220 995324 469272 995376
rect 480812 995324 480864 995376
rect 303528 994720 303580 994772
rect 283472 993828 283524 993880
rect 301780 993828 301832 993880
rect 378324 993828 378376 993880
rect 392676 993828 392728 993880
rect 129096 993692 129148 993744
rect 145012 993760 145064 993812
rect 180156 993760 180208 993812
rect 200028 993760 200080 993812
rect 285956 993760 286008 993812
rect 309324 993760 309376 993812
rect 469312 993760 469364 993812
rect 487804 993760 487856 993812
rect 521384 993760 521436 993812
rect 535552 993760 535604 993812
rect 140504 993692 140556 993744
rect 151820 993692 151872 993744
rect 180800 993692 180852 993744
rect 200120 993692 200172 993744
rect 282828 993692 282880 993744
rect 314936 993692 314988 993744
rect 374460 993692 374512 993744
rect 393320 993692 393372 993744
rect 470876 993692 470928 993744
rect 484124 993692 484176 993744
rect 571616 993692 571668 993744
rect 633992 993692 634044 993744
rect 77024 993624 77076 993676
rect 104164 993624 104216 993676
rect 128452 993624 128504 993676
rect 160284 993624 160336 993676
rect 181444 993624 181496 993676
rect 207572 993624 207624 993676
rect 231584 993624 231636 993676
rect 262220 993624 262272 993676
rect 284116 993624 284168 993676
rect 310612 993624 310664 993676
rect 355968 993624 356020 993676
rect 398840 993624 398892 993676
rect 462780 993624 462832 993676
rect 485964 993624 486016 993676
rect 499488 993624 499540 993676
rect 539232 993624 539284 993676
rect 551652 993624 551704 993676
rect 640708 993624 640760 993676
rect 433524 993556 433576 993608
rect 434628 993556 434680 993608
rect 510712 993556 510764 993608
rect 510896 993556 510948 993608
rect 511908 993556 511960 993608
rect 563152 993556 563204 993608
rect 368572 993488 368624 993540
rect 433432 993488 433484 993540
rect 433616 993488 433668 993540
rect 434812 993488 434864 993540
rect 510620 993488 510672 993540
rect 510804 993488 510856 993540
rect 512092 993488 512144 993540
rect 563060 993488 563112 993540
rect 368756 993420 368808 993472
rect 433340 993420 433392 993472
rect 436192 993420 436244 993472
rect 437940 993420 437992 993472
rect 513380 993420 513432 993472
rect 513472 993420 513524 993472
rect 515220 993420 515272 993472
rect 565820 993420 565872 993472
rect 368388 993352 368440 993404
rect 436100 993352 436152 993404
rect 89628 990768 89680 990820
rect 92500 990768 92552 990820
rect 564256 990768 564308 990820
rect 576308 990768 576360 990820
rect 168380 990632 168432 990684
rect 170404 990632 170456 990684
rect 203156 990632 203208 990684
rect 204168 990632 204220 990684
rect 331220 990632 331272 990684
rect 332692 990632 332744 990684
rect 444380 990632 444432 990684
rect 446220 990632 446272 990684
rect 366180 989680 366232 989732
rect 381636 989680 381688 989732
rect 371148 989612 371200 989664
rect 397828 989612 397880 989664
rect 437756 989612 437808 989664
rect 462780 989612 462832 989664
rect 514852 989612 514904 989664
rect 527640 989612 527692 989664
rect 567108 989612 567160 989664
rect 592500 989612 592552 989664
rect 321468 989544 321520 989596
rect 349160 989544 349212 989596
rect 371332 989544 371384 989596
rect 414112 989544 414164 989596
rect 437388 989544 437440 989596
rect 478972 989544 479024 989596
rect 515036 989544 515088 989596
rect 543832 989544 543884 989596
rect 567476 989544 567528 989596
rect 608784 989544 608836 989596
rect 269212 989476 269264 989528
rect 300492 989476 300544 989528
rect 319076 989476 319128 989528
rect 365444 989476 365496 989528
rect 371516 989476 371568 989528
rect 430304 989476 430356 989528
rect 437572 989476 437624 989528
rect 495164 989476 495216 989528
rect 514668 989476 514720 989528
rect 560116 989476 560168 989528
rect 567292 989476 567344 989528
rect 624976 989476 625028 989528
rect 73436 989408 73488 989460
rect 92960 989408 93012 989460
rect 105820 989408 105872 989460
rect 113272 989408 113324 989460
rect 151820 989408 151872 989460
rect 186964 989408 187016 989460
rect 216588 989408 216640 989460
rect 235632 989408 235684 989460
rect 269028 989408 269080 989460
rect 284300 989408 284352 989460
rect 303528 989408 303580 989460
rect 666560 989408 666612 989460
rect 138296 988728 138348 988780
rect 144828 988728 144880 988780
rect 248328 988116 248380 988168
rect 251824 988116 251876 988168
rect 45468 988048 45520 988100
rect 367192 988048 367244 988100
rect 45744 987980 45796 988032
rect 368756 987980 368808 988032
rect 45560 987912 45612 987964
rect 369860 987912 369912 987964
rect 314292 987844 314344 987896
rect 666836 987844 666888 987896
rect 318892 987776 318944 987828
rect 669228 987776 669280 987828
rect 311808 987708 311860 987760
rect 666652 987708 666704 987760
rect 318708 987640 318760 987692
rect 669320 987640 669372 987692
rect 280068 987572 280120 987624
rect 651380 987572 651432 987624
rect 270408 987504 270460 987556
rect 652852 987504 652904 987556
rect 267648 987436 267700 987488
rect 652668 987436 652720 987488
rect 48228 987368 48280 987420
rect 433524 987368 433576 987420
rect 267556 987300 267608 987352
rect 652760 987300 652812 987352
rect 227628 987232 227680 987284
rect 651472 987232 651524 987284
rect 212632 987164 212684 987216
rect 652944 987164 652996 987216
rect 215300 987096 215352 987148
rect 658280 987096 658332 987148
rect 212724 987028 212776 987080
rect 658188 987028 658240 987080
rect 175188 986960 175240 987012
rect 651564 986960 651616 987012
rect 125508 986892 125560 986944
rect 651656 986892 651708 986944
rect 62672 986824 62724 986876
rect 113364 986824 113416 986876
rect 669596 986824 669648 986876
rect 62488 986756 62540 986808
rect 110512 986756 110564 986808
rect 669412 986756 669464 986808
rect 62304 986688 62356 986740
rect 110604 986688 110656 986740
rect 669504 986688 669556 986740
rect 564532 985464 564584 985516
rect 564716 985464 564768 985516
rect 675668 985464 675720 985516
rect 62856 985396 62908 985448
rect 669688 985396 669740 985448
rect 62396 985328 62448 985380
rect 670056 985328 670108 985380
rect 350448 985056 350500 985108
rect 670976 985056 671028 985108
rect 45652 984988 45704 985040
rect 367100 984988 367152 985040
rect 45928 984920 45980 984972
rect 368572 984920 368624 984972
rect 45836 984852 45888 984904
rect 368388 984852 368440 984904
rect 419080 984852 419132 984904
rect 670884 984852 670936 984904
rect 317512 984784 317564 984836
rect 666744 984784 666796 984836
rect 315948 984716 316000 984768
rect 671988 984716 672040 984768
rect 300768 984648 300820 984700
rect 671068 984648 671120 984700
rect 46112 984580 46164 984632
rect 433616 984580 433668 984632
rect 48320 984512 48372 984564
rect 436192 984512 436244 984564
rect 496636 984512 496688 984564
rect 670792 984512 670844 984564
rect 46388 984444 46440 984496
rect 510804 984444 510856 984496
rect 46204 984376 46256 984428
rect 510896 984376 510948 984428
rect 48412 984308 48464 984360
rect 513472 984308 513524 984360
rect 546408 984308 546460 984360
rect 670700 984308 670752 984360
rect 162860 984240 162912 984292
rect 655428 984240 655480 984292
rect 162952 984172 163004 984224
rect 658464 984172 658516 984224
rect 46020 984104 46072 984156
rect 110420 984104 110472 984156
rect 160468 984104 160520 984156
rect 658372 984104 658424 984156
rect 62212 984036 62264 984088
rect 561036 984036 561088 984088
rect 564348 984036 564400 984088
rect 649908 984036 649960 984088
rect 62120 983968 62172 984020
rect 564532 983968 564584 984020
rect 62028 983900 62080 983952
rect 564440 983900 564492 983952
rect 62580 983084 62632 983136
rect 668952 983084 669004 983136
rect 62764 983016 62816 983068
rect 670240 983016 670292 983068
rect 63132 982948 63184 983000
rect 668584 982948 668636 983000
rect 62948 982880 63000 982932
rect 668492 982880 668544 982932
rect 42340 972884 42392 972936
rect 58440 972884 58492 972936
rect 674840 970096 674892 970148
rect 675668 970096 675720 970148
rect 42156 967240 42208 967292
rect 42340 967240 42392 967292
rect 42064 967036 42116 967088
rect 42800 967036 42852 967088
rect 673552 966356 673604 966408
rect 675392 966356 675444 966408
rect 674748 965540 674800 965592
rect 675392 965540 675444 965592
rect 673460 964996 673512 965048
rect 675484 964996 675536 965048
rect 42156 963976 42208 964028
rect 42984 963976 43036 964028
rect 673644 963296 673696 963348
rect 675392 963296 675444 963348
rect 673920 962684 673972 962736
rect 675484 962684 675536 962736
rect 42156 962616 42208 962668
rect 42892 962616 42944 962668
rect 42156 962072 42208 962124
rect 43076 962072 43128 962124
rect 673828 962004 673880 962056
rect 675392 962004 675444 962056
rect 673736 961324 673788 961376
rect 675392 961324 675444 961376
rect 48504 960508 48556 960560
rect 57980 960508 58032 960560
rect 655612 960508 655664 960560
rect 675024 960508 675076 960560
rect 42892 959624 42944 959676
rect 43628 959624 43680 959676
rect 42064 959488 42116 959540
rect 42892 959488 42944 959540
rect 42156 958876 42208 958928
rect 43260 958876 43312 958928
rect 674472 958808 674524 958860
rect 675392 958808 675444 958860
rect 42064 958468 42116 958520
rect 43352 958468 43404 958520
rect 674288 958332 674340 958384
rect 675392 958332 675444 958384
rect 42064 957720 42116 957772
rect 43168 957720 43220 957772
rect 674380 957720 674432 957772
rect 675484 957720 675536 957772
rect 674564 956972 674616 957024
rect 675392 956972 675444 957024
rect 674656 955680 674708 955732
rect 675484 955680 675536 955732
rect 675024 955476 675076 955528
rect 675484 955476 675536 955528
rect 42156 955340 42208 955392
rect 42708 955340 42760 955392
rect 673920 953980 673972 954032
rect 674748 953980 674800 954032
rect 674748 953844 674800 953896
rect 675392 953844 675444 953896
rect 674840 952144 674892 952196
rect 674840 952008 674892 952060
rect 675392 952008 675444 952060
rect 675668 951736 675720 951788
rect 673920 951056 673972 951108
rect 675760 951056 675812 951108
rect 41972 950784 42024 950836
rect 62672 950784 62724 950836
rect 673460 950580 673512 950632
rect 673644 950580 673696 950632
rect 35624 949560 35676 949612
rect 43628 949560 43680 949612
rect 35716 949492 35768 949544
rect 42892 949492 42944 949544
rect 41512 949424 41564 949476
rect 58440 949424 58492 949476
rect 41788 943032 41840 943084
rect 49700 943032 49752 943084
rect 41788 942692 41840 942744
rect 48504 942692 48556 942744
rect 41788 941468 41840 941520
rect 46020 941468 46072 941520
rect 41788 941332 41840 941384
rect 42708 941332 42760 941384
rect 41880 941196 41932 941248
rect 42708 941196 42760 941248
rect 655796 938816 655848 938868
rect 676220 938816 676272 938868
rect 655704 938680 655756 938732
rect 676312 938680 676364 938732
rect 655520 938544 655572 938596
rect 676128 938544 676180 938596
rect 49700 938340 49752 938392
rect 58440 938340 58492 938392
rect 41154 936504 41206 936556
rect 41696 936504 41748 936556
rect 670332 935756 670384 935808
rect 676220 935756 676272 935808
rect 670148 935688 670200 935740
rect 676036 935688 676088 935740
rect 649908 935620 649960 935672
rect 678980 935620 679032 935672
rect 674748 935552 674800 935604
rect 676036 935552 676088 935604
rect 674472 935484 674524 935536
rect 676128 935484 676180 935536
rect 673644 935416 673696 935468
rect 675944 935416 675996 935468
rect 673552 935348 673604 935400
rect 675852 935348 675904 935400
rect 673736 935280 673788 935332
rect 675944 935280 675996 935332
rect 674840 934940 674892 934992
rect 676036 934940 676088 934992
rect 674656 932832 674708 932884
rect 676036 932832 676088 932884
rect 674012 932764 674064 932816
rect 676128 932764 676180 932816
rect 673828 932696 673880 932748
rect 675944 932696 675996 932748
rect 673920 932628 673972 932680
rect 676128 932628 676180 932680
rect 674288 932220 674340 932272
rect 676128 932220 676180 932272
rect 41788 932016 41840 932068
rect 46020 932016 46072 932068
rect 674380 931676 674432 931728
rect 676036 931676 676088 931728
rect 674564 931268 674616 931320
rect 676036 931268 676088 931320
rect 672080 927392 672132 927444
rect 678980 927392 679032 927444
rect 654876 922224 654928 922276
rect 669872 922224 669924 922276
rect 48596 921816 48648 921868
rect 58440 921816 58492 921868
rect 53840 908080 53892 908132
rect 59176 908080 59228 908132
rect 654876 908080 654928 908132
rect 663800 908080 663852 908132
rect 53932 896996 53984 897048
rect 58440 896996 58492 897048
rect 654876 895500 654928 895552
rect 661132 895500 661184 895552
rect 51080 883192 51132 883244
rect 58440 883192 58492 883244
rect 674656 873468 674708 873520
rect 675392 873468 675444 873520
rect 674748 872652 674800 872704
rect 675392 872652 675444 872704
rect 655152 870748 655204 870800
rect 674932 870748 674984 870800
rect 673644 869796 673696 869848
rect 675392 869796 675444 869848
rect 656808 869592 656860 869644
rect 663708 869592 663760 869644
rect 50988 869388 51040 869440
rect 58440 869388 58492 869440
rect 674196 868980 674248 869032
rect 675392 868980 675444 869032
rect 673736 868504 673788 868556
rect 675392 868504 675444 868556
rect 674288 867756 674340 867808
rect 675392 867756 675444 867808
rect 673828 866464 673880 866516
rect 675392 866464 675444 866516
rect 674932 866260 674984 866312
rect 675392 866260 675444 866312
rect 674012 864628 674064 864680
rect 675392 864628 675444 864680
rect 673920 862792 673972 862844
rect 675484 862792 675536 862844
rect 48688 858372 48740 858424
rect 58440 858372 58492 858424
rect 654692 855652 654744 855704
rect 661040 855652 661092 855704
rect 674656 854224 674708 854276
rect 675576 854224 675628 854276
rect 674748 854156 674800 854208
rect 675760 854156 675812 854208
rect 48780 844568 48832 844620
rect 58440 844568 58492 844620
rect 655060 841916 655112 841968
rect 668768 841916 668820 841968
rect 54024 830764 54076 830816
rect 57980 830764 58032 830816
rect 41788 817640 41840 817692
rect 53932 817640 53984 817692
rect 41788 817300 41840 817352
rect 51080 817300 51132 817352
rect 53748 817096 53800 817148
rect 59176 817096 59228 817148
rect 42708 817028 42760 817080
rect 62304 817028 62356 817080
rect 41154 816960 41206 817012
rect 41788 816960 41840 817012
rect 62488 816960 62540 817012
rect 654140 814716 654192 814768
rect 660948 814716 661000 814768
rect 41788 814240 41840 814292
rect 42892 814240 42944 814292
rect 62672 814240 62724 814292
rect 41788 808664 41840 808716
rect 44088 808664 44140 808716
rect 41788 808256 41840 808308
rect 42616 808256 42668 808308
rect 41788 806012 41840 806064
rect 42708 806012 42760 806064
rect 41972 805944 42024 805996
rect 48504 805944 48556 805996
rect 51080 805944 51132 805996
rect 58440 805944 58492 805996
rect 656808 803224 656860 803276
rect 666468 803224 666520 803276
rect 44272 800436 44324 800488
rect 48596 800436 48648 800488
rect 41880 800164 41932 800216
rect 43904 800164 43956 800216
rect 44088 800164 44140 800216
rect 42340 800028 42392 800080
rect 43904 800028 43956 800080
rect 41880 799960 41932 800012
rect 42156 798124 42208 798176
rect 42892 798124 42944 798176
rect 42892 797988 42944 798040
rect 43352 797988 43404 798040
rect 42616 797852 42668 797904
rect 42432 797580 42484 797632
rect 43352 797852 43404 797904
rect 43720 797852 43772 797904
rect 43720 797716 43772 797768
rect 43904 798124 43956 798176
rect 43904 797988 43956 798040
rect 44180 797988 44232 798040
rect 42156 797240 42208 797292
rect 44272 797240 44324 797292
rect 42156 796288 42208 796340
rect 43076 796288 43128 796340
rect 674748 796288 674800 796340
rect 675760 796288 675812 796340
rect 674564 796220 674616 796272
rect 675576 796220 675628 796272
rect 43076 796152 43128 796204
rect 44088 796152 44140 796204
rect 42156 794996 42208 795048
rect 42708 794996 42760 795048
rect 42156 794248 42208 794300
rect 43260 794248 43312 794300
rect 42156 793772 42208 793824
rect 42432 793772 42484 793824
rect 42156 792956 42208 793008
rect 43904 792956 43956 793008
rect 51264 792140 51316 792192
rect 58072 792140 58124 792192
rect 42156 790644 42208 790696
rect 43628 790644 43680 790696
rect 42156 790100 42208 790152
rect 43996 790100 44048 790152
rect 42156 789420 42208 789472
rect 43168 789420 43220 789472
rect 655060 789352 655112 789404
rect 663892 789352 663944 789404
rect 42156 788808 42208 788860
rect 43536 788808 43588 788860
rect 42156 786972 42208 787024
rect 42984 786972 43036 787024
rect 42064 786224 42116 786276
rect 43076 786224 43128 786276
rect 42156 785612 42208 785664
rect 43444 785612 43496 785664
rect 673460 784932 673512 784984
rect 675392 784932 675444 784984
rect 673552 782892 673604 782944
rect 675484 782892 675536 782944
rect 655520 782416 655572 782468
rect 674656 782416 674708 782468
rect 674288 780580 674340 780632
rect 675484 780580 675536 780632
rect 674472 779764 674524 779816
rect 675484 779764 675536 779816
rect 674196 779288 674248 779340
rect 675392 779288 675444 779340
rect 674380 778744 674432 778796
rect 674748 778744 674800 778796
rect 674748 778608 674800 778660
rect 675484 778608 675536 778660
rect 48596 778336 48648 778388
rect 58440 778336 58492 778388
rect 674380 777316 674432 777368
rect 675392 777316 675444 777368
rect 674656 777044 674708 777096
rect 675392 777044 675444 777096
rect 674564 775480 674616 775532
rect 675392 775480 675444 775532
rect 41512 774732 41564 774784
rect 48780 774732 48832 774784
rect 41512 774392 41564 774444
rect 54024 774392 54076 774444
rect 41512 773916 41564 773968
rect 48688 773916 48740 773968
rect 674656 773848 674708 773900
rect 675208 773848 675260 773900
rect 674656 773576 674708 773628
rect 675484 773576 675536 773628
rect 674472 773372 674524 773424
rect 675668 773372 675720 773424
rect 675208 773304 675260 773356
rect 675576 773304 675628 773356
rect 674748 773100 674800 773152
rect 675484 773100 675536 773152
rect 42892 772828 42944 772880
rect 62856 772828 62908 772880
rect 42064 772760 42116 772812
rect 62396 772760 62448 772812
rect 674288 770516 674340 770568
rect 674564 770516 674616 770568
rect 673552 770244 673604 770296
rect 674196 770244 674248 770296
rect 673460 770176 673512 770228
rect 674288 770176 674340 770228
rect 48780 767320 48832 767372
rect 58440 767320 58492 767372
rect 43628 766368 43680 766420
rect 43904 766368 43956 766420
rect 43628 766232 43680 766284
rect 44088 766232 44140 766284
rect 43260 766096 43312 766148
rect 44088 766096 44140 766148
rect 41512 762832 41564 762884
rect 46296 762832 46348 762884
rect 654784 762764 654836 762816
rect 668860 762764 668912 762816
rect 41788 760520 41840 760572
rect 50988 760520 51040 760572
rect 669872 759568 669924 759620
rect 676220 759568 676272 759620
rect 663800 759432 663852 759484
rect 678980 759432 679032 759484
rect 661132 759296 661184 759348
rect 676128 759296 676180 759348
rect 673368 759092 673420 759144
rect 676036 759092 676088 759144
rect 670516 759024 670568 759076
rect 676312 759024 676364 759076
rect 674012 758956 674064 759008
rect 676036 758956 676088 759008
rect 42064 757596 42116 757648
rect 42984 757596 43036 757648
rect 43444 757460 43496 757512
rect 43996 757460 44048 757512
rect 42156 757392 42208 757444
rect 43536 757392 43588 757444
rect 42708 757324 42760 757376
rect 43996 757324 44048 757376
rect 41880 756984 41932 757036
rect 41880 756712 41932 756764
rect 670608 756440 670660 756492
rect 676220 756440 676272 756492
rect 668400 756372 668452 756424
rect 676312 756372 676364 756424
rect 669964 756304 670016 756356
rect 670148 756304 670200 756356
rect 676128 756304 676180 756356
rect 669872 756236 669924 756288
rect 670332 756236 670384 756288
rect 678980 756236 679032 756288
rect 673920 756168 673972 756220
rect 676036 756168 676088 756220
rect 673644 756100 673696 756152
rect 676128 756100 676180 756152
rect 42432 755488 42484 755540
rect 42156 755420 42208 755472
rect 42156 755148 42208 755200
rect 42156 754876 42208 754928
rect 53840 753516 53892 753568
rect 58348 753516 58400 753568
rect 673828 753448 673880 753500
rect 676036 753448 676088 753500
rect 673736 753244 673788 753296
rect 676036 753244 676088 753296
rect 42156 753040 42208 753092
rect 43076 753040 43128 753092
rect 42156 751748 42208 751800
rect 42892 751748 42944 751800
rect 42156 751068 42208 751120
rect 43260 751068 43312 751120
rect 43260 750932 43312 750984
rect 43720 750932 43772 750984
rect 42064 750592 42116 750644
rect 43168 750592 43220 750644
rect 43168 750456 43220 750508
rect 43996 750456 44048 750508
rect 42156 749776 42208 749828
rect 43352 749776 43404 749828
rect 672172 749776 672224 749828
rect 678980 749776 679032 749828
rect 42616 749640 42668 749692
rect 43352 749640 43404 749692
rect 654876 748960 654928 749012
rect 668676 748960 668728 749012
rect 42156 746920 42208 746972
rect 43260 746920 43312 746972
rect 42156 746716 42208 746768
rect 43352 746716 43404 746768
rect 42156 746240 42208 746292
rect 43168 746240 43220 746292
rect 42156 745424 42208 745476
rect 43628 745424 43680 745476
rect 42156 743724 42208 743776
rect 43444 743724 43496 743776
rect 42156 743044 42208 743096
rect 43904 743044 43956 743096
rect 42156 742568 42208 742620
rect 43996 742568 44048 742620
rect 48688 739712 48740 739764
rect 58440 739712 58492 739764
rect 673920 738420 673972 738472
rect 674656 738420 674708 738472
rect 655520 738284 655572 738336
rect 674656 738284 674708 738336
rect 654784 735972 654836 736024
rect 661132 735972 661184 736024
rect 674012 735428 674064 735480
rect 675392 735428 675444 735480
rect 673644 734952 673696 735004
rect 675392 734952 675444 735004
rect 673828 734340 673880 734392
rect 675392 734340 675444 734392
rect 673552 733592 673604 733644
rect 675392 733592 675444 733644
rect 673736 732300 673788 732352
rect 675392 732300 675444 732352
rect 674656 732028 674708 732080
rect 675392 732028 675444 732080
rect 674012 731892 674064 731944
rect 674656 731892 674708 731944
rect 673920 731824 673972 731876
rect 673920 731552 673972 731604
rect 673644 730464 673696 730516
rect 675392 730464 675444 730516
rect 41512 729648 41564 729700
rect 43536 729648 43588 729700
rect 42524 729512 42576 729564
rect 43076 729512 43128 729564
rect 41788 728832 41840 728884
rect 44364 728832 44416 728884
rect 42524 728696 42576 728748
rect 62396 728696 62448 728748
rect 675668 728628 675720 728680
rect 675668 728356 675720 728408
rect 51172 725908 51224 725960
rect 58440 725908 58492 725960
rect 673368 723120 673420 723172
rect 678980 723120 679032 723172
rect 41512 719584 41564 719636
rect 48596 719584 48648 719636
rect 674196 718088 674248 718140
rect 674840 718088 674892 718140
rect 673920 717952 673972 718004
rect 674196 717952 674248 718004
rect 673644 717612 673696 717664
rect 673920 717612 673972 717664
rect 41328 717544 41380 717596
rect 43720 717544 43772 717596
rect 42524 716592 42576 716644
rect 53748 716592 53800 716644
rect 663708 716116 663760 716168
rect 675944 716116 675996 716168
rect 668768 715708 668820 715760
rect 675944 715708 675996 715760
rect 670516 715300 670568 715352
rect 675944 715300 675996 715352
rect 661040 714960 661092 715012
rect 676036 714960 676088 715012
rect 670148 714892 670200 714944
rect 670516 714892 670568 714944
rect 50988 714824 51040 714876
rect 58440 714824 58492 714876
rect 670240 714824 670292 714876
rect 676036 714824 676088 714876
rect 673092 714008 673144 714060
rect 676036 714008 676088 714060
rect 41880 713804 41932 713856
rect 668400 713668 668452 713720
rect 670332 713668 670384 713720
rect 676036 713668 676088 713720
rect 41880 713532 41932 713584
rect 668952 713192 669004 713244
rect 670516 713192 670568 713244
rect 676036 713192 676088 713244
rect 668768 712784 668820 712836
rect 670608 712784 670660 712836
rect 676036 712784 676088 712836
rect 669044 712376 669096 712428
rect 676036 712376 676088 712428
rect 674748 712036 674800 712088
rect 676036 712036 676088 712088
rect 674564 711968 674616 712020
rect 675944 711968 675996 712020
rect 674288 711900 674340 711952
rect 675852 711900 675904 711952
rect 674196 711832 674248 711884
rect 675760 711832 675812 711884
rect 42156 711628 42208 711680
rect 42892 711628 42944 711680
rect 42984 711356 43036 711408
rect 43628 711356 43680 711408
rect 42156 711084 42208 711136
rect 42524 711084 42576 711136
rect 673828 710812 673880 710864
rect 675484 710812 675536 710864
rect 673552 710676 673604 710728
rect 673828 710676 673880 710728
rect 674656 710676 674708 710728
rect 675576 710676 675628 710728
rect 42156 709860 42208 709912
rect 42800 709860 42852 709912
rect 42800 709724 42852 709776
rect 43260 709724 43312 709776
rect 655980 709724 656032 709776
rect 666928 709724 666980 709776
rect 674472 709248 674524 709300
rect 676036 709248 676088 709300
rect 42156 708568 42208 708620
rect 43168 708568 43220 708620
rect 674380 708228 674432 708280
rect 676036 708228 676088 708280
rect 42156 708024 42208 708076
rect 43904 708024 43956 708076
rect 674840 707820 674892 707872
rect 676036 707820 676088 707872
rect 676036 707412 676088 707464
rect 676956 707412 677008 707464
rect 42156 707344 42208 707396
rect 43812 707344 43864 707396
rect 42156 706732 42208 706784
rect 43260 706732 43312 706784
rect 671804 705100 671856 705152
rect 676036 705100 676088 705152
rect 42248 704828 42300 704880
rect 43076 704828 43128 704880
rect 42064 704216 42116 704268
rect 43996 704216 44048 704268
rect 42064 702856 42116 702908
rect 43720 702856 43772 702908
rect 42064 702380 42116 702432
rect 43444 702380 43496 702432
rect 53748 701020 53800 701072
rect 58624 701020 58676 701072
rect 42156 700408 42208 700460
rect 43536 700408 43588 700460
rect 42156 700000 42208 700052
rect 42892 700000 42944 700052
rect 674564 699728 674616 699780
rect 675576 699728 675628 699780
rect 674748 699660 674800 699712
rect 675484 699660 675536 699712
rect 674656 699592 674708 699644
rect 675668 699592 675720 699644
rect 42064 699388 42116 699440
rect 42800 699388 42852 699440
rect 654692 695512 654744 695564
rect 663708 695512 663760 695564
rect 655520 691364 655572 691416
rect 674472 691364 674524 691416
rect 673736 690412 673788 690464
rect 675392 690412 675444 690464
rect 673184 689120 673236 689172
rect 675484 689120 675536 689172
rect 673000 688576 673052 688628
rect 675392 688576 675444 688628
rect 41512 688372 41564 688424
rect 48688 688372 48740 688424
rect 41696 688032 41748 688084
rect 53840 688032 53892 688084
rect 41788 687692 41840 687744
rect 51172 687692 51224 687744
rect 673276 687284 673328 687336
rect 675392 687284 675444 687336
rect 51080 687216 51132 687268
rect 58440 687216 58492 687268
rect 674472 687012 674524 687064
rect 675484 687012 675536 687064
rect 673828 685448 673880 685500
rect 675392 685448 675444 685500
rect 674288 683612 674340 683664
rect 675484 683612 675536 683664
rect 654876 682932 654928 682984
rect 663800 682932 663852 682984
rect 42800 681640 42852 681692
rect 62948 681640 63000 681692
rect 673092 678988 673144 679040
rect 678980 678988 679032 679040
rect 41788 678308 41840 678360
rect 44088 678308 44140 678360
rect 41788 676608 41840 676660
rect 48688 676608 48740 676660
rect 48872 673480 48924 673532
rect 58440 673480 58492 673532
rect 41328 673412 41380 673464
rect 42892 673412 42944 673464
rect 666468 671508 666520 671560
rect 676220 671508 676272 671560
rect 674748 671236 674800 671288
rect 675208 671236 675260 671288
rect 660948 670760 661000 670812
rect 676036 670760 676088 670812
rect 44180 670692 44232 670744
rect 48780 670692 48832 670744
rect 43812 670624 43864 670676
rect 43996 670624 44048 670676
rect 44088 670624 44140 670676
rect 41880 670556 41932 670608
rect 41972 670556 42024 670608
rect 42708 670556 42760 670608
rect 41880 670352 41932 670404
rect 43812 670420 43864 670472
rect 43996 670420 44048 670472
rect 663892 670556 663944 670608
rect 676036 670556 676088 670608
rect 670240 670284 670292 670336
rect 676220 670284 676272 670336
rect 44180 670148 44232 670200
rect 669136 669740 669188 669792
rect 674472 669740 674524 669792
rect 676036 669740 676088 669792
rect 670516 668652 670568 668704
rect 676220 668652 676272 668704
rect 42064 668448 42116 668500
rect 43904 668448 43956 668500
rect 673092 668040 673144 668092
rect 675944 668040 675996 668092
rect 674748 667904 674800 667956
rect 676036 667904 676088 667956
rect 673920 667836 673972 667888
rect 676128 667836 676180 667888
rect 674564 667768 674616 667820
rect 676036 667768 676088 667820
rect 42156 667700 42208 667752
rect 44088 667700 44140 667752
rect 669044 667700 669096 667752
rect 675944 667700 675996 667752
rect 42156 666680 42208 666732
rect 43720 666680 43772 666732
rect 42156 665388 42208 665440
rect 42708 665388 42760 665440
rect 674656 665116 674708 665168
rect 676036 665116 676088 665168
rect 675208 664708 675260 664760
rect 676036 664708 676088 664760
rect 42156 664640 42208 664692
rect 43536 664640 43588 664692
rect 42156 663960 42208 664012
rect 43996 663960 44048 664012
rect 42156 663552 42208 663604
rect 42892 663552 42944 663604
rect 48964 662396 49016 662448
rect 58440 662396 58492 662448
rect 42156 661036 42208 661088
rect 43812 661036 43864 661088
rect 42156 660492 42208 660544
rect 43444 660492 43496 660544
rect 42156 659880 42208 659932
rect 43260 659880 43312 659932
rect 672356 659676 672408 659728
rect 678980 659676 679032 659728
rect 42156 659200 42208 659252
rect 42984 659200 43036 659252
rect 42156 657228 42208 657280
rect 43628 657228 43680 657280
rect 656164 657024 656216 657076
rect 660948 657024 661000 657076
rect 42156 656820 42208 656872
rect 44088 656820 44140 656872
rect 42156 656140 42208 656192
rect 43076 656140 43128 656192
rect 673552 649544 673604 649596
rect 675392 649544 675444 649596
rect 53840 648592 53892 648644
rect 59176 648592 59228 648644
rect 674656 647708 674708 647760
rect 675484 647708 675536 647760
rect 673460 647300 673512 647352
rect 674748 647300 674800 647352
rect 655520 647164 655572 647216
rect 674748 647164 674800 647216
rect 673920 645396 673972 645448
rect 675392 645396 675444 645448
rect 41512 645124 41564 645176
rect 51080 645124 51132 645176
rect 41512 644784 41564 644836
rect 53748 644784 53800 644836
rect 674564 644784 674616 644836
rect 675392 644784 675444 644836
rect 41788 644512 41840 644564
rect 48872 644512 48924 644564
rect 673644 644104 673696 644156
rect 675392 644104 675444 644156
rect 674380 643356 674432 643408
rect 675392 643356 675444 643408
rect 654876 643084 654928 643136
rect 663892 643084 663944 643136
rect 674012 642064 674064 642116
rect 675392 642064 675444 642116
rect 674748 641860 674800 641912
rect 675392 641860 675444 641912
rect 674196 640228 674248 640280
rect 675392 640228 675444 640280
rect 674656 638800 674708 638852
rect 675208 638664 675260 638716
rect 674564 638392 674616 638444
rect 675484 638392 675536 638444
rect 675208 638188 675260 638240
rect 675668 638188 675720 638240
rect 673092 637848 673144 637900
rect 679164 637848 679216 637900
rect 673460 637508 673512 637560
rect 679072 637508 679124 637560
rect 48872 634788 48924 634840
rect 58440 634788 58492 634840
rect 41512 633224 41564 633276
rect 48780 633224 48832 633276
rect 43628 629280 43680 629332
rect 50988 629280 51040 629332
rect 655060 629280 655112 629332
rect 669044 629280 669096 629332
rect 30288 627852 30340 627904
rect 42524 627852 42576 627904
rect 41788 627376 41840 627428
rect 41788 627036 41840 627088
rect 674472 626492 674524 626544
rect 676036 626492 676088 626544
rect 42156 625268 42208 625320
rect 43720 625268 43772 625320
rect 42156 624656 42208 624708
rect 43628 624656 43680 624708
rect 668860 624112 668912 624164
rect 676220 624112 676272 624164
rect 668676 623976 668728 624028
rect 678980 623976 679032 624028
rect 673368 623908 673420 623960
rect 676036 623908 676088 623960
rect 661132 623840 661184 623892
rect 676312 623840 676364 623892
rect 51080 623772 51132 623824
rect 58440 623772 58492 623824
rect 668584 623772 668636 623824
rect 670608 623772 670660 623824
rect 676128 623772 676180 623824
rect 673828 623704 673880 623756
rect 676036 623704 676088 623756
rect 42156 623432 42208 623484
rect 43076 623432 43128 623484
rect 42064 622140 42116 622192
rect 42524 622140 42576 622192
rect 42156 621460 42208 621512
rect 43260 621460 43312 621512
rect 670240 621052 670292 621104
rect 678980 621052 679032 621104
rect 42064 620984 42116 621036
rect 43168 620984 43220 621036
rect 668492 620984 668544 621036
rect 670516 620984 670568 621036
rect 676220 620984 676272 621036
rect 674288 620916 674340 620968
rect 676036 620916 676088 620968
rect 673736 620848 673788 620900
rect 676128 620848 676180 620900
rect 42064 620168 42116 620220
rect 43904 620168 43956 620220
rect 42248 619012 42300 619064
rect 42892 619012 42944 619064
rect 673276 618196 673328 618248
rect 676036 618196 676088 618248
rect 673184 617924 673236 617976
rect 676220 617924 676272 617976
rect 42156 617856 42208 617908
rect 43812 617856 43864 617908
rect 42064 617312 42116 617364
rect 43444 617312 43496 617364
rect 673000 616700 673052 616752
rect 676220 616700 676272 616752
rect 42248 616020 42300 616072
rect 43536 616020 43588 616072
rect 672448 614592 672500 614644
rect 678980 614592 679032 614644
rect 42156 614184 42208 614236
rect 43352 614184 43404 614236
rect 42156 613640 42208 613692
rect 42984 613640 43036 613692
rect 42156 612960 42208 613012
rect 42800 612960 42852 613012
rect 50988 609968 51040 610020
rect 58440 609968 58492 610020
rect 674472 608744 674524 608796
rect 675668 608744 675720 608796
rect 654600 603032 654652 603084
rect 674656 603032 674708 603084
rect 654324 602148 654376 602200
rect 661040 602148 661092 602200
rect 41512 601876 41564 601928
rect 48872 601876 48924 601928
rect 674288 600380 674340 600432
rect 675484 600380 675536 600432
rect 674748 599564 674800 599616
rect 675484 599564 675536 599616
rect 673736 598952 673788 599004
rect 675392 598952 675444 599004
rect 42432 598884 42484 598936
rect 62764 598884 62816 598936
rect 673460 598408 673512 598460
rect 675484 598408 675536 598460
rect 673828 597116 673880 597168
rect 675392 597116 675444 597168
rect 674656 596844 674708 596896
rect 675392 596844 675444 596896
rect 674472 596572 674524 596624
rect 674748 596572 674800 596624
rect 53748 596164 53800 596216
rect 59176 596164 59228 596216
rect 674472 595280 674524 595332
rect 675392 595280 675444 595332
rect 674380 593648 674432 593700
rect 675484 593648 675536 593700
rect 656808 590656 656860 590708
rect 669136 590656 669188 590708
rect 41512 589976 41564 590028
rect 48872 589976 48924 590028
rect 673368 587868 673420 587920
rect 678980 587868 679032 587920
rect 43352 586712 43404 586764
rect 44088 586712 44140 586764
rect 42800 586576 42852 586628
rect 43352 586576 43404 586628
rect 41144 585148 41196 585200
rect 44180 585148 44232 585200
rect 44272 585148 44324 585200
rect 48964 585148 49016 585200
rect 673368 584264 673420 584316
rect 673552 584264 673604 584316
rect 41880 584196 41932 584248
rect 673552 584128 673604 584180
rect 673920 584128 673972 584180
rect 674748 583992 674800 584044
rect 675668 583992 675720 584044
rect 41880 583924 41932 583976
rect 674472 583856 674524 583908
rect 674748 583856 674800 583908
rect 42432 583720 42484 583772
rect 42800 583720 42852 583772
rect 42892 583720 42944 583772
rect 43076 583720 43128 583772
rect 673460 583720 673512 583772
rect 673828 583720 673880 583772
rect 673920 583652 673972 583704
rect 674380 583652 674432 583704
rect 43076 583584 43128 583636
rect 43260 583584 43312 583636
rect 43260 583448 43312 583500
rect 43996 583448 44048 583500
rect 44088 583448 44140 583500
rect 44088 583108 44140 583160
rect 48964 582360 49016 582412
rect 58440 582360 58492 582412
rect 42156 582088 42208 582140
rect 42708 582088 42760 582140
rect 42156 581272 42208 581324
rect 44272 581272 44324 581324
rect 42156 580252 42208 580304
rect 43352 580252 43404 580304
rect 670608 580184 670660 580236
rect 676036 580184 676088 580236
rect 666928 580048 666980 580100
rect 676128 580048 676180 580100
rect 663800 579912 663852 579964
rect 676220 579912 676272 579964
rect 663708 579776 663760 579828
rect 676312 579776 676364 579828
rect 672540 579232 672592 579284
rect 673276 579232 673328 579284
rect 676220 579232 676272 579284
rect 42156 578960 42208 579012
rect 43536 578960 43588 579012
rect 42156 578416 42208 578468
rect 43720 578416 43772 578468
rect 673092 578416 673144 578468
rect 676220 578416 676272 578468
rect 42156 577804 42208 577856
rect 43628 577804 43680 577856
rect 43628 577668 43680 577720
rect 43996 577668 44048 577720
rect 672632 577600 672684 577652
rect 673184 577600 673236 577652
rect 676220 577600 676272 577652
rect 42156 576920 42208 576972
rect 44088 576920 44140 576972
rect 670516 576920 670568 576972
rect 676220 576920 676272 576972
rect 655060 576852 655112 576904
rect 663708 576852 663760 576904
rect 673368 576852 673420 576904
rect 676036 576852 676088 576904
rect 674196 576784 674248 576836
rect 675944 576784 675996 576836
rect 674564 576716 674616 576768
rect 676036 576716 676088 576768
rect 673460 576648 673512 576700
rect 676128 576648 676180 576700
rect 673552 576036 673604 576088
rect 675944 576036 675996 576088
rect 42156 574676 42208 574728
rect 43904 574676 43956 574728
rect 42156 573792 42208 573844
rect 43168 573792 43220 573844
rect 674012 573588 674064 573640
rect 676036 573588 676088 573640
rect 42156 573452 42208 573504
rect 43628 573452 43680 573504
rect 673644 572772 673696 572824
rect 676036 572772 676088 572824
rect 42064 572636 42116 572688
rect 43812 572636 43864 572688
rect 42064 570868 42116 570920
rect 43076 570868 43128 570920
rect 42156 570256 42208 570308
rect 42984 570256 43036 570308
rect 42064 569576 42116 569628
rect 42892 569576 42944 569628
rect 672540 568556 672592 568608
rect 678980 568556 679032 568608
rect 673552 559512 673604 559564
rect 675484 559512 675536 559564
rect 41512 558764 41564 558816
rect 48964 558764 49016 558816
rect 41420 558492 41472 558544
rect 53748 558492 53800 558544
rect 41512 558424 41564 558476
rect 58440 558424 58492 558476
rect 49056 557540 49108 557592
rect 58348 557540 58400 557592
rect 654324 556112 654376 556164
rect 675300 556112 675352 556164
rect 673920 555228 673972 555280
rect 675392 555228 675444 555280
rect 673460 554548 673512 554600
rect 675392 554548 675444 554600
rect 674012 553732 674064 553784
rect 675392 553732 675444 553784
rect 673644 553188 673696 553240
rect 675392 553188 675444 553240
rect 674196 551896 674248 551948
rect 675392 551896 675444 551948
rect 654692 549244 654744 549296
rect 663800 549244 663852 549296
rect 41512 548632 41564 548684
rect 43536 548632 43588 548684
rect 674564 548292 674616 548344
rect 675392 548292 675444 548344
rect 674656 548224 674708 548276
rect 675300 548224 675352 548276
rect 41604 546864 41656 546916
rect 48964 546864 49016 546916
rect 41512 546728 41564 546780
rect 42800 546728 42852 546780
rect 673092 546252 673144 546304
rect 679072 546252 679124 546304
rect 53840 543736 53892 543788
rect 58348 543736 58400 543788
rect 43720 541696 43772 541748
rect 50988 541696 51040 541748
rect 41788 541016 41840 541068
rect 41788 540744 41840 540796
rect 42064 538908 42116 538960
rect 42708 538908 42760 538960
rect 42156 538092 42208 538144
rect 43720 538092 43772 538144
rect 42064 537072 42116 537124
rect 42984 537072 43036 537124
rect 42984 536936 43036 536988
rect 43168 536936 43220 536988
rect 43168 536800 43220 536852
rect 43352 536800 43404 536852
rect 43352 536664 43404 536716
rect 43628 536664 43680 536716
rect 654876 536392 654928 536444
rect 666468 536392 666520 536444
rect 42156 535780 42208 535832
rect 42800 535780 42852 535832
rect 663892 535712 663944 535764
rect 676220 535712 676272 535764
rect 660948 535576 661000 535628
rect 676036 535576 676088 535628
rect 42064 535032 42116 535084
rect 43260 535032 43312 535084
rect 673276 534896 673328 534948
rect 676036 534896 676088 534948
rect 42156 534420 42208 534472
rect 43536 534420 43588 534472
rect 42156 533944 42208 533996
rect 43352 533944 43404 533996
rect 673184 533264 673236 533316
rect 676036 533264 676088 533316
rect 669044 532856 669096 532908
rect 678980 532856 679032 532908
rect 670056 532788 670108 532840
rect 675852 532788 675904 532840
rect 676128 532788 676180 532840
rect 674748 532652 674800 532704
rect 676036 532652 676088 532704
rect 672816 532584 672868 532636
rect 673368 532584 673420 532636
rect 676220 532584 676272 532636
rect 42156 531428 42208 531480
rect 43904 531428 43956 531480
rect 674288 531088 674340 531140
rect 676036 531088 676088 531140
rect 42156 530680 42208 530732
rect 43996 530680 44048 530732
rect 42156 530272 42208 530324
rect 43076 530272 43128 530324
rect 674472 529864 674524 529916
rect 676036 529864 676088 529916
rect 42156 529456 42208 529508
rect 43168 529456 43220 529508
rect 674380 529456 674432 529508
rect 676036 529456 676088 529508
rect 673736 527824 673788 527876
rect 676036 527824 676088 527876
rect 42156 527212 42208 527264
rect 43444 527212 43496 527264
rect 42064 527144 42116 527196
rect 43812 527144 43864 527196
rect 673828 527076 673880 527128
rect 676036 527076 676088 527128
rect 42156 526600 42208 526652
rect 42984 526600 43036 526652
rect 672632 524424 672684 524476
rect 678980 524424 679032 524476
rect 677498 524356 677550 524408
rect 679072 524356 679124 524408
rect 675852 523948 675904 524000
rect 676128 523948 676180 524000
rect 654140 522452 654192 522504
rect 661224 522452 661276 522504
rect 51264 518916 51316 518968
rect 58440 518916 58492 518968
rect 654876 510824 654928 510876
rect 670516 510824 670568 510876
rect 50988 505112 51040 505164
rect 58440 505112 58492 505164
rect 656808 497632 656860 497684
rect 663892 497632 663944 497684
rect 675576 492192 675628 492244
rect 676036 492192 676088 492244
rect 669136 491648 669188 491700
rect 676036 491648 676088 491700
rect 663708 491512 663760 491564
rect 676036 491512 676088 491564
rect 661040 491376 661092 491428
rect 675944 491376 675996 491428
rect 49148 491308 49200 491360
rect 57980 491308 58032 491360
rect 676220 491240 676272 491292
rect 677508 491240 677560 491292
rect 669688 488520 669740 488572
rect 675668 488520 675720 488572
rect 675944 488520 675996 488572
rect 674656 488180 674708 488232
rect 676036 488180 676088 488232
rect 673552 487908 673604 487960
rect 675668 487908 675720 487960
rect 673920 487092 673972 487144
rect 676036 487092 676088 487144
rect 669688 485800 669740 485852
rect 675576 485800 675628 485852
rect 674564 485732 674616 485784
rect 676036 485732 676088 485784
rect 674196 485460 674248 485512
rect 676036 485460 676088 485512
rect 654876 483012 654928 483064
rect 669136 483012 669188 483064
rect 673644 482944 673696 482996
rect 676036 482944 676088 482996
rect 673460 482876 673512 482928
rect 675668 482876 675720 482928
rect 672724 480700 672776 480752
rect 676036 480700 676088 480752
rect 51172 480224 51224 480276
rect 58440 480224 58492 480276
rect 675944 478592 675996 478644
rect 676036 478388 676088 478440
rect 654876 470772 654928 470824
rect 660948 470772 661000 470824
rect 54024 466420 54076 466472
rect 58716 466420 58768 466472
rect 654232 457444 654284 457496
rect 667020 457444 667072 457496
rect 53748 452616 53800 452668
rect 59176 452616 59228 452668
rect 654416 444456 654468 444508
rect 663984 444456 664036 444508
rect 51080 438880 51132 438932
rect 58440 438880 58492 438932
rect 41788 430788 41840 430840
rect 59268 430788 59320 430840
rect 654692 430584 654744 430636
rect 663708 430584 663760 430636
rect 53932 427864 53984 427916
rect 58256 427864 58308 427916
rect 41788 427796 41840 427848
rect 44088 427796 44140 427848
rect 62764 427796 62816 427848
rect 41788 419432 41840 419484
rect 46664 419432 46716 419484
rect 655060 416780 655112 416832
rect 661040 416780 661092 416832
rect 41880 416304 41932 416356
rect 43076 416304 43128 416356
rect 49240 413992 49292 414044
rect 58440 413992 58492 414044
rect 42156 413108 42208 413160
rect 42340 413108 42392 413160
rect 42800 411340 42852 411392
rect 42156 411272 42208 411324
rect 675760 411068 675812 411120
rect 676128 411068 676180 411120
rect 42156 410660 42208 410712
rect 49056 410660 49108 410712
rect 42156 409436 42208 409488
rect 42984 409436 43036 409488
rect 42064 408144 42116 408196
rect 42524 408144 42576 408196
rect 42156 407464 42208 407516
rect 43168 407464 43220 407516
rect 42064 406988 42116 407040
rect 43076 406988 43128 407040
rect 42156 406172 42208 406224
rect 43444 406172 43496 406224
rect 654876 403996 654928 404048
rect 661132 403996 661184 404048
rect 42156 403860 42208 403912
rect 43996 403860 44048 403912
rect 666468 403384 666520 403436
rect 676220 403384 676272 403436
rect 42156 403316 42208 403368
rect 43536 403316 43588 403368
rect 663800 403248 663852 403300
rect 676220 403248 676272 403300
rect 661224 403112 661276 403164
rect 675944 403112 675996 403164
rect 42156 402500 42208 402552
rect 43720 402500 43772 402552
rect 43812 402432 43864 402484
rect 43812 402228 43864 402280
rect 42156 402024 42208 402076
rect 43352 402024 43404 402076
rect 675116 400392 675168 400444
rect 676128 400392 676180 400444
rect 49056 400188 49108 400240
rect 58440 400188 58492 400240
rect 42156 399984 42208 400036
rect 42892 399984 42944 400036
rect 42156 399440 42208 399492
rect 43720 399440 43772 399492
rect 674380 399440 674432 399492
rect 676036 399440 676088 399492
rect 42156 398760 42208 398812
rect 43260 398760 43312 398812
rect 674472 398216 674524 398268
rect 676036 398216 676088 398268
rect 673828 397604 673880 397656
rect 675944 397604 675996 397656
rect 674288 397536 674340 397588
rect 676128 397536 676180 397588
rect 674656 397468 674708 397520
rect 676036 397468 676088 397520
rect 673460 396584 673512 396636
rect 676036 396584 676088 396636
rect 673552 395360 673604 395412
rect 675944 395360 675996 395412
rect 675024 394952 675076 395004
rect 676036 394952 676088 395004
rect 673644 394816 673696 394868
rect 675944 394816 675996 394868
rect 674932 394748 674984 394800
rect 676128 394748 676180 394800
rect 675208 394680 675260 394732
rect 676036 394680 676088 394732
rect 672908 392096 672960 392148
rect 679072 392096 679124 392148
rect 673736 392028 673788 392080
rect 676128 392028 676180 392080
rect 674012 391960 674064 392012
rect 676036 391960 676088 392012
rect 674748 390532 674800 390584
rect 675760 390532 675812 390584
rect 674564 390464 674616 390516
rect 675668 390464 675720 390516
rect 654324 389852 654376 389904
rect 666468 389852 666520 389904
rect 53840 389172 53892 389224
rect 57980 389172 58032 389224
rect 41512 387948 41564 388000
rect 51172 387948 51224 388000
rect 41512 387608 41564 387660
rect 54024 387608 54076 387660
rect 41512 387132 41564 387184
rect 49148 387132 49200 387184
rect 42800 386384 42852 386436
rect 63132 386384 63184 386436
rect 675760 386384 675812 386436
rect 675760 386112 675812 386164
rect 674472 384956 674524 385008
rect 675300 384956 675352 385008
rect 675208 384072 675260 384124
rect 675300 383868 675352 383920
rect 674656 383120 674708 383172
rect 675392 383120 675444 383172
rect 674380 382984 674432 383036
rect 674656 382984 674708 383036
rect 675024 382440 675076 382492
rect 675392 382440 675444 382492
rect 674932 381896 674984 381948
rect 675392 381896 675444 381948
rect 673828 379448 673880 379500
rect 675300 379448 675352 379500
rect 656808 378156 656860 378208
rect 670056 378156 670108 378208
rect 674012 378156 674064 378208
rect 675484 378156 675536 378208
rect 673644 378088 673696 378140
rect 675300 378088 675352 378140
rect 673736 376932 673788 376984
rect 675484 376932 675536 376984
rect 673552 376864 673604 376916
rect 675300 376864 675352 376916
rect 41604 376048 41656 376100
rect 46848 376048 46900 376100
rect 49148 375368 49200 375420
rect 58440 375368 58492 375420
rect 675116 374076 675168 374128
rect 675300 374076 675352 374128
rect 674288 373872 674340 373924
rect 675392 373872 675444 373924
rect 675300 372852 675352 372904
rect 675300 372648 675352 372700
rect 673460 372036 673512 372088
rect 675392 372036 675444 372088
rect 41512 371424 41564 371476
rect 42708 371424 42760 371476
rect 674748 370744 674800 370796
rect 675760 370744 675812 370796
rect 674564 370676 674616 370728
rect 675668 370676 675720 370728
rect 42156 369928 42208 369980
rect 42340 369928 42392 369980
rect 42156 368092 42208 368144
rect 42800 368092 42852 368144
rect 42156 366800 42208 366852
rect 50988 366800 51040 366852
rect 42156 366256 42208 366308
rect 42892 366256 42944 366308
rect 42892 366120 42944 366172
rect 43444 366120 43496 366172
rect 42156 364964 42208 365016
rect 42708 364964 42760 365016
rect 42156 364420 42208 364472
rect 43168 364420 43220 364472
rect 656808 364420 656860 364472
rect 669044 364420 669096 364472
rect 42156 363808 42208 363860
rect 43076 363808 43128 363860
rect 43076 363672 43128 363724
rect 43628 363672 43680 363724
rect 42156 363128 42208 363180
rect 43904 363128 43956 363180
rect 51172 361564 51224 361616
rect 58440 361564 58492 361616
rect 42064 360680 42116 360732
rect 43260 360680 43312 360732
rect 42156 359932 42208 359984
rect 43628 359932 43680 359984
rect 42156 359456 42208 359508
rect 43076 359456 43128 359508
rect 42064 358640 42116 358692
rect 42984 358640 43036 358692
rect 673276 357008 673328 357060
rect 675760 357008 675812 357060
rect 42064 356940 42116 356992
rect 43352 356940 43404 356992
rect 670516 356464 670568 356516
rect 675944 356464 675996 356516
rect 42156 356396 42208 356448
rect 42892 356396 42944 356448
rect 669136 356328 669188 356380
rect 676036 356328 676088 356380
rect 663892 356192 663944 356244
rect 675852 356192 675904 356244
rect 673368 356124 673420 356176
rect 676036 356124 676088 356176
rect 669596 356056 669648 356108
rect 673000 356056 673052 356108
rect 673276 356056 673328 356108
rect 673184 355376 673236 355428
rect 676036 355376 676088 355428
rect 673276 354560 673328 354612
rect 676036 354560 676088 354612
rect 669504 353472 669556 353524
rect 673092 353472 673144 353524
rect 673276 353472 673328 353524
rect 673828 353472 673880 353524
rect 676036 353472 676088 353524
rect 669412 353336 669464 353388
rect 673184 353336 673236 353388
rect 674104 353268 674156 353320
rect 676036 353268 676088 353320
rect 673000 351772 673052 351824
rect 673276 351772 673328 351824
rect 674196 351432 674248 351484
rect 676036 351432 676088 351484
rect 673460 351024 673512 351076
rect 675944 351024 675996 351076
rect 673920 350616 673972 350668
rect 675944 350616 675996 350668
rect 654876 350548 654928 350600
rect 669504 350548 669556 350600
rect 674288 350548 674340 350600
rect 676036 350548 676088 350600
rect 673736 349800 673788 349852
rect 676036 349800 676088 349852
rect 673644 348984 673696 349036
rect 675944 348984 675996 349036
rect 673552 347828 673604 347880
rect 675944 347828 675996 347880
rect 50988 347760 51040 347812
rect 58440 347760 58492 347812
rect 674012 347760 674064 347812
rect 676036 347760 676088 347812
rect 673000 347216 673052 347268
rect 676036 347216 676088 347268
rect 44180 344972 44232 345024
rect 48412 344972 48464 345024
rect 41512 344700 41564 344752
rect 43536 344700 43588 344752
rect 41788 344428 41840 344480
rect 53932 344428 53984 344480
rect 41604 344292 41656 344344
rect 49240 344292 49292 344344
rect 41604 343884 41656 343936
rect 51080 343884 51132 343936
rect 41788 343340 41840 343392
rect 44180 343340 44232 343392
rect 674104 340960 674156 341012
rect 675484 340960 675536 341012
rect 673828 339532 673880 339584
rect 675484 339532 675536 339584
rect 674196 337900 674248 337952
rect 675484 337900 675536 337952
rect 674288 337220 674340 337272
rect 675392 337220 675444 337272
rect 48412 336744 48464 336796
rect 58440 336744 58492 336796
rect 655060 336744 655112 336796
rect 666928 336744 666980 336796
rect 673920 336540 673972 336592
rect 675392 336540 675444 336592
rect 674012 335860 674064 335912
rect 675484 335860 675536 335912
rect 673460 333548 673512 333600
rect 675392 333548 675444 333600
rect 673644 332936 673696 332988
rect 675392 332936 675444 332988
rect 41512 332800 41564 332852
rect 46204 332800 46256 332852
rect 673736 332392 673788 332444
rect 675392 332392 675444 332444
rect 673552 331576 673604 331628
rect 675392 331576 675444 331628
rect 33048 330080 33100 330132
rect 41880 330080 41932 330132
rect 32864 329944 32916 329996
rect 42892 329944 42944 329996
rect 32956 329876 33008 329928
rect 43352 329876 43404 329928
rect 32680 329808 32732 329860
rect 42800 329808 42852 329860
rect 41880 326952 41932 327004
rect 41880 326748 41932 326800
rect 42064 324912 42116 324964
rect 42800 324912 42852 324964
rect 42800 324776 42852 324828
rect 43076 324776 43128 324828
rect 43168 324776 43220 324828
rect 43168 324572 43220 324624
rect 654876 323892 654928 323944
rect 669136 323892 669188 323944
rect 53932 323484 53984 323536
rect 58164 323484 58216 323536
rect 42156 323280 42208 323332
rect 42616 323280 42668 323332
rect 42064 323076 42116 323128
rect 42892 323076 42944 323128
rect 42156 321784 42208 321836
rect 43168 321784 43220 321836
rect 42156 321036 42208 321088
rect 43352 321036 43404 321088
rect 42156 320560 42208 320612
rect 42984 320560 43036 320612
rect 42616 320084 42668 320136
rect 53748 320084 53800 320136
rect 42156 317432 42208 317484
rect 42800 317432 42852 317484
rect 658464 314576 658516 314628
rect 671160 314576 671212 314628
rect 667020 313692 667072 313744
rect 676036 313692 676088 313744
rect 663984 312876 664036 312928
rect 676036 312876 676088 312928
rect 673276 312468 673328 312520
rect 676036 312468 676088 312520
rect 671160 312060 671212 312112
rect 672264 312060 672316 312112
rect 676036 312060 676088 312112
rect 660948 311992 661000 312044
rect 676220 311992 676272 312044
rect 658372 311788 658424 311840
rect 671160 311788 671212 311840
rect 673368 311652 673420 311704
rect 676036 311652 676088 311704
rect 654140 311244 654192 311296
rect 669412 311244 669464 311296
rect 674748 310972 674800 311024
rect 676036 310972 676088 311024
rect 673184 310836 673236 310888
rect 676036 310836 676088 310888
rect 655428 310428 655480 310480
rect 673276 310428 673328 310480
rect 676036 310428 676088 310480
rect 673092 310020 673144 310072
rect 676036 310020 676088 310072
rect 671160 309612 671212 309664
rect 671896 309612 671948 309664
rect 676036 309612 676088 309664
rect 674196 309136 674248 309188
rect 676036 309136 676088 309188
rect 673552 308048 673604 308100
rect 676036 308048 676088 308100
rect 673460 306484 673512 306536
rect 675944 306484 675996 306536
rect 674472 306416 674524 306468
rect 676036 306416 676088 306468
rect 673920 306348 673972 306400
rect 676128 306348 676180 306400
rect 674656 306008 674708 306060
rect 676036 306008 676088 306060
rect 673644 305056 673696 305108
rect 676128 305056 676180 305108
rect 673736 304648 673788 304700
rect 676128 304648 676180 304700
rect 673828 303832 673880 303884
rect 675852 303832 675904 303884
rect 674012 303764 674064 303816
rect 675944 303764 675996 303816
rect 674564 303696 674616 303748
rect 676128 303696 676180 303748
rect 41512 301588 41564 301640
rect 49148 301588 49200 301640
rect 675208 300976 675260 301028
rect 675484 300976 675536 301028
rect 41788 300908 41840 300960
rect 51172 300908 51224 300960
rect 673092 300840 673144 300892
rect 678980 300840 679032 300892
rect 655612 298256 655664 298308
rect 669596 298256 669648 298308
rect 675760 296148 675812 296200
rect 675760 295944 675812 295996
rect 675208 295060 675260 295112
rect 675392 295060 675444 295112
rect 674196 294516 674248 294568
rect 675392 294516 675444 294568
rect 674472 292884 674524 292936
rect 675392 292884 675444 292936
rect 674656 292272 674708 292324
rect 675392 292272 675444 292324
rect 41788 292000 41840 292052
rect 43352 292000 43404 292052
rect 41788 291592 41840 291644
rect 43536 291592 43588 291644
rect 41880 291116 41932 291168
rect 42708 291116 42760 291168
rect 674564 291048 674616 291100
rect 675392 291048 675444 291100
rect 41788 289824 41840 289876
rect 43168 289824 43220 289876
rect 673920 288532 673972 288584
rect 675392 288532 675444 288584
rect 674012 287920 674064 287972
rect 675392 287920 675444 287972
rect 673736 287172 673788 287224
rect 675484 287172 675536 287224
rect 673828 286560 673880 286612
rect 675392 286560 675444 286612
rect 32680 285744 32732 285796
rect 42800 285744 42852 285796
rect 32864 285676 32916 285728
rect 42984 285676 43036 285728
rect 32772 285608 32824 285660
rect 42892 285608 42944 285660
rect 673644 285540 673696 285592
rect 675484 285540 675536 285592
rect 655336 284724 655388 284776
rect 670516 284724 670568 284776
rect 673552 283704 673604 283756
rect 675484 283704 675536 283756
rect 42156 283568 42208 283620
rect 42708 283568 42760 283620
rect 42432 283296 42484 283348
rect 42708 283296 42760 283348
rect 673460 281868 673512 281920
rect 675392 281868 675444 281920
rect 42156 281732 42208 281784
rect 42800 281732 42852 281784
rect 42156 281052 42208 281104
rect 49056 281052 49108 281104
rect 42156 279828 42208 279880
rect 43076 279828 43128 279880
rect 42064 278604 42116 278656
rect 43168 278604 43220 278656
rect 46480 278536 46532 278588
rect 672816 278536 672868 278588
rect 46572 278468 46624 278520
rect 670240 278468 670292 278520
rect 46756 278400 46808 278452
rect 670424 278400 670476 278452
rect 62580 278332 62632 278384
rect 670148 278332 670200 278384
rect 62764 278264 62816 278316
rect 668768 278264 668820 278316
rect 62948 278196 63000 278248
rect 670332 278196 670384 278248
rect 62396 278128 62448 278180
rect 669688 278128 669740 278180
rect 63132 278060 63184 278112
rect 669780 278060 669832 278112
rect 63224 277992 63276 278044
rect 669872 277992 669924 278044
rect 63316 277924 63368 277976
rect 669964 277924 670016 277976
rect 42156 277856 42208 277908
rect 43260 277856 43312 277908
rect 42156 277380 42208 277432
rect 43536 277380 43588 277432
rect 42064 276700 42116 276752
rect 42984 276700 43036 276752
rect 345112 275952 345164 276004
rect 471336 275952 471388 276004
rect 343732 275884 343784 275936
rect 467840 275884 467892 275936
rect 349068 275816 349120 275868
rect 482008 275816 482060 275868
rect 350356 275748 350408 275800
rect 485504 275748 485556 275800
rect 354404 275680 354456 275732
rect 496176 275680 496228 275732
rect 355784 275612 355836 275664
rect 499764 275612 499816 275664
rect 358452 275544 358504 275596
rect 506848 275544 506900 275596
rect 361120 275476 361172 275528
rect 513932 275476 513984 275528
rect 364064 275408 364116 275460
rect 521016 275408 521068 275460
rect 366456 275340 366508 275392
rect 528100 275340 528152 275392
rect 369124 275272 369176 275324
rect 535184 275272 535236 275324
rect 371792 275204 371844 275256
rect 542268 275204 542320 275256
rect 374920 275136 374972 275188
rect 550548 275136 550600 275188
rect 377588 275068 377640 275120
rect 557632 275068 557684 275120
rect 380256 275000 380308 275052
rect 564716 275000 564768 275052
rect 382924 274932 382976 274984
rect 571800 274932 571852 274984
rect 385592 274864 385644 274916
rect 578884 274864 578936 274916
rect 318892 274796 318944 274848
rect 401600 274796 401652 274848
rect 403900 274796 403952 274848
rect 320180 274728 320232 274780
rect 405188 274728 405240 274780
rect 406568 274728 406620 274780
rect 411444 274796 411496 274848
rect 620284 274796 620336 274848
rect 321008 274660 321060 274712
rect 407488 274660 407540 274712
rect 409236 274660 409288 274712
rect 627368 274728 627420 274780
rect 322848 274592 322900 274644
rect 411076 274592 411128 274644
rect 634452 274660 634504 274712
rect 641628 274592 641680 274644
rect 342536 274524 342588 274576
rect 464252 274524 464304 274576
rect 341064 274456 341116 274508
rect 460664 274456 460716 274508
rect 337108 274388 337160 274440
rect 450084 274388 450136 274440
rect 335728 274320 335780 274372
rect 446496 274320 446548 274372
rect 42156 274252 42208 274304
rect 42892 274252 42944 274304
rect 334348 274252 334400 274304
rect 427084 274252 427136 274304
rect 333428 274184 333480 274236
rect 439412 274184 439464 274236
rect 332140 274116 332192 274168
rect 437020 274116 437072 274168
rect 351828 274048 351880 274100
rect 432328 274048 432380 274100
rect 331680 273980 331732 274032
rect 435916 273980 435968 274032
rect 327724 273912 327776 273964
rect 425244 273912 425296 273964
rect 329104 273844 329156 273896
rect 428832 273844 428884 273896
rect 326804 273776 326856 273828
rect 42064 273708 42116 273760
rect 42708 273708 42760 273760
rect 325424 273708 325476 273760
rect 418160 273708 418212 273760
rect 326344 273640 326396 273692
rect 427084 273776 427136 273828
rect 443000 273776 443052 273828
rect 323676 273572 323728 273624
rect 422852 273640 422904 273692
rect 330392 273504 330444 273556
rect 351828 273504 351880 273556
rect 414572 273504 414624 273556
rect 421656 273504 421708 273556
rect 401140 273436 401192 273488
rect 411444 273436 411496 273488
rect 155684 273096 155736 273148
rect 225880 273164 225932 273216
rect 263232 273164 263284 273216
rect 266728 273164 266780 273216
rect 292120 273164 292172 273216
rect 330668 273164 330720 273216
rect 339500 273164 339552 273216
rect 344836 273164 344888 273216
rect 362776 273164 362828 273216
rect 491484 273164 491536 273216
rect 177856 273096 177908 273148
rect 149796 273028 149848 273080
rect 224408 273028 224460 273080
rect 150992 272960 151044 273012
rect 223948 272960 224000 273012
rect 42156 272892 42208 272944
rect 43352 272892 43404 272944
rect 143908 272892 143960 272944
rect 221280 272892 221332 272944
rect 148600 272824 148652 272876
rect 223212 272824 223264 272876
rect 146208 272756 146260 272808
rect 223028 272756 223080 272808
rect 145012 272688 145064 272740
rect 222200 272688 222252 272740
rect 139124 272620 139176 272672
rect 220360 272620 220412 272672
rect 136824 272552 136876 272604
rect 218612 272552 218664 272604
rect 137928 272484 137980 272536
rect 219440 272484 219492 272536
rect 132040 272416 132092 272468
rect 217692 272416 217744 272468
rect 129648 272348 129700 272400
rect 215668 272348 215720 272400
rect 124956 272280 125008 272332
rect 215024 272280 215076 272332
rect 117872 272212 117924 272264
rect 205548 272212 205600 272264
rect 264428 273096 264480 273148
rect 267188 273096 267240 273148
rect 292580 273096 292632 273148
rect 331864 273096 331916 273148
rect 331956 273096 332008 273148
rect 337752 273096 337804 273148
rect 355324 273096 355376 273148
rect 243176 273028 243228 273080
rect 259184 273028 259236 273080
rect 260932 273028 260984 273080
rect 265808 273028 265860 273080
rect 293408 273028 293460 273080
rect 334164 273028 334216 273080
rect 358820 273028 358872 273080
rect 498568 273096 498620 273148
rect 293868 272960 293920 273012
rect 335360 272960 335412 273012
rect 344008 272960 344060 273012
rect 362592 272960 362644 273012
rect 363144 273028 363196 273080
rect 497372 273028 497424 273080
rect 498844 273028 498896 273080
rect 617984 273028 618036 273080
rect 504456 272960 504508 273012
rect 239588 272892 239640 272944
rect 257804 272892 257856 272944
rect 304908 272892 304960 272944
rect 332508 272892 332560 272944
rect 357992 272892 358044 272944
rect 505652 272892 505704 272944
rect 236092 272824 236144 272876
rect 256424 272824 256476 272876
rect 307852 272824 307904 272876
rect 348424 272824 348476 272876
rect 354864 272824 354916 272876
rect 362868 272824 362920 272876
rect 234896 272756 234948 272808
rect 256056 272756 256108 272808
rect 300768 272756 300820 272808
rect 353116 272756 353168 272808
rect 360660 272756 360712 272808
rect 512736 272824 512788 272876
rect 363236 272756 363288 272808
rect 511540 272756 511592 272808
rect 511632 272756 511684 272808
rect 610808 272756 610860 272808
rect 237288 272688 237340 272740
rect 257160 272688 257212 272740
rect 296076 272688 296128 272740
rect 341340 272688 341392 272740
rect 344928 272688 344980 272740
rect 300676 272620 300728 272672
rect 351920 272620 351972 272672
rect 353024 272620 353076 272672
rect 362776 272620 362828 272672
rect 470140 272688 470192 272740
rect 471980 272688 472032 272740
rect 625068 272688 625120 272740
rect 363144 272620 363196 272672
rect 518624 272620 518676 272672
rect 232504 272552 232556 272604
rect 255136 272552 255188 272604
rect 301412 272552 301464 272604
rect 355508 272552 355560 272604
rect 368204 272552 368256 272604
rect 532792 272552 532844 272604
rect 295248 272484 295300 272536
rect 338948 272484 339000 272536
rect 342812 272484 342864 272536
rect 465448 272484 465500 272536
rect 466276 272484 466328 272536
rect 632152 272484 632204 272536
rect 230204 272416 230256 272468
rect 254216 272416 254268 272468
rect 301872 272416 301924 272468
rect 356704 272416 356756 272468
rect 360568 272416 360620 272468
rect 363236 272416 363288 272468
rect 373172 272416 373224 272468
rect 545856 272416 545908 272468
rect 303528 272348 303580 272400
rect 360200 272348 360252 272400
rect 376668 272348 376720 272400
rect 555240 272348 555292 272400
rect 295064 272280 295116 272332
rect 331956 272280 332008 272332
rect 332508 272280 332560 272332
rect 346032 272280 346084 272332
rect 351828 272280 351880 272332
rect 458364 272280 458416 272332
rect 459468 272280 459520 272332
rect 639236 272280 639288 272332
rect 227076 272212 227128 272264
rect 303344 272212 303396 272264
rect 359004 272212 359056 272264
rect 382004 272212 382056 272264
rect 569500 272212 569552 272264
rect 93032 272144 93084 272196
rect 184940 272144 184992 272196
rect 188804 272144 188856 272196
rect 234804 272144 234856 272196
rect 238484 272144 238536 272196
rect 257252 272144 257304 272196
rect 306288 272144 306340 272196
rect 367284 272144 367336 272196
rect 384672 272144 384724 272196
rect 576584 272144 576636 272196
rect 104900 272076 104952 272128
rect 202696 272076 202748 272128
rect 205364 272076 205416 272128
rect 240140 272076 240192 272128
rect 308956 272076 309008 272128
rect 374368 272076 374420 272128
rect 387340 272076 387392 272128
rect 583668 272076 583720 272128
rect 89536 272008 89588 272060
rect 178040 272008 178092 272060
rect 178132 272008 178184 272060
rect 197268 272008 197320 272060
rect 199476 272008 199528 272060
rect 242624 272008 242676 272060
rect 284208 272008 284260 272060
rect 309416 272008 309468 272060
rect 311624 272008 311676 272060
rect 381544 272008 381596 272060
rect 394608 272008 394660 272060
rect 590752 272008 590804 272060
rect 75276 271940 75328 271992
rect 195428 271940 195480 271992
rect 201776 271940 201828 271992
rect 243544 271940 243596 271992
rect 66996 271872 67048 271924
rect 192484 271872 192536 271924
rect 65892 271804 65944 271856
rect 192116 271804 192168 271856
rect 120264 271736 120316 271788
rect 156788 271736 156840 271788
rect 156880 271736 156932 271788
rect 177856 271736 177908 271788
rect 177948 271736 178000 271788
rect 194508 271736 194560 271788
rect 130844 271668 130896 271720
rect 197176 271804 197228 271856
rect 198280 271804 198332 271856
rect 242256 271872 242308 271924
rect 194692 271668 194744 271720
rect 240876 271804 240928 271856
rect 244372 271804 244424 271856
rect 259552 271940 259604 271992
rect 285404 271940 285456 271992
rect 312912 271940 312964 271992
rect 314292 271940 314344 271992
rect 388628 271940 388680 271992
rect 395436 271940 395488 271992
rect 604920 271940 604972 271992
rect 208492 271668 208544 271720
rect 226524 271736 226576 271788
rect 241980 271736 242032 271788
rect 258724 271872 258776 271924
rect 290280 271872 290332 271924
rect 325976 271872 326028 271924
rect 326712 271872 326764 271924
rect 402796 271872 402848 271924
rect 402888 271872 402940 271924
rect 619088 271872 619140 271924
rect 240784 271668 240836 271720
rect 258264 271804 258316 271856
rect 289544 271804 289596 271856
rect 323584 271804 323636 271856
rect 325608 271804 325660 271856
rect 409880 271804 409932 271856
rect 412824 271804 412876 271856
rect 633348 271804 633400 271856
rect 163964 271600 164016 271652
rect 229744 271600 229796 271652
rect 233700 271600 233752 271652
rect 255596 271736 255648 271788
rect 262128 271736 262180 271788
rect 266268 271736 266320 271788
rect 291752 271736 291804 271788
rect 329472 271736 329524 271788
rect 340236 271736 340288 271788
rect 351828 271736 351880 271788
rect 246764 271668 246816 271720
rect 260472 271668 260524 271720
rect 290740 271668 290792 271720
rect 327080 271668 327132 271720
rect 336740 271668 336792 271720
rect 343640 271668 343692 271720
rect 247868 271600 247920 271652
rect 260932 271600 260984 271652
rect 289820 271600 289872 271652
rect 324780 271600 324832 271652
rect 350264 271600 350316 271652
rect 484308 271736 484360 271788
rect 352380 271668 352432 271720
rect 486700 271668 486752 271720
rect 165160 271532 165212 271584
rect 229468 271532 229520 271584
rect 245568 271532 245620 271584
rect 250168 271532 250220 271584
rect 250260 271532 250312 271584
rect 261852 271532 261904 271584
rect 291200 271532 291252 271584
rect 328276 271532 328328 271584
rect 348240 271532 348292 271584
rect 479616 271600 479668 271652
rect 352104 271532 352156 271584
rect 477224 271532 477276 271584
rect 158076 271464 158128 271516
rect 177948 271464 178000 271516
rect 178132 271464 178184 271516
rect 228824 271464 228876 271516
rect 231400 271464 231452 271516
rect 254676 271464 254728 271516
rect 255044 271464 255096 271516
rect 263600 271464 263652 271516
rect 289360 271464 289412 271516
rect 322388 271464 322440 271516
rect 342168 271464 342220 271516
rect 171048 271396 171100 271448
rect 232412 271396 232464 271448
rect 258540 271396 258592 271448
rect 264888 271396 264940 271448
rect 288532 271396 288584 271448
rect 321192 271396 321244 271448
rect 347596 271396 347648 271448
rect 351920 271396 351972 271448
rect 463056 271464 463108 271516
rect 355968 271396 356020 271448
rect 472532 271396 472584 271448
rect 172244 271328 172296 271380
rect 162768 271260 162820 271312
rect 178132 271260 178184 271312
rect 180064 271328 180116 271380
rect 231492 271328 231544 271380
rect 257344 271328 257396 271380
rect 264520 271328 264572 271380
rect 287612 271328 287664 271380
rect 318800 271328 318852 271380
rect 339408 271328 339460 271380
rect 455972 271328 456024 271380
rect 231768 271260 231820 271312
rect 256148 271260 256200 271312
rect 264060 271260 264112 271312
rect 286784 271260 286836 271312
rect 316500 271260 316552 271312
rect 336464 271260 336516 271312
rect 448888 271260 448940 271312
rect 178040 271192 178092 271244
rect 188620 271192 188672 271244
rect 197268 271192 197320 271244
rect 231952 271192 232004 271244
rect 251456 271192 251508 271244
rect 262220 271192 262272 271244
rect 288164 271192 288216 271244
rect 319996 271192 320048 271244
rect 337476 271192 337528 271244
rect 451280 271192 451332 271244
rect 179328 271124 179380 271176
rect 234528 271124 234580 271176
rect 249064 271124 249116 271176
rect 261392 271124 261444 271176
rect 287152 271124 287204 271176
rect 317696 271124 317748 271176
rect 333980 271124 334032 271176
rect 441804 271124 441856 271176
rect 169852 271056 169904 271108
rect 180064 271056 180116 271108
rect 182916 271056 182968 271108
rect 232044 271056 232096 271108
rect 253848 271056 253900 271108
rect 263140 271056 263192 271108
rect 266820 271056 266872 271108
rect 268016 271056 268068 271108
rect 286692 271056 286744 271108
rect 315304 271056 315356 271108
rect 334808 271056 334860 271108
rect 444196 271056 444248 271108
rect 176936 270988 176988 271040
rect 226432 270988 226484 271040
rect 226616 270988 226668 271040
rect 252928 270988 252980 271040
rect 331312 270988 331364 271040
rect 434720 270988 434772 271040
rect 175832 270920 175884 270972
rect 179328 270920 179380 270972
rect 185216 270920 185268 270972
rect 234712 270920 234764 270972
rect 250168 270920 250220 270972
rect 260012 270920 260064 270972
rect 285864 270920 285916 270972
rect 314108 270920 314160 270972
rect 329932 270920 329984 270972
rect 431132 270920 431184 270972
rect 186412 270852 186464 270904
rect 232136 270852 232188 270904
rect 327264 270852 327316 270904
rect 424048 270852 424100 270904
rect 190000 270784 190052 270836
rect 232504 270784 232556 270836
rect 259736 270784 259788 270836
rect 265348 270784 265400 270836
rect 329012 270784 329064 270836
rect 340144 270784 340196 270836
rect 340328 270784 340380 270836
rect 416964 270784 417016 270836
rect 187608 270716 187660 270768
rect 202788 270716 202840 270768
rect 206744 270716 206796 270768
rect 229376 270716 229428 270768
rect 326436 270716 326488 270768
rect 395712 270716 395764 270768
rect 191196 270648 191248 270700
rect 206744 270580 206796 270632
rect 192300 270512 192352 270564
rect 198648 270512 198700 270564
rect 202788 270512 202840 270564
rect 230204 270648 230256 270700
rect 252652 270648 252704 270700
rect 262864 270648 262916 270700
rect 331128 270648 331180 270700
rect 377956 270648 378008 270700
rect 229008 270580 229060 270632
rect 253756 270580 253808 270632
rect 324596 270580 324648 270632
rect 340328 270580 340380 270632
rect 352012 270580 352064 270632
rect 394516 270580 394568 270632
rect 227812 270512 227864 270564
rect 253388 270512 253440 270564
rect 357440 270512 357492 270564
rect 385040 270512 385092 270564
rect 411812 270512 411864 270564
rect 413100 270512 413152 270564
rect 154488 270444 154540 270496
rect 206468 270444 206520 270496
rect 147404 270376 147456 270428
rect 222660 270444 222712 270496
rect 225420 270444 225472 270496
rect 252468 270444 252520 270496
rect 265624 270444 265676 270496
rect 267556 270444 267608 270496
rect 269856 270444 269908 270496
rect 271512 270444 271564 270496
rect 272064 270444 272116 270496
rect 277492 270444 277544 270496
rect 304080 270444 304132 270496
rect 344008 270444 344060 270496
rect 346860 270444 346912 270496
rect 476120 270444 476172 270496
rect 140320 270308 140372 270360
rect 208032 270308 208084 270360
rect 141516 270240 141568 270292
rect 220820 270376 220872 270428
rect 224224 270376 224276 270428
rect 252008 270376 252060 270428
rect 270316 270376 270368 270428
rect 272708 270376 272760 270428
rect 272984 270376 273036 270428
rect 279792 270376 279844 270428
rect 294328 270376 294380 270428
rect 336556 270376 336608 270428
rect 348608 270376 348660 270428
rect 480812 270376 480864 270428
rect 208308 270308 208360 270360
rect 219992 270308 220044 270360
rect 220728 270308 220780 270360
rect 250720 270308 250772 270360
rect 270684 270308 270736 270360
rect 273904 270308 273956 270360
rect 274272 270308 274324 270360
rect 283380 270308 283432 270360
rect 296996 270308 297048 270360
rect 336740 270308 336792 270360
rect 349528 270308 349580 270360
rect 483204 270308 483256 270360
rect 135628 270172 135680 270224
rect 219072 270240 219124 270292
rect 221924 270240 221976 270292
rect 251088 270240 251140 270292
rect 271144 270240 271196 270292
rect 275100 270240 275152 270292
rect 277400 270240 277452 270292
rect 291660 270240 291712 270292
rect 297456 270240 297508 270292
rect 339500 270240 339552 270292
rect 351276 270240 351328 270292
rect 487896 270240 487948 270292
rect 208400 270172 208452 270224
rect 218152 270172 218204 270224
rect 218336 270172 218388 270224
rect 249800 270172 249852 270224
rect 272524 270172 272576 270224
rect 278688 270172 278740 270224
rect 278780 270172 278832 270224
rect 290464 270172 290516 270224
rect 296536 270172 296588 270224
rect 342444 270172 342496 270224
rect 352196 270172 352248 270224
rect 490288 270172 490340 270224
rect 133236 270104 133288 270156
rect 134432 270036 134484 270088
rect 208216 270036 208268 270088
rect 215944 270104 215996 270156
rect 248880 270104 248932 270156
rect 273720 270104 273772 270156
rect 280988 270104 281040 270156
rect 217324 270036 217376 270088
rect 223120 270036 223172 270088
rect 251548 270036 251600 270088
rect 271604 270036 271656 270088
rect 276296 270036 276348 270088
rect 278688 270036 278740 270088
rect 295156 270104 295208 270156
rect 298284 270104 298336 270156
rect 347228 270104 347280 270156
rect 350908 270104 350960 270156
rect 352380 270104 352432 270156
rect 353576 270104 353628 270156
rect 493784 270104 493836 270156
rect 126152 269968 126204 270020
rect 119068 269900 119120 269952
rect 211896 269900 211948 269952
rect 213644 269968 213696 270020
rect 248052 269968 248104 270020
rect 278320 269968 278372 270020
rect 294052 270036 294104 270088
rect 299204 270036 299256 270088
rect 349620 270036 349672 270088
rect 281540 269968 281592 270020
rect 292856 269968 292908 270020
rect 345480 269968 345532 270020
rect 355968 270036 356020 270088
rect 356244 270036 356296 270088
rect 500868 270036 500920 270088
rect 351736 269968 351788 270020
rect 363788 269968 363840 270020
rect 364708 269968 364760 270020
rect 214656 269900 214708 269952
rect 217140 269900 217192 269952
rect 249340 269900 249392 269952
rect 276940 269900 276992 269952
rect 278780 269900 278832 269952
rect 279608 269900 279660 269952
rect 297548 269900 297600 269952
rect 305460 269900 305512 269952
rect 366088 269900 366140 269952
rect 367376 269900 367428 269952
rect 382464 269968 382516 270020
rect 515128 269968 515180 270020
rect 110788 269832 110840 269884
rect 209688 269832 209740 269884
rect 210056 269832 210108 269884
rect 246672 269832 246724 269884
rect 279148 269832 279200 269884
rect 296352 269832 296404 269884
rect 306748 269832 306800 269884
rect 369676 269832 369728 269884
rect 370044 269832 370096 269884
rect 523408 269900 523460 269952
rect 114284 269764 114336 269816
rect 211068 269764 211120 269816
rect 214840 269764 214892 269816
rect 248420 269764 248472 269816
rect 280528 269764 280580 269816
rect 299940 269764 299992 269816
rect 307208 269764 307260 269816
rect 370872 269764 370924 269816
rect 109592 269696 109644 269748
rect 208860 269696 208912 269748
rect 212448 269696 212500 269748
rect 247592 269696 247644 269748
rect 280068 269696 280120 269748
rect 298744 269696 298796 269748
rect 308128 269696 308180 269748
rect 373264 269764 373316 269816
rect 530492 269832 530544 269884
rect 537576 269764 537628 269816
rect 375380 269696 375432 269748
rect 102508 269628 102560 269680
rect 206192 269628 206244 269680
rect 209136 269628 209188 269680
rect 246212 269628 246264 269680
rect 277860 269628 277912 269680
rect 281540 269628 281592 269680
rect 281816 269628 281868 269680
rect 303436 269628 303488 269680
rect 343272 269628 343324 269680
rect 352288 269628 352340 269680
rect 361580 269628 361632 269680
rect 382280 269628 382332 269680
rect 382464 269696 382516 269748
rect 544660 269696 544712 269748
rect 551744 269628 551796 269680
rect 188620 269560 188672 269612
rect 200764 269560 200816 269612
rect 207756 269560 207808 269612
rect 245752 269560 245804 269612
rect 281448 269560 281500 269612
rect 302332 269560 302384 269612
rect 310796 269560 310848 269612
rect 380348 269560 380400 269612
rect 380716 269560 380768 269612
rect 565912 269560 565964 269612
rect 94228 269492 94280 269544
rect 202604 269492 202656 269544
rect 202972 269492 203024 269544
rect 226340 269492 226392 269544
rect 226432 269492 226484 269544
rect 234160 269492 234212 269544
rect 280988 269492 281040 269544
rect 301136 269492 301188 269544
rect 312084 269492 312136 269544
rect 383844 269492 383896 269544
rect 386052 269492 386104 269544
rect 580080 269492 580132 269544
rect 198648 269424 198700 269476
rect 239956 269424 240008 269476
rect 282736 269424 282788 269476
rect 305828 269424 305880 269476
rect 313464 269424 313516 269476
rect 387432 269424 387484 269476
rect 388720 269424 388772 269476
rect 587164 269424 587216 269476
rect 74080 269356 74132 269408
rect 195888 269356 195940 269408
rect 204168 269356 204220 269408
rect 244464 269356 244516 269408
rect 282276 269356 282328 269408
rect 304632 269356 304684 269408
rect 314844 269356 314896 269408
rect 390928 269356 390980 269408
rect 394056 269356 394108 269408
rect 601424 269356 601476 269408
rect 80060 269288 80112 269340
rect 197268 269288 197320 269340
rect 197360 269288 197412 269340
rect 241796 269288 241848 269340
rect 283656 269288 283708 269340
rect 308220 269288 308272 269340
rect 315212 269288 315264 269340
rect 392124 269288 392176 269340
rect 396724 269288 396776 269340
rect 608508 269288 608560 269340
rect 81256 269220 81308 269272
rect 198096 269220 198148 269272
rect 200580 269220 200632 269272
rect 243084 269220 243136 269272
rect 283196 269220 283248 269272
rect 307024 269220 307076 269272
rect 317880 269220 317932 269272
rect 399208 269220 399260 269272
rect 399392 269220 399444 269272
rect 615592 269220 615644 269272
rect 71780 269152 71832 269204
rect 194600 269152 194652 269204
rect 195796 269152 195848 269204
rect 241336 269152 241388 269204
rect 284944 269152 284996 269204
rect 311716 269152 311768 269204
rect 320548 269152 320600 269204
rect 406292 269152 406344 269204
rect 411444 269152 411496 269204
rect 647516 269152 647568 269204
rect 193496 269084 193548 269136
rect 240416 269084 240468 269136
rect 284484 269084 284536 269136
rect 310520 269084 310572 269136
rect 323216 269084 323268 269136
rect 411812 269084 411864 269136
rect 411904 269084 411956 269136
rect 648712 269084 648764 269136
rect 152188 269016 152240 269068
rect 224868 269016 224920 269068
rect 226340 269016 226392 269068
rect 244004 269016 244056 269068
rect 292948 269016 293000 269068
rect 333060 269016 333112 269068
rect 159272 268948 159324 269000
rect 227536 268948 227588 269000
rect 232136 268948 232188 269000
rect 237288 268948 237340 269000
rect 269396 268948 269448 269000
rect 270408 268948 270460 269000
rect 295616 268948 295668 269000
rect 329012 268948 329064 269000
rect 330852 268948 330904 269000
rect 351828 269016 351880 269068
rect 345940 268948 345992 269000
rect 473728 269016 473780 269068
rect 352288 268948 352340 269000
rect 466644 268948 466696 269000
rect 160468 268880 160520 268932
rect 228456 268880 228508 268932
rect 230204 268880 230256 268932
rect 238208 268880 238260 268932
rect 309876 268880 309928 268932
rect 331128 268880 331180 268932
rect 161572 268812 161624 268864
rect 227996 268812 228048 268864
rect 229376 268812 229428 268864
rect 239588 268812 239640 268864
rect 328644 268812 328696 268864
rect 351920 268880 351972 268932
rect 352104 268880 352156 268932
rect 468944 268880 468996 268932
rect 341524 268812 341576 268864
rect 461860 268812 461912 268864
rect 166356 268744 166408 268796
rect 230204 268744 230256 268796
rect 340604 268744 340656 268796
rect 459560 268744 459612 268796
rect 167552 268676 167604 268728
rect 231124 268676 231176 268728
rect 273812 268676 273864 268728
rect 282184 268676 282236 268728
rect 338856 268676 338908 268728
rect 454776 268676 454828 268728
rect 173440 268608 173492 268660
rect 232872 268608 232924 268660
rect 168656 268540 168708 268592
rect 230664 268540 230716 268592
rect 156788 268472 156840 268524
rect 212816 268472 212868 268524
rect 219532 268472 219584 268524
rect 250260 268608 250312 268660
rect 337936 268608 337988 268660
rect 452476 268608 452528 268660
rect 240140 268540 240192 268592
rect 244924 268540 244976 268592
rect 336188 268540 336240 268592
rect 447692 268540 447744 268592
rect 335268 268472 335320 268524
rect 445300 268472 445352 268524
rect 174636 268404 174688 268456
rect 233792 268404 233844 268456
rect 234804 268404 234856 268456
rect 239128 268404 239180 268456
rect 276480 268404 276532 268456
rect 289268 268404 289320 268456
rect 325976 268404 326028 268456
rect 332784 268404 332836 268456
rect 333520 268404 333572 268456
rect 440608 268404 440660 268456
rect 179328 268336 179380 268388
rect 233332 268336 233384 268388
rect 275192 268336 275244 268388
rect 285772 268336 285824 268388
rect 309416 268336 309468 268388
rect 332508 268336 332560 268388
rect 332600 268336 332652 268388
rect 438216 268336 438268 268388
rect 180524 268268 180576 268320
rect 235540 268268 235592 268320
rect 274732 268268 274784 268320
rect 284576 268268 284628 268320
rect 312544 268268 312596 268320
rect 181720 268200 181772 268252
rect 236460 268200 236512 268252
rect 275652 268200 275704 268252
rect 286876 268200 286928 268252
rect 316132 268200 316184 268252
rect 206560 268132 206612 268184
rect 245292 268132 245344 268184
rect 316592 268132 316644 268184
rect 326436 268132 326488 268184
rect 184112 268064 184164 268116
rect 236920 268064 236972 268116
rect 82360 267996 82412 268048
rect 198556 267996 198608 268048
rect 201316 267996 201368 268048
rect 203892 267996 203944 268048
rect 206468 267996 206520 268048
rect 225328 267996 225380 268048
rect 231952 267996 232004 268048
rect 235080 267996 235132 268048
rect 319260 267996 319312 268048
rect 326712 267996 326764 268048
rect 197176 267928 197228 267980
rect 216864 267928 216916 267980
rect 232044 267928 232096 267980
rect 235724 267928 235776 267980
rect 298744 267928 298796 267980
rect 307852 267928 307904 267980
rect 321928 267928 321980 267980
rect 325608 267928 325660 267980
rect 351828 268268 351880 268320
rect 433524 268268 433576 268320
rect 332692 268200 332744 268252
rect 426440 268200 426492 268252
rect 351920 268132 351972 268184
rect 427636 268132 427688 268184
rect 332784 268064 332836 268116
rect 420552 268064 420604 268116
rect 663708 268064 663760 268116
rect 676220 268064 676272 268116
rect 357440 267996 357492 268048
rect 357532 267996 357584 268048
rect 358728 267996 358780 268048
rect 372712 267996 372764 268048
rect 382464 267996 382516 268048
rect 390008 267996 390060 268048
rect 394608 267996 394660 268048
rect 400772 267996 400824 268048
rect 402888 267996 402940 268048
rect 406108 267996 406160 268048
rect 412824 267996 412876 268048
rect 352012 267928 352064 267980
rect 661132 267928 661184 267980
rect 676036 267928 676088 267980
rect 88340 267860 88392 267912
rect 201224 267860 201276 267912
rect 211252 267860 211304 267912
rect 247132 267860 247184 267912
rect 276296 267860 276348 267912
rect 288072 267860 288124 267912
rect 297916 267860 297968 267912
rect 304908 267860 304960 267912
rect 328000 267860 328052 267912
rect 332692 267860 332744 267912
rect 344192 267860 344244 267912
rect 352104 267860 352156 267912
rect 95424 267792 95476 267844
rect 203524 267792 203576 267844
rect 205548 267792 205600 267844
rect 212356 267792 212408 267844
rect 234712 267792 234764 267844
rect 237748 267792 237800 267844
rect 304540 267792 304592 267844
rect 351736 267792 351788 267844
rect 202696 267724 202748 267776
rect 206560 267724 206612 267776
rect 232504 267724 232556 267776
rect 238668 267724 238720 267776
rect 332508 267724 332560 267776
rect 376760 267724 376812 267776
rect 661040 267724 661092 267776
rect 676128 267724 676180 267776
rect 359740 267656 359792 267708
rect 510344 267656 510396 267708
rect 674748 267656 674800 267708
rect 676036 267656 676088 267708
rect 362408 267588 362460 267640
rect 517428 267588 517480 267640
rect 365076 267520 365128 267572
rect 524512 267520 524564 267572
rect 367744 267452 367796 267504
rect 531596 267452 531648 267504
rect 672264 267452 672316 267504
rect 675944 267452 675996 267504
rect 370504 267384 370556 267436
rect 538772 267384 538824 267436
rect 373540 267316 373592 267368
rect 547052 267316 547104 267368
rect 374460 267248 374512 267300
rect 549352 267248 549404 267300
rect 376208 267180 376260 267232
rect 554136 267180 554188 267232
rect 299664 267112 299716 267164
rect 350724 267112 350776 267164
rect 375840 267112 375892 267164
rect 552940 267112 552992 267164
rect 300952 267044 301004 267096
rect 354312 267044 354364 267096
rect 377128 267044 377180 267096
rect 556436 267044 556488 267096
rect 302332 266976 302384 267028
rect 357900 266976 357952 267028
rect 378508 266976 378560 267028
rect 560024 266976 560076 267028
rect 303712 266908 303764 266960
rect 361396 266908 361448 266960
rect 378876 266908 378928 266960
rect 561220 266908 561272 266960
rect 305000 266840 305052 266892
rect 364984 266840 365036 266892
rect 379796 266840 379848 266892
rect 563520 266840 563572 266892
rect 306380 266772 306432 266824
rect 368480 266772 368532 266824
rect 381636 266772 381688 266824
rect 568304 266772 568356 266824
rect 307668 266704 307720 266756
rect 372068 266704 372120 266756
rect 381176 266704 381228 266756
rect 567108 266704 567160 266756
rect 309048 266636 309100 266688
rect 375564 266636 375616 266688
rect 382464 266636 382516 266688
rect 570696 266636 570748 266688
rect 123760 266568 123812 266620
rect 214196 266568 214248 266620
rect 310336 266568 310388 266620
rect 379152 266568 379204 266620
rect 384304 266568 384356 266620
rect 575388 266568 575440 266620
rect 116676 266500 116728 266552
rect 211528 266500 211580 266552
rect 311716 266500 311768 266552
rect 382648 266500 382700 266552
rect 383844 266500 383896 266552
rect 574192 266500 574244 266552
rect 72976 266432 73028 266484
rect 195060 266432 195112 266484
rect 313004 266432 313056 266484
rect 386236 266432 386288 266484
rect 389180 266432 389232 266484
rect 588360 266432 588412 266484
rect 113180 266364 113232 266416
rect 210148 266364 210200 266416
rect 315672 266364 315724 266416
rect 68192 266296 68244 266348
rect 193220 266296 193272 266348
rect 317052 266296 317104 266348
rect 382188 266296 382240 266348
rect 392308 266364 392360 266416
rect 596640 266364 596692 266416
rect 393320 266296 393372 266348
rect 394976 266296 395028 266348
rect 603724 266296 603776 266348
rect 652944 266296 652996 266348
rect 675668 266296 675720 266348
rect 357072 266228 357124 266280
rect 503260 266228 503312 266280
rect 353116 266160 353168 266212
rect 492588 266160 492640 266212
rect 351736 266092 351788 266144
rect 489092 266092 489144 266144
rect 673276 266092 673328 266144
rect 676220 266092 676272 266144
rect 347780 266024 347832 266076
rect 478420 266024 478472 266076
rect 346400 265956 346452 266008
rect 474924 265956 474976 266008
rect 339776 265888 339828 265940
rect 457168 265888 457220 265940
rect 338396 265820 338448 265872
rect 453580 265820 453632 265872
rect 317512 265752 317564 265804
rect 382096 265752 382148 265804
rect 382188 265752 382240 265804
rect 396908 265752 396960 265804
rect 397644 265752 397696 265804
rect 511632 265752 511684 265804
rect 329472 265684 329524 265736
rect 429936 265684 429988 265736
rect 382280 265616 382332 265668
rect 398012 265616 398064 265668
rect 400312 265616 400364 265668
rect 498844 265616 498896 265668
rect 325516 265548 325568 265600
rect 419356 265548 419408 265600
rect 324136 265480 324188 265532
rect 415768 265480 415820 265532
rect 322940 265412 322992 265464
rect 412272 265412 412324 265464
rect 321468 265344 321520 265396
rect 408684 265344 408736 265396
rect 674748 265344 674800 265396
rect 676036 265344 676088 265396
rect 318340 265276 318392 265328
rect 400404 265276 400456 265328
rect 402980 265276 403032 265328
rect 471980 265276 472032 265328
rect 314384 265208 314436 265260
rect 389732 265208 389784 265260
rect 319720 265140 319772 265192
rect 403992 265140 404044 265192
rect 658280 265004 658332 265056
rect 675760 265004 675812 265056
rect 671896 264936 671948 264988
rect 676220 264936 676272 264988
rect 674196 263032 674248 263084
rect 676036 263032 676088 263084
rect 674012 262488 674064 262540
rect 676128 262488 676180 262540
rect 673736 262284 673788 262336
rect 676128 262284 676180 262336
rect 416780 262216 416832 262268
rect 571708 262216 571760 262268
rect 674288 262216 674340 262268
rect 676036 262216 676088 262268
rect 674104 261808 674156 261860
rect 676036 261808 676088 261860
rect 673460 260176 673512 260228
rect 675576 260176 675628 260228
rect 673552 259700 673604 259752
rect 675576 259700 675628 259752
rect 674472 259632 674524 259684
rect 676128 259632 676180 259684
rect 674380 259564 674432 259616
rect 675944 259564 675996 259616
rect 675024 259496 675076 259548
rect 676128 259496 676180 259548
rect 675208 259428 675260 259480
rect 676036 259428 676088 259480
rect 41512 258340 41564 258392
rect 48412 258340 48464 258392
rect 41512 258000 41564 258052
rect 53932 258000 53984 258052
rect 41512 257524 41564 257576
rect 50988 257524 51040 257576
rect 41788 256844 41840 256896
rect 45836 256844 45888 256896
rect 672816 256844 672868 256896
rect 678980 256844 679032 256896
rect 673644 256776 673696 256828
rect 676128 256776 676180 256828
rect 52276 256708 52328 256760
rect 184940 256708 184992 256760
rect 416780 256708 416832 256760
rect 571800 256708 571852 256760
rect 673828 256708 673880 256760
rect 676036 256708 676088 256760
rect 674748 255280 674800 255332
rect 675668 255280 675720 255332
rect 674656 255212 674708 255264
rect 675760 255212 675812 255264
rect 416780 253920 416832 253972
rect 571524 253920 571576 253972
rect 416780 251200 416832 251252
rect 574100 251200 574152 251252
rect 675760 251200 675812 251252
rect 675760 250928 675812 250980
rect 675208 250384 675260 250436
rect 675484 250384 675536 250436
rect 33048 249772 33100 249824
rect 43628 249772 43680 249824
rect 674196 249568 674248 249620
rect 675392 249568 675444 249620
rect 416780 248412 416832 248464
rect 574192 248412 574244 248464
rect 674288 247868 674340 247920
rect 675484 247868 675536 247920
rect 41512 247664 41564 247716
rect 45928 247664 45980 247716
rect 41512 247256 41564 247308
rect 45836 247256 45888 247308
rect 674472 247256 674524 247308
rect 675392 247256 675444 247308
rect 674380 246508 674432 246560
rect 675392 246508 675444 246560
rect 41512 246440 41564 246492
rect 45744 246440 45796 246492
rect 675116 246032 675168 246084
rect 675392 246032 675444 246084
rect 52184 245624 52236 245676
rect 184940 245624 184992 245676
rect 416780 245624 416832 245676
rect 571616 245624 571668 245676
rect 42708 244468 42760 244520
rect 43536 244468 43588 244520
rect 32956 244400 33008 244452
rect 43076 244400 43128 244452
rect 33048 244332 33100 244384
rect 42892 244332 42944 244384
rect 31668 244264 31720 244316
rect 42708 244264 42760 244316
rect 32864 244196 32916 244248
rect 42984 244196 43036 244248
rect 673736 243584 673788 243636
rect 675300 243584 675352 243636
rect 42432 243312 42484 243364
rect 43812 243312 43864 243364
rect 43352 243108 43404 243160
rect 43628 243108 43680 243160
rect 42800 242972 42852 243024
rect 43352 242972 43404 243024
rect 673828 242904 673880 242956
rect 675300 242904 675352 242956
rect 38292 242836 38344 242888
rect 42800 242836 42852 242888
rect 673552 242156 673604 242208
rect 675392 242156 675444 242208
rect 674380 241884 674432 241936
rect 675300 241884 675352 241936
rect 673644 241544 673696 241596
rect 675392 241544 675444 241596
rect 673460 240524 673512 240576
rect 675392 240524 675444 240576
rect 42156 240320 42208 240372
rect 42432 240320 42484 240372
rect 42156 238416 42208 238468
rect 42708 238416 42760 238468
rect 52092 237396 52144 237448
rect 184940 237396 184992 237448
rect 674472 236852 674524 236904
rect 675392 236852 675444 236904
rect 42156 236648 42208 236700
rect 42892 236648 42944 236700
rect 674748 235560 674800 235612
rect 675668 235560 675720 235612
rect 674656 235492 674708 235544
rect 675760 235492 675812 235544
rect 42156 235356 42208 235408
rect 42800 235356 42852 235408
rect 42156 234608 42208 234660
rect 43260 234608 43312 234660
rect 42156 234200 42208 234252
rect 43168 234200 43220 234252
rect 42156 233316 42208 233368
rect 43720 233316 43772 233368
rect 42156 231072 42208 231124
rect 43628 231072 43680 231124
rect 48872 231072 48924 231124
rect 654140 231072 654192 231124
rect 48964 231004 49016 231056
rect 656992 231004 657044 231056
rect 46664 230936 46716 230988
rect 656900 230936 656952 230988
rect 46848 230868 46900 230920
rect 659752 230868 659804 230920
rect 46204 230800 46256 230852
rect 659660 230800 659712 230852
rect 46388 230732 46440 230784
rect 662696 230732 662748 230784
rect 46112 230664 46164 230716
rect 662420 230664 662472 230716
rect 45928 230596 45980 230648
rect 662512 230596 662564 230648
rect 42156 230528 42208 230580
rect 43076 230528 43128 230580
rect 45836 230528 45888 230580
rect 662604 230528 662656 230580
rect 45744 230460 45796 230512
rect 662788 230460 662840 230512
rect 45376 230392 45428 230444
rect 662880 230392 662932 230444
rect 350172 230256 350224 230308
rect 423864 230256 423916 230308
rect 351644 230188 351696 230240
rect 427176 230188 427228 230240
rect 348792 230120 348844 230172
rect 420460 230120 420512 230172
rect 347320 230052 347372 230104
rect 417148 230052 417200 230104
rect 354496 229984 354548 230036
rect 433892 229984 433944 230036
rect 355876 229916 355928 229968
rect 437296 229916 437348 229968
rect 42156 229848 42208 229900
rect 42984 229848 43036 229900
rect 357348 229848 357400 229900
rect 440700 229848 440752 229900
rect 360200 229780 360252 229832
rect 447416 229780 447468 229832
rect 364064 229712 364116 229764
rect 455788 229712 455840 229764
rect 365536 229644 365588 229696
rect 459192 229644 459244 229696
rect 368388 229576 368440 229628
rect 466000 229576 466052 229628
rect 371608 229508 371660 229560
rect 474280 229508 474332 229560
rect 370504 229440 370556 229492
rect 473452 229440 473504 229492
rect 371240 229372 371292 229424
rect 472624 229372 472676 229424
rect 374092 229304 374144 229356
rect 479340 229304 479392 229356
rect 376208 229236 376260 229288
rect 487160 229236 487212 229288
rect 393688 229168 393740 229220
rect 528376 229168 528428 229220
rect 396908 229100 396960 229152
rect 535552 229100 535604 229152
rect 42156 229032 42208 229084
rect 43352 229032 43404 229084
rect 156144 229032 156196 229084
rect 235356 229032 235408 229084
rect 247040 229032 247092 229084
rect 273904 229032 273956 229084
rect 296352 229032 296404 229084
rect 298468 229032 298520 229084
rect 304540 229032 304592 229084
rect 316132 229032 316184 229084
rect 368020 229032 368072 229084
rect 369768 229032 369820 229084
rect 386236 229032 386288 229084
rect 460940 229032 460992 229084
rect 152832 228964 152884 229016
rect 233976 228964 234028 229016
rect 239956 228964 240008 229016
rect 265348 228964 265400 229016
rect 290740 228964 290792 229016
rect 292396 228964 292448 229016
rect 293224 228964 293276 229016
rect 294604 228964 294656 229016
rect 297456 228964 297508 229016
rect 299388 228964 299440 229016
rect 304172 228964 304224 229016
rect 314660 228964 314712 229016
rect 343456 228964 343508 229016
rect 381084 228964 381136 229016
rect 395068 228964 395120 229016
rect 477500 228964 477552 229016
rect 156972 228896 157024 228948
rect 237196 228896 237248 228948
rect 239220 228896 239272 228948
rect 266728 228896 266780 228948
rect 297824 228896 297876 228948
rect 301872 228896 301924 228948
rect 305644 228896 305696 228948
rect 317880 228896 317932 228948
rect 320272 228896 320324 228948
rect 342168 228896 342220 228948
rect 342352 228896 342404 228948
rect 383752 228896 383804 228948
rect 388720 228896 388772 228948
rect 469864 228896 469916 228948
rect 150256 228828 150308 228880
rect 234344 228828 234396 228880
rect 240692 228828 240744 228880
rect 269580 228828 269632 228880
rect 308496 228828 308548 228880
rect 324596 228828 324648 228880
rect 340604 228828 340656 228880
rect 385224 228828 385276 228880
rect 392952 228828 393004 228880
rect 474740 228828 474792 228880
rect 146024 228760 146076 228812
rect 231124 228760 231176 228812
rect 245292 228760 245344 228812
rect 273536 228760 273588 228812
rect 310612 228760 310664 228812
rect 332140 228760 332192 228812
rect 340880 228760 340932 228812
rect 383660 228760 383712 228812
rect 390836 228760 390888 228812
rect 473268 228760 473320 228812
rect 151728 228692 151780 228744
rect 234712 228692 234764 228744
rect 241980 228692 242032 228744
rect 272156 228692 272208 228744
rect 298836 228692 298888 228744
rect 302700 228692 302752 228744
rect 307392 228692 307444 228744
rect 322940 228692 322992 228744
rect 336648 228692 336700 228744
rect 380992 228692 381044 228744
rect 397276 228692 397328 228744
rect 480260 228692 480312 228744
rect 143448 228624 143500 228676
rect 231492 228624 231544 228676
rect 239864 228624 239916 228676
rect 268200 228624 268252 228676
rect 306656 228624 306708 228676
rect 323768 228624 323820 228676
rect 328828 228624 328880 228676
rect 345388 228624 345440 228676
rect 376576 228624 376628 228676
rect 465908 228624 465960 228676
rect 138480 228556 138532 228608
rect 229008 228556 229060 228608
rect 240140 228556 240192 228608
rect 271052 228556 271104 228608
rect 308128 228556 308180 228608
rect 327080 228556 327132 228608
rect 337752 228556 337804 228608
rect 383844 228556 383896 228608
rect 388352 228556 388404 228608
rect 408316 228556 408368 228608
rect 410892 228556 410944 228608
rect 411168 228556 411220 228608
rect 145196 228488 145248 228540
rect 231860 228488 231912 228540
rect 238576 228488 238628 228540
rect 270684 228488 270736 228540
rect 303528 228488 303580 228540
rect 315304 228488 315356 228540
rect 317420 228488 317472 228540
rect 338120 228488 338172 228540
rect 341984 228488 342036 228540
rect 394608 228488 394660 228540
rect 409052 228488 409104 228540
rect 516232 228556 516284 228608
rect 417332 228488 417384 228540
rect 518900 228488 518952 228540
rect 136824 228420 136876 228472
rect 228640 228420 228692 228472
rect 235264 228420 235316 228472
rect 269304 228420 269356 228472
rect 306012 228420 306064 228472
rect 319536 228420 319588 228472
rect 324872 228420 324924 228472
rect 365812 228420 365864 228472
rect 380808 228420 380860 228472
rect 497832 228420 497884 228472
rect 131764 228352 131816 228404
rect 226156 228352 226208 228404
rect 227628 228352 227680 228404
rect 267096 228352 267148 228404
rect 309508 228352 309560 228404
rect 330484 228352 330536 228404
rect 338028 228352 338080 228404
rect 378140 228352 378192 228404
rect 383384 228352 383436 228404
rect 503720 228352 503772 228404
rect 125048 228284 125100 228336
rect 223304 228284 223356 228336
rect 223488 228284 223540 228336
rect 263876 228284 263928 228336
rect 307760 228284 307812 228336
rect 325700 228284 325752 228336
rect 330576 228284 330628 228336
rect 379244 228284 379296 228336
rect 385500 228284 385552 228336
rect 508780 228284 508832 228336
rect 130108 228216 130160 228268
rect 225788 228216 225840 228268
rect 229376 228216 229428 228268
rect 267464 228216 267516 228268
rect 309232 228216 309284 228268
rect 328828 228216 328880 228268
rect 333428 228216 333480 228268
rect 385960 228216 386012 228268
rect 387616 228216 387668 228268
rect 513840 228216 513892 228268
rect 123392 228148 123444 228200
rect 222936 228148 222988 228200
rect 231676 228148 231728 228200
rect 267832 228148 267884 228200
rect 300952 228148 301004 228200
rect 310244 228148 310296 228200
rect 310520 228148 310572 228200
rect 329656 228148 329708 228200
rect 339132 228148 339184 228200
rect 391848 228148 391900 228200
rect 399392 228148 399444 228200
rect 541624 228148 541676 228200
rect 108212 228080 108264 228132
rect 216128 228080 216180 228132
rect 216680 228080 216732 228132
rect 261024 228080 261076 228132
rect 308864 228080 308916 228132
rect 326252 228080 326304 228132
rect 334900 228080 334952 228132
rect 389088 228080 389140 228132
rect 407212 228080 407264 228132
rect 417332 228080 417384 228132
rect 78772 228012 78824 228064
rect 202604 228012 202656 228064
rect 209688 228012 209740 228064
rect 258172 228012 258224 228064
rect 259368 228012 259420 228064
rect 276020 228012 276072 228064
rect 311716 228012 311768 228064
rect 332968 228012 333020 228064
rect 336280 228012 336332 228064
rect 388996 228012 389048 228064
rect 400496 228012 400548 228064
rect 544108 228080 544160 228132
rect 417516 228012 417568 228064
rect 545212 228012 545264 228064
rect 65340 227944 65392 227996
rect 196900 227944 196952 227996
rect 199016 227944 199068 227996
rect 254308 227944 254360 227996
rect 254400 227944 254452 227996
rect 275652 227944 275704 227996
rect 302792 227944 302844 227996
rect 311164 227944 311216 227996
rect 311348 227944 311400 227996
rect 331312 227944 331364 227996
rect 342720 227944 342772 227996
rect 395160 227944 395212 227996
rect 402612 227944 402664 227996
rect 549260 227944 549312 227996
rect 77944 227876 77996 227928
rect 203064 227876 203116 227928
rect 203248 227876 203300 227928
rect 255320 227876 255372 227928
rect 257252 227876 257304 227928
rect 277492 227876 277544 227928
rect 301688 227876 301740 227928
rect 309416 227876 309468 227928
rect 312728 227876 312780 227928
rect 334716 227876 334768 227928
rect 338396 227876 338448 227928
rect 395252 227876 395304 227928
rect 404728 227876 404780 227928
rect 554228 227876 554280 227928
rect 72056 227808 72108 227860
rect 199752 227808 199804 227860
rect 204076 227808 204128 227860
rect 257160 227808 257212 227860
rect 261484 227808 261536 227860
rect 278872 227808 278924 227860
rect 303804 227808 303856 227860
rect 317420 227808 317472 227860
rect 318800 227808 318852 227860
rect 64512 227740 64564 227792
rect 197636 227740 197688 227792
rect 197728 227740 197780 227792
rect 254032 227740 254084 227792
rect 254216 227740 254268 227792
rect 277124 227740 277176 227792
rect 304908 227740 304960 227792
rect 318708 227740 318760 227792
rect 341248 227808 341300 227860
rect 397644 227808 397696 227860
rect 406844 227808 406896 227860
rect 559288 227808 559340 227860
rect 339776 227740 339828 227792
rect 345940 227740 345992 227792
rect 408224 227740 408276 227792
rect 409328 227740 409380 227792
rect 565452 227740 565504 227792
rect 52736 227672 52788 227724
rect 192944 227672 192996 227724
rect 193036 227672 193088 227724
rect 251824 227672 251876 227724
rect 252008 227672 252060 227724
rect 276388 227672 276440 227724
rect 312084 227672 312136 227724
rect 335544 227672 335596 227724
rect 341616 227672 341668 227724
rect 402152 227672 402204 227724
rect 410432 227672 410484 227724
rect 567936 227672 567988 227724
rect 158720 227604 158772 227656
rect 237564 227604 237616 227656
rect 243636 227604 243688 227656
rect 272432 227604 272484 227656
rect 305276 227604 305328 227656
rect 320364 227604 320416 227656
rect 320640 227604 320692 227656
rect 165436 227536 165488 227588
rect 240416 227536 240468 227588
rect 250352 227536 250404 227588
rect 275284 227536 275336 227588
rect 307024 227536 307076 227588
rect 321192 227536 321244 227588
rect 332048 227604 332100 227656
rect 369676 227604 369728 227656
rect 381912 227604 381964 227656
rect 453672 227604 453724 227656
rect 356060 227536 356112 227588
rect 356612 227536 356664 227588
rect 372896 227536 372948 227588
rect 384028 227536 384080 227588
rect 455420 227536 455472 227588
rect 162768 227468 162820 227520
rect 238208 227468 238260 227520
rect 253664 227468 253716 227520
rect 276756 227468 276808 227520
rect 303160 227468 303212 227520
rect 312820 227468 312872 227520
rect 324504 227468 324556 227520
rect 345296 227468 345348 227520
rect 353024 227468 353076 227520
rect 410984 227468 411036 227520
rect 42064 227400 42116 227452
rect 43536 227400 43588 227452
rect 163688 227400 163740 227452
rect 240048 227400 240100 227452
rect 257344 227400 257396 227452
rect 264612 227400 264664 227452
rect 264704 227400 264756 227452
rect 275008 227400 275060 227452
rect 325976 227400 326028 227452
rect 345112 227400 345164 227452
rect 372988 227400 373040 227452
rect 433156 227400 433208 227452
rect 167092 227332 167144 227384
rect 241428 227332 241480 227384
rect 251272 227332 251324 227384
rect 271420 227332 271472 227384
rect 323124 227332 323176 227384
rect 342812 227332 342864 227384
rect 358728 227332 358780 227384
rect 415308 227332 415360 227384
rect 172152 227264 172204 227316
rect 243268 227264 243320 227316
rect 248512 227264 248564 227316
rect 268568 227264 268620 227316
rect 295248 227264 295300 227316
rect 296812 227264 296864 227316
rect 298744 227264 298796 227316
rect 301044 227264 301096 227316
rect 302424 227264 302476 227316
rect 313648 227264 313700 227316
rect 374828 227264 374880 227316
rect 433248 227264 433300 227316
rect 169576 227196 169628 227248
rect 241060 227196 241112 227248
rect 251180 227196 251232 227248
rect 272800 227196 272852 227248
rect 302056 227196 302108 227248
rect 311992 227196 312044 227248
rect 370136 227196 370188 227248
rect 428372 227196 428424 227248
rect 173624 227128 173676 227180
rect 244280 227128 244332 227180
rect 248604 227128 248656 227180
rect 269948 227128 270000 227180
rect 333060 227128 333112 227180
rect 347780 227128 347832 227180
rect 367284 227128 367336 227180
rect 422300 227128 422352 227180
rect 178868 227060 178920 227112
rect 246120 227060 246172 227112
rect 254124 227060 254176 227112
rect 274272 227060 274324 227112
rect 331680 227060 331732 227112
rect 347872 227060 347924 227112
rect 364432 227060 364484 227112
rect 416780 227060 416832 227112
rect 176384 226992 176436 227044
rect 243912 226992 243964 227044
rect 248420 226992 248472 227044
rect 265716 226992 265768 227044
rect 322020 226992 322072 227044
rect 359096 226992 359148 227044
rect 361580 226992 361632 227044
rect 415492 226992 415544 227044
rect 180524 226924 180576 226976
rect 247132 226924 247184 226976
rect 254308 226924 254360 226976
rect 271788 226924 271840 226976
rect 345204 226924 345256 226976
rect 376668 226924 376720 226976
rect 379060 226924 379112 226976
rect 387524 226924 387576 226976
rect 399024 226924 399076 226976
rect 438860 226924 438912 226976
rect 190368 226856 190420 226908
rect 251456 226856 251508 226908
rect 257804 226856 257856 226908
rect 274640 226856 274692 226908
rect 300676 226856 300728 226908
rect 308588 226856 308640 226908
rect 359832 226856 359884 226908
rect 400220 226856 400272 226908
rect 400772 226856 400824 226908
rect 417516 226856 417568 226908
rect 42156 226788 42208 226840
rect 43904 226788 43956 226840
rect 185584 226788 185636 226840
rect 186412 226720 186464 226772
rect 233884 226720 233936 226772
rect 192944 226652 192996 226704
rect 234068 226788 234120 226840
rect 248236 226788 248288 226840
rect 248696 226788 248748 226840
rect 264704 226788 264756 226840
rect 299572 226788 299624 226840
rect 306932 226788 306984 226840
rect 323492 226788 323544 226840
rect 362408 226788 362460 226840
rect 363052 226788 363104 226840
rect 371516 226788 371568 226840
rect 373356 226788 373408 226840
rect 395988 226788 396040 226840
rect 407580 226788 407632 226840
rect 449624 226856 449676 226908
rect 417700 226788 417752 226840
rect 441620 226788 441672 226840
rect 258448 226720 258500 226772
rect 273168 226720 273220 226772
rect 299204 226720 299256 226772
rect 305276 226720 305328 226772
rect 306380 226720 306432 226772
rect 322020 226720 322072 226772
rect 371976 226720 372028 226772
rect 400404 226720 400456 226772
rect 405464 226720 405516 226772
rect 444564 226720 444616 226772
rect 248972 226652 249024 226704
rect 298100 226652 298152 226704
rect 303620 226652 303672 226704
rect 369584 226652 369636 226704
rect 402980 226652 403032 226704
rect 409696 226652 409748 226704
rect 451188 226652 451240 226704
rect 237288 226584 237340 226636
rect 256792 226584 256844 226636
rect 296720 226584 296772 226636
rect 300216 226584 300268 226636
rect 300308 226584 300360 226636
rect 306380 226584 306432 226636
rect 395804 226584 395856 226636
rect 434628 226584 434680 226636
rect 251088 226516 251140 226568
rect 254032 226516 254084 226568
rect 270316 226516 270368 226568
rect 301320 226516 301372 226568
rect 307760 226516 307812 226568
rect 334532 226516 334584 226568
rect 351920 226516 351972 226568
rect 378692 226516 378744 226568
rect 397460 226516 397512 226568
rect 401140 226516 401192 226568
rect 417700 226516 417752 226568
rect 246304 226448 246356 226500
rect 258540 226448 258592 226500
rect 389364 226448 389416 226500
rect 408408 226448 408460 226500
rect 394792 226380 394844 226432
rect 411168 226380 411220 226432
rect 197912 226312 197964 226364
rect 207940 226312 207992 226364
rect 253940 226312 253992 226364
rect 268936 226312 268988 226364
rect 299940 226312 299992 226364
rect 304356 226312 304408 226364
rect 309876 226312 309928 226364
rect 327908 226312 327960 226364
rect 151084 226244 151136 226296
rect 233608 226244 233660 226296
rect 353760 226244 353812 226296
rect 434812 226244 434864 226296
rect 154488 226176 154540 226228
rect 235080 226176 235132 226228
rect 352288 226176 352340 226228
rect 431408 226176 431460 226228
rect 433248 226176 433300 226228
rect 483020 226176 483072 226228
rect 144368 226108 144420 226160
rect 230756 226108 230808 226160
rect 355140 226108 355192 226160
rect 438124 226108 438176 226160
rect 147772 226040 147824 226092
rect 232228 226040 232280 226092
rect 359464 226040 359516 226092
rect 448244 226040 448296 226092
rect 465908 226040 465960 226092
rect 487804 226040 487856 226092
rect 141056 225972 141108 226024
rect 229100 225972 229152 226024
rect 362316 225972 362368 226024
rect 137652 225904 137704 225956
rect 227904 225904 227956 225956
rect 362684 225904 362736 225956
rect 452660 225904 452712 225956
rect 453672 225972 453724 226024
rect 500684 225972 500736 226024
rect 454960 225904 455012 225956
rect 455420 225904 455472 225956
rect 505744 225904 505796 225956
rect 134248 225836 134300 225888
rect 226524 225836 226576 225888
rect 366916 225836 366968 225888
rect 462504 225836 462556 225888
rect 469864 225836 469916 225888
rect 516416 225904 516468 225956
rect 518900 225904 518952 225956
rect 560392 225904 560444 225956
rect 516232 225836 516284 225888
rect 564348 225836 564400 225888
rect 130936 225768 130988 225820
rect 225052 225768 225104 225820
rect 365168 225768 365220 225820
rect 461676 225768 461728 225820
rect 474740 225768 474792 225820
rect 526444 225768 526496 225820
rect 127532 225700 127584 225752
rect 223672 225700 223724 225752
rect 230112 225700 230164 225752
rect 249616 225700 249668 225752
rect 363696 225700 363748 225752
rect 458456 225700 458508 225752
rect 460940 225700 460992 225752
rect 510712 225700 510764 225752
rect 516140 225700 516192 225752
rect 566832 225700 566884 225752
rect 119160 225632 119212 225684
rect 219716 225632 219768 225684
rect 230296 225632 230348 225684
rect 249984 225632 250036 225684
rect 344468 225632 344520 225684
rect 369584 225632 369636 225684
rect 369768 225632 369820 225684
rect 468392 225632 468444 225684
rect 473268 225632 473320 225684
rect 521660 225632 521712 225684
rect 124128 225564 124180 225616
rect 222200 225564 222252 225616
rect 234528 225564 234580 225616
rect 253848 225564 253900 225616
rect 366548 225564 366600 225616
rect 465080 225564 465132 225616
rect 477500 225564 477552 225616
rect 531504 225564 531556 225616
rect 114100 225496 114152 225548
rect 217968 225496 218020 225548
rect 218060 225496 218112 225548
rect 245384 225496 245436 225548
rect 355508 225496 355560 225548
rect 433524 225496 433576 225548
rect 434628 225496 434680 225548
rect 532792 225496 532844 225548
rect 117504 225428 117556 225480
rect 219348 225428 219400 225480
rect 228456 225428 228508 225480
rect 266452 225428 266504 225480
rect 339868 225428 339920 225480
rect 371240 225428 371292 225480
rect 372620 225428 372672 225480
rect 476028 225428 476080 225480
rect 480260 225428 480312 225480
rect 536564 225428 536616 225480
rect 107384 225360 107436 225412
rect 215116 225360 215168 225412
rect 218428 225360 218480 225412
rect 262128 225360 262180 225412
rect 356980 225360 357032 225412
rect 105728 225292 105780 225344
rect 214012 225292 214064 225344
rect 221740 225292 221792 225344
rect 263600 225292 263652 225344
rect 358360 225292 358412 225344
rect 429016 225292 429068 225344
rect 438860 225360 438912 225412
rect 541440 225360 541492 225412
rect 439044 225292 439096 225344
rect 441620 225292 441672 225344
rect 545764 225292 545816 225344
rect 90548 225224 90600 225276
rect 197912 225224 197964 225276
rect 198188 225224 198240 225276
rect 253572 225224 253624 225276
rect 357992 225224 358044 225276
rect 100668 225156 100720 225208
rect 212264 225156 212316 225208
rect 225144 225156 225196 225208
rect 264980 225156 265032 225208
rect 317788 225156 317840 225208
rect 348976 225156 349028 225208
rect 361212 225156 361264 225208
rect 444564 225224 444616 225276
rect 557448 225224 557500 225276
rect 103980 225088 104032 225140
rect 213644 225088 213696 225140
rect 215024 225088 215076 225140
rect 260748 225088 260800 225140
rect 319168 225088 319220 225140
rect 352380 225088 352432 225140
rect 360844 225088 360896 225140
rect 444104 225088 444156 225140
rect 444840 225156 444892 225208
rect 449624 225156 449676 225208
rect 561220 225156 561272 225208
rect 449072 225088 449124 225140
rect 451188 225088 451240 225140
rect 566004 225088 566056 225140
rect 95608 225020 95660 225072
rect 209504 225020 209556 225072
rect 211712 225020 211764 225072
rect 259276 225020 259328 225072
rect 313464 225020 313516 225072
rect 338856 225020 338908 225072
rect 344100 225020 344152 225072
rect 408684 225020 408736 225072
rect 408960 225020 409012 225072
rect 563704 225020 563756 225072
rect 88892 224952 88944 225004
rect 206836 224952 206888 225004
rect 208308 224952 208360 225004
rect 257896 224952 257948 225004
rect 316316 224952 316368 225004
rect 345664 224952 345716 225004
rect 345848 224952 345900 225004
rect 410800 224952 410852 225004
rect 73712 224884 73764 224936
rect 200856 224884 200908 224936
rect 201408 224884 201460 224936
rect 255044 224884 255096 224936
rect 314936 224884 314988 224936
rect 342444 224884 342496 224936
rect 343732 224884 343784 224936
rect 411168 224952 411220 225004
rect 411536 224952 411588 225004
rect 570236 224952 570288 225004
rect 411076 224884 411128 224936
rect 568580 224884 568632 224936
rect 161204 224816 161256 224868
rect 237932 224816 237984 224868
rect 354128 224816 354180 224868
rect 432236 224816 432288 224868
rect 433156 224816 433208 224868
rect 477776 224816 477828 224868
rect 157800 224748 157852 224800
rect 236460 224748 236512 224800
rect 349436 224748 349488 224800
rect 425060 224748 425112 224800
rect 428372 224748 428424 224800
rect 470968 224748 471020 224800
rect 167920 224680 167972 224732
rect 240784 224680 240836 224732
rect 352656 224680 352708 224732
rect 428924 224680 428976 224732
rect 429016 224680 429068 224732
rect 442356 224680 442408 224732
rect 444104 224680 444156 224732
rect 451556 224680 451608 224732
rect 164608 224612 164660 224664
rect 239312 224612 239364 224664
rect 350908 224612 350960 224664
rect 428004 224612 428056 224664
rect 170956 224544 171008 224596
rect 242164 224544 242216 224596
rect 349804 224544 349856 224596
rect 409696 224544 409748 224596
rect 174636 224476 174688 224528
rect 243360 224476 243412 224528
rect 346584 224476 346636 224528
rect 409604 224476 409656 224528
rect 181352 224408 181404 224460
rect 246488 224408 246540 224460
rect 348056 224408 348108 224460
rect 421288 224544 421340 224596
rect 422300 224544 422352 224596
rect 464252 224544 464304 224596
rect 416780 224476 416832 224528
rect 457444 224476 457496 224528
rect 410800 224408 410852 224460
rect 412088 224408 412140 224460
rect 178040 224340 178092 224392
rect 245016 224340 245068 224392
rect 340236 224340 340288 224392
rect 371148 224340 371200 224392
rect 372896 224340 372948 224392
rect 441620 224340 441672 224392
rect 184756 224272 184808 224324
rect 247868 224272 247920 224324
rect 348424 224272 348476 224324
rect 418804 224272 418856 224324
rect 188160 224204 188212 224256
rect 249340 224204 249392 224256
rect 346952 224204 347004 224256
rect 415400 224204 415452 224256
rect 415492 224204 415544 224256
rect 450728 224204 450780 224256
rect 191472 224136 191524 224188
rect 250720 224136 250772 224188
rect 339500 224136 339552 224188
rect 394792 224136 394844 224188
rect 402980 224136 403032 224188
rect 469220 224136 469272 224188
rect 139308 224068 139360 224120
rect 194876 224068 194928 224120
rect 194968 224068 195020 224120
rect 252192 224068 252244 224120
rect 335176 224068 335228 224120
rect 391020 224068 391072 224120
rect 400220 224068 400272 224120
rect 445668 224068 445720 224120
rect 155868 224000 155920 224052
rect 209596 224000 209648 224052
rect 236828 224000 236880 224052
rect 343088 224000 343140 224052
rect 368112 224000 368164 224052
rect 376668 224000 376720 224052
rect 204904 223932 204956 223984
rect 256424 223932 256476 223984
rect 383752 223932 383804 223984
rect 407856 223932 407908 223984
rect 409696 224000 409748 224052
rect 422300 224000 422352 224052
rect 414572 223932 414624 223984
rect 204260 223864 204312 223916
rect 252468 223864 252520 223916
rect 383660 223864 383712 223916
rect 404452 223864 404504 223916
rect 415308 223864 415360 223916
rect 444380 223864 444432 223916
rect 189724 223796 189776 223848
rect 232504 223796 232556 223848
rect 395160 223796 395212 223848
rect 405740 223796 405792 223848
rect 410984 223796 411036 223848
rect 430580 223796 430632 223848
rect 209412 223728 209464 223780
rect 213092 223728 213144 223780
rect 242532 223728 242584 223780
rect 409604 223728 409656 223780
rect 417976 223728 418028 223780
rect 171048 223660 171100 223712
rect 206560 223660 206612 223712
rect 215208 223660 215260 223712
rect 239680 223660 239732 223712
rect 182180 223592 182232 223644
rect 192300 223592 192352 223644
rect 140136 223524 140188 223576
rect 230020 223592 230072 223644
rect 278688 223524 278740 223576
rect 287796 223524 287848 223576
rect 318432 223524 318484 223576
rect 348148 223592 348200 223644
rect 408224 223592 408276 223644
rect 414020 223592 414072 223644
rect 433524 223592 433576 223644
rect 435640 223592 435692 223644
rect 347780 223524 347832 223576
rect 383660 223524 383712 223576
rect 386512 223524 386564 223576
rect 511356 223524 511408 223576
rect 674564 223524 674616 223576
rect 675852 223524 675904 223576
rect 153660 223456 153712 223508
rect 235724 223456 235776 223508
rect 322388 223456 322440 223508
rect 360752 223456 360804 223508
rect 495808 223456 495860 223508
rect 607588 223456 607640 223508
rect 87144 223388 87196 223440
rect 171048 223388 171100 223440
rect 177212 223388 177264 223440
rect 245752 223388 245804 223440
rect 146944 223320 146996 223372
rect 232872 223320 232924 223372
rect 326988 223320 327040 223372
rect 343640 223388 343692 223440
rect 361764 223388 361816 223440
rect 387248 223388 387300 223440
rect 513380 223388 513432 223440
rect 368296 223320 368348 223372
rect 389732 223320 389784 223372
rect 518900 223320 518952 223372
rect 543556 223320 543608 223372
rect 616420 223320 616472 223372
rect 148600 223252 148652 223304
rect 233240 223252 233292 223304
rect 246672 223252 246724 223304
rect 256056 223252 256108 223304
rect 269672 223252 269724 223304
rect 284576 223252 284628 223304
rect 324136 223252 324188 223304
rect 343456 223252 343508 223304
rect 343548 223252 343600 223304
rect 364340 223252 364392 223304
rect 391940 223252 391992 223304
rect 523960 223252 524012 223304
rect 552020 223252 552072 223304
rect 553676 223252 553728 223304
rect 618260 223252 618312 223304
rect 60280 223184 60332 223236
rect 139308 223184 139360 223236
rect 141884 223184 141936 223236
rect 230388 223184 230440 223236
rect 135168 223116 135220 223168
rect 227536 223116 227588 223168
rect 133420 223048 133472 223100
rect 227168 223048 227220 223100
rect 231032 223048 231084 223100
rect 248512 223184 248564 223236
rect 326344 223184 326396 223236
rect 369124 223184 369176 223236
rect 394056 223184 394108 223236
rect 529020 223184 529072 223236
rect 545764 223184 545816 223236
rect 616880 223184 616932 223236
rect 242808 223116 242860 223168
rect 258448 223116 258500 223168
rect 328460 223116 328512 223168
rect 371700 223116 371752 223168
rect 396172 223116 396224 223168
rect 533988 223116 534040 223168
rect 535552 223116 535604 223168
rect 536104 223116 536156 223168
rect 615040 223116 615092 223168
rect 246764 223048 246816 223100
rect 248420 223048 248472 223100
rect 271420 223048 271472 223100
rect 285680 223048 285732 223100
rect 325608 223048 325660 223100
rect 364984 223048 365036 223100
rect 398656 223048 398708 223100
rect 539876 223048 539928 223100
rect 560208 223048 560260 223100
rect 619180 223048 619232 223100
rect 128360 222980 128412 223032
rect 224684 222980 224736 223032
rect 236092 222980 236144 223032
rect 254032 222980 254084 223032
rect 263784 222980 263836 223032
rect 280988 222980 281040 223032
rect 324044 222980 324096 223032
rect 343548 222980 343600 223032
rect 343640 222980 343692 223032
rect 367468 222980 367520 223032
rect 398288 222980 398340 223032
rect 539048 222980 539100 223032
rect 541440 222980 541492 223032
rect 615960 222980 616012 223032
rect 126704 222912 126756 222964
rect 224040 222912 224092 222964
rect 232688 222912 232740 222964
rect 253940 222912 253992 222964
rect 266360 222912 266412 222964
rect 283196 222912 283248 222964
rect 326620 222912 326672 222964
rect 370872 222912 370924 222964
rect 371240 222912 371292 222964
rect 398564 222912 398616 222964
rect 399760 222912 399812 222964
rect 543096 222912 543148 222964
rect 119988 222844 120040 222896
rect 221464 222844 221516 222896
rect 224316 222844 224368 222896
rect 246764 222844 246816 222896
rect 246856 222844 246908 222896
rect 256700 222844 256752 222896
rect 257068 222844 257120 222896
rect 278136 222844 278188 222896
rect 327356 222844 327408 222896
rect 370044 222844 370096 222896
rect 371148 222844 371200 222896
rect 400404 222844 400456 222896
rect 401876 222844 401928 222896
rect 547512 222844 547564 222896
rect 566004 222844 566056 222896
rect 620560 222844 620612 222896
rect 116584 222776 116636 222828
rect 220084 222776 220136 222828
rect 222568 222776 222620 222828
rect 91376 222708 91428 222760
rect 209044 222708 209096 222760
rect 257344 222776 257396 222828
rect 261300 222776 261352 222828
rect 281356 222776 281408 222828
rect 330208 222776 330260 222828
rect 376760 222776 376812 222828
rect 401508 222776 401560 222828
rect 546684 222776 546736 222828
rect 549352 222776 549404 222828
rect 551100 222776 551152 222828
rect 617800 222776 617852 222828
rect 82176 222640 82228 222692
rect 203984 222640 204036 222692
rect 215852 222640 215904 222692
rect 246856 222640 246908 222692
rect 258908 222708 258960 222760
rect 262956 222708 263008 222760
rect 281724 222708 281776 222760
rect 328092 222708 328144 222760
rect 374184 222708 374236 222760
rect 402244 222708 402296 222760
rect 548340 222708 548392 222760
rect 567936 222708 567988 222760
rect 635464 222708 635516 222760
rect 85488 222572 85540 222624
rect 205456 222572 205508 222624
rect 209136 222572 209188 222624
rect 260472 222640 260524 222692
rect 279608 222640 279660 222692
rect 329472 222640 329524 222692
rect 377588 222640 377640 222692
rect 403624 222640 403676 222692
rect 552020 222640 552072 222692
rect 568580 222640 568632 222692
rect 621020 222640 621072 222692
rect 75368 222504 75420 222556
rect 201132 222504 201184 222556
rect 205824 222504 205876 222556
rect 257528 222572 257580 222624
rect 262128 222572 262180 222624
rect 280712 222572 280764 222624
rect 68652 222436 68704 222488
rect 198280 222436 198332 222488
rect 202420 222436 202472 222488
rect 246672 222436 246724 222488
rect 53564 222368 53616 222420
rect 182180 222368 182232 222420
rect 188988 222368 189040 222420
rect 264612 222504 264664 222556
rect 282828 222504 282880 222556
rect 249524 222436 249576 222488
rect 259368 222436 259420 222488
rect 272248 222436 272300 222488
rect 284944 222572 284996 222624
rect 331588 222572 331640 222624
rect 378416 222572 378468 222624
rect 405832 222572 405884 222624
rect 556712 222572 556764 222624
rect 557448 222572 557500 222624
rect 618720 222572 618772 222624
rect 283196 222504 283248 222556
rect 290280 222504 290332 222556
rect 325240 222436 325292 222488
rect 343640 222504 343692 222556
rect 343732 222504 343784 222556
rect 375380 222504 375432 222556
rect 380992 222504 381044 222556
rect 394700 222504 394752 222556
rect 403992 222504 404044 222556
rect 552112 222504 552164 222556
rect 556528 222504 556580 222556
rect 561220 222504 561272 222556
rect 66168 222300 66220 222352
rect 198648 222300 198700 222352
rect 200764 222300 200816 222352
rect 243728 222300 243780 222352
rect 247868 222368 247920 222420
rect 254400 222368 254452 222420
rect 254584 222368 254636 222420
rect 278504 222368 278556 222420
rect 327724 222368 327776 222420
rect 372620 222436 372672 222488
rect 382280 222436 382332 222488
rect 396264 222436 396316 222488
rect 406476 222436 406528 222488
rect 558828 222436 558880 222488
rect 560208 222436 560260 222488
rect 560392 222436 560444 222488
rect 343548 222368 343600 222420
rect 375932 222368 375984 222420
rect 378140 222368 378192 222420
rect 397736 222368 397788 222420
rect 406200 222368 406252 222420
rect 407948 222368 408000 222420
rect 561772 222368 561824 222420
rect 250076 222300 250128 222352
rect 259368 222300 259420 222352
rect 280344 222300 280396 222352
rect 310980 222300 311032 222352
rect 333980 222300 334032 222352
rect 339776 222300 339828 222352
rect 349804 222300 349856 222352
rect 349896 222300 349948 222352
rect 385132 222300 385184 222352
rect 385224 222300 385276 222352
rect 402980 222300 403032 222352
rect 557540 222300 557592 222352
rect 563704 222436 563756 222488
rect 620100 222436 620152 222488
rect 619640 222368 619692 222420
rect 634084 222300 634136 222352
rect 61936 222232 61988 222284
rect 195428 222232 195480 222284
rect 195704 222232 195756 222284
rect 253204 222232 253256 222284
rect 314200 222232 314252 222284
rect 338028 222232 338080 222284
rect 338120 222232 338172 222284
rect 346492 222232 346544 222284
rect 59176 222164 59228 222216
rect 195796 222164 195848 222216
rect 207480 222164 207532 222216
rect 246304 222164 246356 222216
rect 257896 222164 257948 222216
rect 279976 222164 280028 222216
rect 281448 222164 281500 222216
rect 289912 222164 289964 222216
rect 313096 222164 313148 222216
rect 336740 222164 336792 222216
rect 337384 222164 337436 222216
rect 393596 222232 393648 222284
rect 394608 222232 394660 222284
rect 406200 222232 406252 222284
rect 408132 222232 408184 222284
rect 562876 222232 562928 222284
rect 565452 222232 565504 222284
rect 635004 222232 635056 222284
rect 346676 222164 346728 222216
rect 391940 222164 391992 222216
rect 397644 222164 397696 222216
rect 401968 222164 402020 222216
rect 410892 222164 410944 222216
rect 569316 222164 569368 222216
rect 652852 222164 652904 222216
rect 674656 222164 674708 222216
rect 675760 222164 675812 222216
rect 155316 222096 155368 222148
rect 235816 222096 235868 222148
rect 93768 222028 93820 222080
rect 155868 222028 155920 222080
rect 232596 222028 232648 222080
rect 244648 222096 244700 222148
rect 251088 222096 251140 222148
rect 254216 222096 254268 222148
rect 273076 222096 273128 222148
rect 286048 222096 286100 222148
rect 321652 222096 321704 222148
rect 356520 222096 356572 222148
rect 383016 222096 383068 222148
rect 503536 222096 503588 222148
rect 538864 222096 538916 222148
rect 615500 222096 615552 222148
rect 160376 221960 160428 222012
rect 238300 222028 238352 222080
rect 243728 222028 243780 222080
rect 255688 222028 255740 222080
rect 320916 222028 320968 222080
rect 357348 222028 357400 222080
rect 384396 222028 384448 222080
rect 506296 222028 506348 222080
rect 555056 222028 555108 222080
rect 633164 222028 633216 222080
rect 237748 221960 237800 222012
rect 251272 221960 251324 222012
rect 322756 221960 322808 222012
rect 358268 221960 358320 222012
rect 380532 221960 380584 222012
rect 497372 221960 497424 222012
rect 499028 221960 499080 222012
rect 552112 221960 552164 222012
rect 552848 221960 552900 222012
rect 632704 221960 632756 222012
rect 170496 221892 170548 221944
rect 242900 221892 242952 221944
rect 319812 221892 319864 221944
rect 354036 221892 354088 221944
rect 387524 221892 387576 221944
rect 396172 221892 396224 221944
rect 396264 221892 396316 221944
rect 501236 221892 501288 221944
rect 532792 221892 532844 221944
rect 533436 221892 533488 221944
rect 614580 221892 614632 221944
rect 168748 221824 168800 221876
rect 241796 221824 241848 221876
rect 244464 221824 244516 221876
rect 254124 221824 254176 221876
rect 274732 221824 274784 221876
rect 287060 221824 287112 221876
rect 287152 221824 287204 221876
rect 289268 221824 289320 221876
rect 318064 221824 318116 221876
rect 350632 221824 350684 221876
rect 377956 221824 378008 221876
rect 491300 221824 491352 221876
rect 547512 221824 547564 221876
rect 631784 221824 631836 221876
rect 175464 221756 175516 221808
rect 232596 221756 232648 221808
rect 234344 221756 234396 221808
rect 248604 221756 248656 221808
rect 255412 221756 255464 221808
rect 277860 221756 277912 221808
rect 182088 221688 182140 221740
rect 183928 221620 183980 221672
rect 239404 221688 239456 221740
rect 254308 221688 254360 221740
rect 258816 221688 258868 221740
rect 279240 221688 279292 221740
rect 183100 221552 183152 221604
rect 235632 221552 235684 221604
rect 159548 221484 159600 221536
rect 209596 221484 209648 221536
rect 214196 221484 214248 221536
rect 240968 221620 241020 221672
rect 235908 221552 235960 221604
rect 246580 221620 246632 221672
rect 273904 221620 273956 221672
rect 285312 221756 285364 221808
rect 321284 221756 321336 221808
rect 354864 221756 354916 221808
rect 379428 221756 379480 221808
rect 494520 221756 494572 221808
rect 530676 221756 530728 221808
rect 614028 221756 614080 221808
rect 283932 221688 283984 221740
rect 289544 221688 289596 221740
rect 319904 221688 319956 221740
rect 351460 221688 351512 221740
rect 377680 221688 377732 221740
rect 490288 221688 490340 221740
rect 545212 221688 545264 221740
rect 631324 221688 631376 221740
rect 287060 221620 287112 221672
rect 288532 221620 288584 221672
rect 316684 221620 316736 221672
rect 347320 221620 347372 221672
rect 351920 221620 351972 221672
rect 383752 221620 383804 221672
rect 383844 221620 383896 221672
rect 396080 221620 396132 221672
rect 396172 221620 396224 221672
rect 494152 221620 494204 221672
rect 495808 221620 495860 221672
rect 528376 221620 528428 221672
rect 613568 221620 613620 221672
rect 241152 221552 241204 221604
rect 251180 221552 251232 221604
rect 268844 221552 268896 221604
rect 283564 221552 283616 221604
rect 313832 221552 313884 221604
rect 340604 221552 340656 221604
rect 345388 221552 345440 221604
rect 373356 221552 373408 221604
rect 375472 221552 375524 221604
rect 484400 221552 484452 221604
rect 543096 221552 543148 221604
rect 630864 221552 630916 221604
rect 166264 221416 166316 221468
rect 215208 221416 215260 221468
rect 220084 221416 220136 221468
rect 240968 221484 241020 221536
rect 247500 221484 247552 221536
rect 270408 221484 270460 221536
rect 283840 221484 283892 221536
rect 284852 221484 284904 221536
rect 291384 221484 291436 221536
rect 317052 221484 317104 221536
rect 345020 221484 345072 221536
rect 345112 221484 345164 221536
rect 366640 221484 366692 221536
rect 374460 221484 374512 221536
rect 480996 221484 481048 221536
rect 532700 221484 532752 221536
rect 532976 221484 533028 221536
rect 628932 221484 628984 221536
rect 187240 221348 187292 221400
rect 230296 221348 230348 221400
rect 235540 221348 235592 221400
rect 236920 221348 236972 221400
rect 240692 221348 240744 221400
rect 248788 221416 248840 221468
rect 275560 221416 275612 221468
rect 286416 221416 286468 221468
rect 286508 221416 286560 221468
rect 291752 221416 291804 221468
rect 315212 221416 315264 221468
rect 343916 221416 343968 221468
rect 345296 221416 345348 221468
rect 363236 221416 363288 221468
rect 368756 221416 368808 221468
rect 467564 221416 467616 221468
rect 535460 221416 535512 221468
rect 538036 221416 538088 221468
rect 629944 221416 629996 221468
rect 246948 221348 247000 221400
rect 256240 221348 256292 221400
rect 261484 221348 261536 221400
rect 267188 221348 267240 221400
rect 282460 221348 282512 221400
rect 289084 221348 289136 221400
rect 292120 221348 292172 221400
rect 292396 221348 292448 221400
rect 293500 221348 293552 221400
rect 314568 221348 314620 221400
rect 339684 221348 339736 221400
rect 342812 221348 342864 221400
rect 359924 221348 359976 221400
rect 365904 221348 365956 221400
rect 460940 221348 460992 221400
rect 507952 221348 508004 221400
rect 609888 221348 609940 221400
rect 172980 221280 173032 221332
rect 213092 221280 213144 221332
rect 233516 221280 233568 221332
rect 239864 221280 239916 221332
rect 280620 221280 280672 221332
rect 288164 221280 288216 221332
rect 289728 221280 289780 221332
rect 293132 221280 293184 221332
rect 294972 221280 295024 221332
rect 295616 221280 295668 221332
rect 315948 221280 316000 221332
rect 343088 221280 343140 221332
rect 371516 221280 371568 221332
rect 454132 221280 454184 221332
rect 510712 221280 510764 221332
rect 610348 221280 610400 221332
rect 192300 221212 192352 221264
rect 193036 221212 193088 221264
rect 149428 221144 149480 221196
rect 189724 221144 189776 221196
rect 189816 221144 189868 221196
rect 230112 221212 230164 221264
rect 230204 221212 230256 221264
rect 239220 221212 239272 221264
rect 277308 221212 277360 221264
rect 286692 221212 286744 221264
rect 315580 221212 315632 221264
rect 341432 221212 341484 221264
rect 342168 221212 342220 221264
rect 199936 221144 199988 221196
rect 234528 221144 234580 221196
rect 246120 221144 246172 221196
rect 257804 221144 257856 221196
rect 279792 221144 279844 221196
rect 288900 221144 288952 221196
rect 312360 221144 312412 221196
rect 337200 221144 337252 221196
rect 337292 221144 337344 221196
rect 346676 221144 346728 221196
rect 347872 221212 347924 221264
rect 380072 221212 380124 221264
rect 383752 221212 383804 221264
rect 386788 221212 386840 221264
rect 388996 221212 389048 221264
rect 392676 221212 392728 221264
rect 402152 221212 402204 221264
rect 403624 221212 403676 221264
rect 353300 221144 353352 221196
rect 369584 221144 369636 221196
rect 410340 221144 410392 221196
rect 179696 221076 179748 221128
rect 217968 221076 218020 221128
rect 206652 221008 206704 221060
rect 237288 221076 237340 221128
rect 252928 221076 252980 221128
rect 257252 221076 257304 221128
rect 265532 221076 265584 221128
rect 282092 221076 282144 221128
rect 282368 221076 282420 221128
rect 287152 221076 287204 221128
rect 288256 221076 288308 221128
rect 292764 221076 292816 221128
rect 329840 221076 329892 221128
rect 343732 221076 343784 221128
rect 368112 221076 368164 221128
rect 407028 221076 407080 221128
rect 226800 221008 226852 221060
rect 239956 221008 240008 221060
rect 278136 221008 278188 221060
rect 287060 221008 287112 221060
rect 287336 221008 287388 221060
rect 291016 221008 291068 221060
rect 329196 221008 329248 221060
rect 343548 221008 343600 221060
rect 196532 220940 196584 220992
rect 204260 220940 204312 220992
rect 213368 220940 213420 220992
rect 237104 220940 237156 220992
rect 268016 220940 268068 220992
rect 284208 220940 284260 220992
rect 285680 220940 285732 220992
rect 290648 220940 290700 220992
rect 291568 220940 291620 220992
rect 294236 220940 294288 220992
rect 334164 220940 334216 220992
rect 349896 220940 349948 220992
rect 381176 220940 381228 220992
rect 409512 221008 409564 221060
rect 394792 220940 394844 220992
rect 401140 220940 401192 220992
rect 162032 220872 162084 220924
rect 238944 220872 238996 220924
rect 276480 220872 276532 220924
rect 287428 220872 287480 220924
rect 369676 220872 369728 220924
rect 382648 220872 382700 220924
rect 391848 220872 391900 220924
rect 399484 220872 399536 220924
rect 400496 220872 400548 220924
rect 476856 221212 476908 221264
rect 527548 221212 527600 221264
rect 628012 221212 628064 221264
rect 411904 221144 411956 221196
rect 485228 221144 485280 221196
rect 505744 221144 505796 221196
rect 609428 221144 609480 221196
rect 670056 221144 670108 221196
rect 675944 221144 675996 221196
rect 503536 221076 503588 221128
rect 608968 221076 609020 221128
rect 517244 221008 517296 221060
rect 517888 221008 517940 221060
rect 626172 221008 626224 221060
rect 669044 221008 669096 221060
rect 676036 221008 676088 221060
rect 500684 220940 500736 220992
rect 608508 220940 608560 220992
rect 499028 220872 499080 220924
rect 608048 220872 608100 220924
rect 194048 220804 194100 220856
rect 252836 220804 252888 220856
rect 385408 220804 385460 220856
rect 507952 220804 508004 220856
rect 548340 220804 548392 220856
rect 617340 220804 617392 220856
rect 666468 220804 666520 220856
rect 675668 220804 675720 220856
rect 347688 220736 347740 220788
rect 419724 220736 419776 220788
rect 571708 220736 571760 220788
rect 572720 220736 572772 220788
rect 574100 220736 574152 220788
rect 575204 220736 575256 220788
rect 351276 220668 351328 220720
rect 425520 220668 425572 220720
rect 571616 220668 571668 220720
rect 573548 220668 573600 220720
rect 352012 220600 352064 220652
rect 429752 220600 429804 220652
rect 353392 220532 353444 220584
rect 433340 220532 433392 220584
rect 356244 220464 356296 220516
rect 439780 220464 439832 220516
rect 355048 220396 355100 220448
rect 436468 220396 436520 220448
rect 359372 220328 359424 220380
rect 446588 220328 446640 220380
rect 139308 220260 139360 220312
rect 228272 220260 228324 220312
rect 357716 220260 357768 220312
rect 443184 220260 443236 220312
rect 142712 220192 142764 220244
rect 229652 220192 229704 220244
rect 361948 220192 362000 220244
rect 453304 220192 453356 220244
rect 135996 220124 136048 220176
rect 226616 220124 226668 220176
rect 360568 220124 360620 220176
rect 449900 220124 449952 220176
rect 132408 220056 132460 220108
rect 225420 220056 225472 220108
rect 364800 220056 364852 220108
rect 460020 220056 460072 220108
rect 129280 219988 129332 220040
rect 223948 219988 224000 220040
rect 363420 219988 363472 220040
rect 456616 219988 456668 220040
rect 125876 219920 125928 219972
rect 222292 219920 222344 219972
rect 367652 219920 367704 219972
rect 466736 219920 466788 219972
rect 122472 219852 122524 219904
rect 221096 219852 221148 219904
rect 366272 219852 366324 219904
rect 463700 219852 463752 219904
rect 58624 219784 58676 219836
rect 193772 219784 193824 219836
rect 369308 219784 369360 219836
rect 470140 219784 470192 219836
rect 48504 219716 48556 219768
rect 648528 219716 648580 219768
rect 46020 219648 46072 219700
rect 647148 219648 647200 219700
rect 48596 219580 48648 219632
rect 651288 219580 651340 219632
rect 652760 219580 652812 219632
rect 46296 219512 46348 219564
rect 649908 219512 649960 219564
rect 675576 219512 675628 219564
rect 676036 219512 676088 219564
rect 48688 219444 48740 219496
rect 652760 219444 652812 219496
rect 48780 219376 48832 219428
rect 654140 219376 654192 219428
rect 349160 219308 349212 219360
rect 423036 219308 423088 219360
rect 652668 219308 652720 219360
rect 674840 219308 674892 219360
rect 676036 219308 676088 219360
rect 350540 219240 350592 219292
rect 426348 219240 426400 219292
rect 344836 219172 344888 219224
rect 412916 219172 412968 219224
rect 346308 219104 346360 219156
rect 416228 219104 416280 219156
rect 523408 218492 523460 218544
rect 612648 218492 612700 218544
rect 525800 218424 525852 218476
rect 613108 218424 613160 218476
rect 520832 218356 520884 218408
rect 612188 218356 612240 218408
rect 518716 218288 518768 218340
rect 611728 218288 611780 218340
rect 674104 218288 674156 218340
rect 676036 218288 676088 218340
rect 513472 218220 513524 218272
rect 515772 218220 515824 218272
rect 611268 218220 611320 218272
rect 662604 218220 662656 218272
rect 663984 218220 664036 218272
rect 490288 218152 490340 218204
rect 607128 218152 607180 218204
rect 487160 218084 487212 218136
rect 606668 218084 606720 218136
rect 662604 218084 662656 218136
rect 662880 218084 662932 218136
rect 673460 218084 673512 218136
rect 675944 218084 675996 218136
rect 46940 218016 46992 218068
rect 671160 218016 671212 218068
rect 674380 218016 674432 218068
rect 676036 218016 676088 218068
rect 418160 217948 418212 218000
rect 418620 217948 418672 218000
rect 646964 217948 647016 218000
rect 651656 217948 651708 218000
rect 642732 217880 642784 217932
rect 651380 217880 651432 217932
rect 662512 217880 662564 217932
rect 664444 217880 664496 217932
rect 644112 217812 644164 217864
rect 651472 217812 651524 217864
rect 570696 217404 570748 217456
rect 635924 217404 635976 217456
rect 563060 217336 563112 217388
rect 634544 217336 634596 217388
rect 558184 217268 558236 217320
rect 633624 217268 633676 217320
rect 550640 217200 550692 217252
rect 632244 217200 632296 217252
rect 540520 217132 540572 217184
rect 630404 217132 630456 217184
rect 535368 217064 535420 217116
rect 629484 217064 629536 217116
rect 673644 217064 673696 217116
rect 675944 217064 675996 217116
rect 530308 216996 530360 217048
rect 628472 216996 628524 217048
rect 513472 216928 513524 216980
rect 610808 216928 610860 216980
rect 525432 216860 525484 216912
rect 627552 216860 627604 216912
rect 418528 216792 418580 216844
rect 639696 216792 639748 216844
rect 41420 216724 41472 216776
rect 59268 216724 59320 216776
rect 418436 216724 418488 216776
rect 640616 216724 640668 216776
rect 41604 216656 41656 216708
rect 59452 216656 59504 216708
rect 418620 216656 418672 216708
rect 640156 216656 640208 216708
rect 645584 216656 645636 216708
rect 651564 216656 651616 216708
rect 674196 216656 674248 216708
rect 676036 216656 676088 216708
rect 41512 216588 41564 216640
rect 59360 216588 59412 216640
rect 417884 216588 417936 216640
rect 641076 216588 641128 216640
rect 492496 216520 492548 216572
rect 504456 216520 504508 216572
rect 505008 216520 505060 216572
rect 495992 216452 496044 216504
rect 484216 216384 484268 216436
rect 486700 216384 486752 216436
rect 490104 216384 490156 216436
rect 500224 216384 500276 216436
rect 504456 216384 504508 216436
rect 520372 216520 520424 216572
rect 626632 216520 626684 216572
rect 515220 216452 515272 216504
rect 625712 216452 625764 216504
rect 510252 216384 510304 216436
rect 624792 216384 624844 216436
rect 623872 216316 623924 216368
rect 622492 216248 622544 216300
rect 673552 216248 673604 216300
rect 675944 216248 675996 216300
rect 622032 216180 622084 216232
rect 637856 216112 637908 216164
rect 636384 216044 636436 216096
rect 638316 215976 638368 216028
rect 638776 215908 638828 215960
rect 48228 215840 48280 215892
rect 666192 215840 666244 215892
rect 31668 215772 31720 215824
rect 665272 215772 665324 215824
rect 29184 215704 29236 215756
rect 665732 215704 665784 215756
rect 580172 215568 580224 215620
rect 599768 215568 599820 215620
rect 673920 215432 673972 215484
rect 675852 215432 675904 215484
rect 674288 215364 674340 215416
rect 675944 215364 675996 215416
rect 674472 215296 674524 215348
rect 676036 215296 676088 215348
rect 656900 215092 656952 215144
rect 657912 215092 657964 215144
rect 659660 215092 659712 215144
rect 660764 215092 660816 215144
rect 673828 214616 673880 214668
rect 676036 214616 676088 214668
rect 41512 214208 41564 214260
rect 43444 214208 43496 214260
rect 41420 213868 41472 213920
rect 45560 213868 45612 213920
rect 674012 213800 674064 213852
rect 676036 213800 676088 213852
rect 582288 212576 582340 212628
rect 599952 212576 600004 212628
rect 673736 212576 673788 212628
rect 675944 212576 675996 212628
rect 580264 212508 580316 212560
rect 599860 212508 599912 212560
rect 675208 212508 675260 212560
rect 676036 212508 676088 212560
rect 651288 212440 651340 212492
rect 651380 212440 651432 212492
rect 673184 212032 673236 212084
rect 676036 212032 676088 212084
rect 662420 210876 662472 210928
rect 662696 210876 662748 210928
rect 581644 209856 581696 209908
rect 600044 209856 600096 209908
rect 580540 209788 580592 209840
rect 599124 209788 599176 209840
rect 579712 207068 579764 207120
rect 601516 207068 601568 207120
rect 582288 207000 582340 207052
rect 601424 207000 601476 207052
rect 674564 206116 674616 206168
rect 674840 206116 674892 206168
rect 674840 205980 674892 206032
rect 675392 205980 675444 206032
rect 675760 205980 675812 206032
rect 674656 205708 674708 205760
rect 675208 205708 675260 205760
rect 674380 205504 674432 205556
rect 675300 205504 675352 205556
rect 674380 205368 674432 205420
rect 674472 205164 674524 205216
rect 675300 205164 675352 205216
rect 674104 204552 674156 204604
rect 675300 204552 675352 204604
rect 582288 204280 582340 204332
rect 599952 204280 600004 204332
rect 674196 202716 674248 202768
rect 675484 202716 675536 202768
rect 674288 201832 674340 201884
rect 675392 201832 675444 201884
rect 581092 201560 581144 201612
rect 599952 201560 600004 201612
rect 580724 201492 580776 201544
rect 598940 201492 598992 201544
rect 673920 201492 673972 201544
rect 675392 201492 675444 201544
rect 674012 200676 674064 200728
rect 675392 200676 675444 200728
rect 33048 200200 33100 200252
rect 41880 200200 41932 200252
rect 581092 200064 581144 200116
rect 599952 200064 600004 200116
rect 32956 199996 33008 200048
rect 42524 199996 42576 200048
rect 582288 198704 582340 198756
rect 599124 198704 599176 198756
rect 673644 198364 673696 198416
rect 675392 198364 675444 198416
rect 673736 197548 673788 197600
rect 675484 197548 675536 197600
rect 41880 197412 41932 197464
rect 582288 197344 582340 197396
rect 599860 197344 599912 197396
rect 580724 197276 580776 197328
rect 599952 197276 600004 197328
rect 41880 197140 41932 197192
rect 673828 197004 673880 197056
rect 675392 197004 675444 197056
rect 674656 196528 674708 196580
rect 675392 196528 675444 196580
rect 674472 196392 674524 196444
rect 674656 196392 674708 196444
rect 674840 195304 674892 195356
rect 675392 195304 675444 195356
rect 42156 195236 42208 195288
rect 42524 195236 42576 195288
rect 674380 195168 674432 195220
rect 674840 195168 674892 195220
rect 582196 194624 582248 194676
rect 599124 194624 599176 194676
rect 582288 194556 582340 194608
rect 599952 194556 600004 194608
rect 42064 193468 42116 193520
rect 42892 193468 42944 193520
rect 673460 193468 673512 193520
rect 675392 193468 675444 193520
rect 42156 192176 42208 192228
rect 42800 192176 42852 192228
rect 582196 191836 582248 191888
rect 599124 191836 599176 191888
rect 582288 191768 582340 191820
rect 599952 191768 600004 191820
rect 673552 191632 673604 191684
rect 675392 191632 675444 191684
rect 42064 191428 42116 191480
rect 43076 191428 43128 191480
rect 42156 190952 42208 191004
rect 42984 190952 43036 191004
rect 579804 190408 579856 190460
rect 599860 190408 599912 190460
rect 582196 187620 582248 187672
rect 601608 187620 601660 187672
rect 582288 187552 582340 187604
rect 600964 187552 601016 187604
rect 580264 184832 580316 184884
rect 599952 184832 600004 184884
rect 580908 184764 580960 184816
rect 601424 184764 601476 184816
rect 666652 183880 666704 183932
rect 667020 183880 667072 183932
rect 580632 182112 580684 182164
rect 600044 182112 600096 182164
rect 580540 182044 580592 182096
rect 599860 182044 599912 182096
rect 580724 179324 580776 179376
rect 599952 179324 600004 179376
rect 666836 179324 666888 179376
rect 671436 179324 671488 179376
rect 674748 179324 674800 179376
rect 675852 179324 675904 179376
rect 581092 179256 581144 179308
rect 599768 179256 599820 179308
rect 669504 177080 669556 177132
rect 675944 177080 675996 177132
rect 669136 176944 669188 176996
rect 676036 176944 676088 176996
rect 671436 176876 671488 176928
rect 673276 176876 673328 176928
rect 675944 176876 675996 176928
rect 666928 176808 666980 176860
rect 675760 176808 675812 176860
rect 581000 176672 581052 176724
rect 598940 176672 598992 176724
rect 581460 176604 581512 176656
rect 600044 176604 600096 176656
rect 666744 176604 666796 176656
rect 671344 176604 671396 176656
rect 674840 176604 674892 176656
rect 676036 176604 676088 176656
rect 667020 176536 667072 176588
rect 672172 176536 672224 176588
rect 674656 176332 674708 176384
rect 676036 176332 676088 176384
rect 673368 175992 673420 176044
rect 675944 175992 675996 176044
rect 674564 175516 674616 175568
rect 676036 175516 676088 175568
rect 671344 175244 671396 175296
rect 672264 175244 672316 175296
rect 675944 175244 675996 175296
rect 671896 174428 671948 174480
rect 672172 174428 672224 174480
rect 676036 174428 676088 174480
rect 580816 173884 580868 173936
rect 599952 173884 600004 173936
rect 674104 173884 674156 173936
rect 676036 173884 676088 173936
rect 579712 173816 579764 173868
rect 599860 173816 599912 173868
rect 582288 173748 582340 173800
rect 600136 173748 600188 173800
rect 674656 171640 674708 171692
rect 676036 171640 676088 171692
rect 673736 171300 673788 171352
rect 675944 171300 675996 171352
rect 582196 171164 582248 171216
rect 599952 171164 600004 171216
rect 674564 171164 674616 171216
rect 675944 171164 675996 171216
rect 579896 171096 579948 171148
rect 599860 171096 599912 171148
rect 674840 171096 674892 171148
rect 676036 171096 676088 171148
rect 582012 171028 582064 171080
rect 599768 171028 599820 171080
rect 580540 170960 580592 171012
rect 599676 170960 599728 171012
rect 673460 170008 673512 170060
rect 675944 170008 675996 170060
rect 673644 169192 673696 169244
rect 675944 169192 675996 169244
rect 673828 168716 673880 168768
rect 675944 168716 675996 168768
rect 674748 168648 674800 168700
rect 676036 168648 676088 168700
rect 579712 168512 579764 168564
rect 599952 168512 600004 168564
rect 673552 168512 673604 168564
rect 675852 168512 675904 168564
rect 582104 168444 582156 168496
rect 599032 168444 599084 168496
rect 580172 168376 580224 168428
rect 599768 168376 599820 168428
rect 582288 168308 582340 168360
rect 600320 168308 600372 168360
rect 672172 168240 672224 168292
rect 676036 168240 676088 168292
rect 672356 167832 672408 167884
rect 676036 167832 676088 167884
rect 672080 167016 672132 167068
rect 676036 167016 676088 167068
rect 581276 165724 581328 165776
rect 599860 165724 599912 165776
rect 580356 165656 580408 165708
rect 600044 165656 600096 165708
rect 581920 165588 581972 165640
rect 599952 165588 600004 165640
rect 581828 165520 581880 165572
rect 601148 165520 601200 165572
rect 581460 162936 581512 162988
rect 599860 162936 599912 162988
rect 581000 162868 581052 162920
rect 599952 162868 600004 162920
rect 675760 160964 675812 161016
rect 675760 160760 675812 160812
rect 581184 160216 581236 160268
rect 600044 160216 600096 160268
rect 580908 160148 580960 160200
rect 599952 160148 600004 160200
rect 580540 160080 580592 160132
rect 599860 160080 599912 160132
rect 674840 159876 674892 159928
rect 675392 159876 675444 159928
rect 674104 159332 674156 159384
rect 675484 159332 675536 159384
rect 674656 157700 674708 157752
rect 675484 157700 675536 157752
rect 582012 157496 582064 157548
rect 599952 157496 600004 157548
rect 581092 157428 581144 157480
rect 599860 157428 599912 157480
rect 580816 157360 580868 157412
rect 598940 157360 598992 157412
rect 674564 156884 674616 156936
rect 675392 156884 675444 156936
rect 674748 155660 674800 155712
rect 675484 155660 675536 155712
rect 582196 154640 582248 154692
rect 599952 154640 600004 154692
rect 580724 154572 580776 154624
rect 599860 154572 599912 154624
rect 673736 153348 673788 153400
rect 675392 153348 675444 153400
rect 673828 152532 673880 152584
rect 675392 152532 675444 152584
rect 673644 151988 673696 152040
rect 675392 151988 675444 152040
rect 582288 151920 582340 151972
rect 599860 151920 599912 151972
rect 581828 151852 581880 151904
rect 599952 151852 600004 151904
rect 582104 151784 582156 151836
rect 600044 151784 600096 151836
rect 673552 151376 673604 151428
rect 675392 151376 675444 151428
rect 673460 150356 673512 150408
rect 675392 150356 675444 150408
rect 581920 149200 581972 149252
rect 598940 149200 598992 149252
rect 581552 149132 581604 149184
rect 599860 149132 599912 149184
rect 581368 149064 581420 149116
rect 599952 149064 600004 149116
rect 581460 146344 581512 146396
rect 599952 146344 600004 146396
rect 580632 146276 580684 146328
rect 599860 146276 599912 146328
rect 581736 143692 581788 143744
rect 599952 143692 600004 143744
rect 581276 143624 581328 143676
rect 599860 143624 599912 143676
rect 579712 143556 579764 143608
rect 600044 143556 600096 143608
rect 581644 140904 581696 140956
rect 599860 140904 599912 140956
rect 581000 140836 581052 140888
rect 599952 140836 600004 140888
rect 581184 140768 581236 140820
rect 599308 140768 599360 140820
rect 581092 138116 581144 138168
rect 599952 138116 600004 138168
rect 579804 138048 579856 138100
rect 599860 138048 599912 138100
rect 580080 137980 580132 138032
rect 599768 137980 599820 138032
rect 580172 135328 580224 135380
rect 599952 135328 600004 135380
rect 579896 135260 579948 135312
rect 599860 135260 599912 135312
rect 670516 132880 670568 132932
rect 676220 132880 676272 132932
rect 669596 132744 669648 132796
rect 676128 132744 676180 132796
rect 580908 132608 580960 132660
rect 599860 132608 599912 132660
rect 669412 132608 669464 132660
rect 676036 132608 676088 132660
rect 580264 132540 580316 132592
rect 599952 132540 600004 132592
rect 579988 132472 580040 132524
rect 600044 132472 600096 132524
rect 673276 132268 673328 132320
rect 676220 132268 676272 132320
rect 670792 131656 670844 131708
rect 676036 131656 676088 131708
rect 673368 131452 673420 131504
rect 676220 131452 676272 131504
rect 672448 130840 672500 130892
rect 676036 130840 676088 130892
rect 672264 130636 672316 130688
rect 676220 130636 676272 130688
rect 670884 130024 670936 130076
rect 676036 130024 676088 130076
rect 580724 129888 580776 129940
rect 599768 129888 599820 129940
rect 580356 129820 580408 129872
rect 599860 129820 599912 129872
rect 669320 129820 669372 129872
rect 670792 129820 670844 129872
rect 580540 129752 580592 129804
rect 599952 129752 600004 129804
rect 669228 129752 669280 129804
rect 670884 129752 670936 129804
rect 671896 129684 671948 129736
rect 676036 129684 676088 129736
rect 671988 129412 672040 129464
rect 676220 129412 676272 129464
rect 674380 127712 674432 127764
rect 676036 127712 676088 127764
rect 580816 127032 580868 127084
rect 599952 127032 600004 127084
rect 673644 127032 673696 127084
rect 675944 127032 675996 127084
rect 580448 126964 580500 127016
rect 599860 126964 599912 127016
rect 674564 126964 674616 127016
rect 676036 126964 676088 127016
rect 673552 124516 673604 124568
rect 675668 124516 675720 124568
rect 674748 124448 674800 124500
rect 675944 124448 675996 124500
rect 674472 124380 674524 124432
rect 675852 124380 675904 124432
rect 582288 124312 582340 124364
rect 600044 124312 600096 124364
rect 674656 124312 674708 124364
rect 676128 124312 676180 124364
rect 582012 124244 582064 124296
rect 599952 124244 600004 124296
rect 675116 124244 675168 124296
rect 675944 124244 675996 124296
rect 580632 124176 580684 124228
rect 599768 124176 599820 124228
rect 675208 124176 675260 124228
rect 676036 124176 676088 124228
rect 673828 123224 673880 123276
rect 676036 123224 676088 123276
rect 672908 123088 672960 123140
rect 676036 123088 676088 123140
rect 671620 122680 671672 122732
rect 676036 122680 676088 122732
rect 672264 121864 672316 121916
rect 676036 121864 676088 121916
rect 582104 121592 582156 121644
rect 599860 121592 599912 121644
rect 581920 121524 581972 121576
rect 599952 121524 600004 121576
rect 582196 121456 582248 121508
rect 600044 121456 600096 121508
rect 673736 121456 673788 121508
rect 675944 121456 675996 121508
rect 583668 118804 583720 118856
rect 599952 118804 600004 118856
rect 581828 118736 581880 118788
rect 600044 118736 600096 118788
rect 581552 118668 581604 118720
rect 599860 118668 599912 118720
rect 581736 116016 581788 116068
rect 599860 116016 599912 116068
rect 581276 115948 581328 116000
rect 599952 115948 600004 116000
rect 675760 115744 675812 115796
rect 675760 115540 675812 115592
rect 675208 114996 675260 115048
rect 675392 114996 675444 115048
rect 674380 114180 674432 114232
rect 675392 114180 675444 114232
rect 581644 113228 581696 113280
rect 599952 113228 600004 113280
rect 581460 113160 581512 113212
rect 599860 113160 599912 113212
rect 674564 112344 674616 112396
rect 675392 112344 675444 112396
rect 674748 111868 674800 111920
rect 675392 111868 675444 111920
rect 674656 111120 674708 111172
rect 675392 111120 675444 111172
rect 675116 110644 675168 110696
rect 675392 110644 675444 110696
rect 581368 110508 581420 110560
rect 599952 110508 600004 110560
rect 581000 110440 581052 110492
rect 599768 110440 599820 110492
rect 673644 108196 673696 108248
rect 675484 108196 675536 108248
rect 581184 107652 581236 107704
rect 599952 107652 600004 107704
rect 673828 107516 673880 107568
rect 675392 107516 675444 107568
rect 673552 106972 673604 107024
rect 675392 106972 675444 107024
rect 673736 106360 673788 106412
rect 675392 106360 675444 106412
rect 674472 105136 674524 105188
rect 675484 105136 675536 105188
rect 581092 104864 581144 104916
rect 599952 104864 600004 104916
rect 657728 99764 657780 99816
rect 660902 99764 660954 99816
rect 580908 99356 580960 99408
rect 599952 99356 600004 99408
rect 633072 96568 633124 96620
rect 635280 96568 635332 96620
rect 636292 96568 636344 96620
rect 640984 96568 641036 96620
rect 655980 96568 656032 96620
rect 659568 96568 659620 96620
rect 661868 96568 661920 96620
rect 663064 96568 663116 96620
rect 633808 96500 633860 96552
rect 636384 96500 636436 96552
rect 637028 96500 637080 96552
rect 642364 96500 642416 96552
rect 654692 96500 654744 96552
rect 658280 96500 658332 96552
rect 659108 96500 659160 96552
rect 662512 96500 662564 96552
rect 634452 96432 634504 96484
rect 637580 96432 637632 96484
rect 652024 96432 652076 96484
rect 661960 96432 662012 96484
rect 635740 96364 635792 96416
rect 639880 96364 639932 96416
rect 631140 96024 631192 96076
rect 632106 96024 632158 96076
rect 632428 96024 632480 96076
rect 634406 96024 634458 96076
rect 635096 96024 635148 96076
rect 639006 96024 639058 96076
rect 647516 96024 647568 96076
rect 652760 96024 652812 96076
rect 631784 95888 631836 95940
rect 632980 95888 633032 95940
rect 640064 95888 640116 95940
rect 646044 95888 646096 95940
rect 646780 95888 646832 95940
rect 663340 95888 663392 95940
rect 638868 95820 638920 95872
rect 646228 95820 646280 95872
rect 614764 95752 614816 95804
rect 620008 95616 620060 95668
rect 623504 95616 623556 95668
rect 607220 95548 607272 95600
rect 608968 95548 609020 95600
rect 610256 95548 610308 95600
rect 611544 95548 611596 95600
rect 613016 95548 613068 95600
rect 614856 95548 614908 95600
rect 618260 95548 618312 95600
rect 620100 95548 620152 95600
rect 621204 95548 621256 95600
rect 622676 95548 622728 95600
rect 623780 95548 623832 95600
rect 624608 95548 624660 95600
rect 621296 95480 621348 95532
rect 623320 95480 623372 95532
rect 616144 95412 616196 95464
rect 623228 95412 623280 95464
rect 596180 95344 596232 95396
rect 612924 95344 612976 95396
rect 619364 95344 619416 95396
rect 622124 95344 622176 95396
rect 578148 95276 578200 95328
rect 606392 95276 606444 95328
rect 575664 95208 575716 95260
rect 610348 95208 610400 95260
rect 618720 95208 618772 95260
rect 622676 95208 622728 95260
rect 639604 95752 639656 95804
rect 645952 95752 646004 95804
rect 637488 95684 637540 95736
rect 640524 95684 640576 95736
rect 640892 95684 640944 95736
rect 645860 95684 645912 95736
rect 641628 95616 641680 95668
rect 642824 95616 642876 95668
rect 652668 95616 652720 95668
rect 663800 95616 663852 95668
rect 638316 95548 638368 95600
rect 642272 95548 642324 95600
rect 642916 95548 642968 95600
rect 646412 95548 646464 95600
rect 648160 95548 648212 95600
rect 656992 95548 657044 95600
rect 659200 95548 659252 95600
rect 642732 95480 642784 95532
rect 660580 95480 660632 95532
rect 661408 95480 661460 95532
rect 648620 95344 648672 95396
rect 650736 95344 650788 95396
rect 656624 95344 656676 95396
rect 663156 95344 663208 95396
rect 646136 95276 646188 95328
rect 663432 95276 663484 95328
rect 657084 95208 657136 95260
rect 657912 95208 657964 95260
rect 665180 95140 665232 95192
rect 617432 94936 617484 94988
rect 623320 94936 623372 94988
rect 643100 94936 643152 94988
rect 644848 94936 644900 94988
rect 645952 94868 646004 94920
rect 646228 94868 646280 94920
rect 618076 94800 618128 94852
rect 621940 94800 621992 94852
rect 651840 94800 651892 94852
rect 653404 94800 653456 94852
rect 648712 94664 648764 94716
rect 649448 94664 649500 94716
rect 653312 94664 653364 94716
rect 663708 94664 663760 94716
rect 657268 94596 657320 94648
rect 663524 94596 663576 94648
rect 616788 94528 616840 94580
rect 623136 94528 623188 94580
rect 648896 94528 648948 94580
rect 650092 94528 650144 94580
rect 656900 94528 656952 94580
rect 658556 94528 658608 94580
rect 648068 94460 648120 94512
rect 659844 94460 659896 94512
rect 660396 94460 660448 94512
rect 643560 94188 643612 94240
rect 644204 94052 644256 94104
rect 654048 94052 654100 94104
rect 649356 93984 649408 94036
rect 656900 93984 656952 94036
rect 605748 93848 605800 93900
rect 613568 93848 613620 93900
rect 644756 93848 644808 93900
rect 652944 93848 652996 93900
rect 607312 93780 607364 93832
rect 612188 93780 612240 93832
rect 601700 90992 601752 91044
rect 609980 91060 610032 91112
rect 657084 88816 657136 88868
rect 658004 88816 658056 88868
rect 659476 88816 659528 88868
rect 663616 88816 663668 88868
rect 648896 85484 648948 85536
rect 657728 85484 657780 85536
rect 651840 85416 651892 85468
rect 658832 85416 658884 85468
rect 648712 85348 648764 85400
rect 660672 85348 660724 85400
rect 648620 85280 648672 85332
rect 657176 85280 657228 85332
rect 643100 85212 643152 85264
rect 660120 85212 660172 85264
rect 646412 85144 646464 85196
rect 661408 85144 661460 85196
rect 586428 84600 586480 84652
rect 600320 84600 600372 84652
rect 583852 84532 583904 84584
rect 600504 84532 600556 84584
rect 583760 84464 583812 84516
rect 600688 84464 600740 84516
rect 582288 84396 582340 84448
rect 600228 84396 600280 84448
rect 582196 84328 582248 84380
rect 600412 84328 600464 84380
rect 582012 84260 582064 84312
rect 600596 84260 600648 84312
rect 582104 84192 582156 84244
rect 600780 84192 600832 84244
rect 581920 84124 581972 84176
rect 600872 84124 600924 84176
rect 579620 82628 579672 82680
rect 583668 82628 583720 82680
rect 591948 80792 592000 80844
rect 596180 80792 596232 80844
rect 600228 78480 600280 78532
rect 610348 78480 610400 78532
rect 605840 77800 605892 77852
rect 607312 77800 607364 77852
rect 600044 74468 600096 74520
rect 605748 74468 605800 74520
rect 590660 73108 590712 73160
rect 601608 73108 601660 73160
rect 598940 69028 598992 69080
rect 605840 69028 605892 69080
rect 583668 66240 583720 66292
rect 590660 66240 590712 66292
rect 580540 66172 580592 66224
rect 586428 66172 586480 66224
rect 590660 64812 590712 64864
rect 600044 64812 600096 64864
rect 600320 63520 600372 63572
rect 607496 63520 607548 63572
rect 590752 62092 590804 62144
rect 598940 62092 598992 62144
rect 595076 60800 595128 60852
rect 600228 60800 600280 60852
rect 578240 60664 578292 60716
rect 583668 60732 583720 60784
rect 579620 60460 579672 60512
rect 583760 60460 583812 60512
rect 579620 58624 579672 58676
rect 583852 58624 583904 58676
rect 582564 58080 582616 58132
rect 591948 58080 592000 58132
rect 586428 57944 586480 57996
rect 590660 57944 590712 57996
rect 590752 57944 590804 57996
rect 585140 57876 585192 57928
rect 587900 55224 587952 55276
rect 595076 55224 595128 55276
rect 582564 53592 582616 53644
rect 571340 53524 571392 53576
rect 346860 52368 346912 52420
rect 642916 52368 642968 52420
rect 52092 51008 52144 51060
rect 213828 51008 213880 51060
rect 346492 51008 346544 51060
rect 587992 51008 588044 51060
rect 600320 51008 600372 51060
rect 579620 49784 579672 49836
rect 585140 49784 585192 49836
rect 578608 49716 578660 49768
rect 587900 49716 587952 49768
rect 478144 48424 478196 48476
rect 518808 48424 518860 48476
rect 149244 48356 149296 48408
rect 150256 48356 150308 48408
rect 218060 48356 218112 48408
rect 412640 48356 412692 48408
rect 494060 48356 494112 48408
rect 216128 48288 216180 48340
rect 521844 48288 521896 48340
rect 552020 48288 552072 48340
rect 575664 48288 575716 48340
rect 52276 47064 52328 47116
rect 149244 47064 149296 47116
rect 574836 46928 574888 46980
rect 578240 46928 578292 46980
rect 218060 46860 218112 46912
rect 642640 46860 642692 46912
rect 494060 46792 494112 46844
rect 502248 46792 502300 46844
rect 460664 45840 460716 45892
rect 610256 45840 610308 45892
rect 367100 45772 367152 45824
rect 607404 45772 607456 45824
rect 311900 45704 311952 45756
rect 607588 45704 607640 45756
rect 85120 45636 85172 45688
rect 475660 45636 475712 45688
rect 540888 45636 540940 45688
rect 578608 45636 578660 45688
rect 233148 45568 233200 45620
rect 642824 45568 642876 45620
rect 212448 45500 212500 45552
rect 639328 45500 639380 45552
rect 311900 44140 311952 44192
rect 367100 44140 367152 44192
rect 563612 44140 563664 44192
rect 578148 44140 578200 44192
rect 310428 44072 310480 44124
rect 365168 44072 365220 44124
rect 474464 44072 474516 44124
rect 586428 44072 586480 44124
rect 419724 44004 419776 44056
rect 540888 44004 540940 44056
rect 405556 43936 405608 43988
rect 607220 43936 607272 43988
rect 230940 43868 230992 43920
rect 613016 43868 613068 43920
rect 230388 43800 230440 43852
rect 618260 43800 618312 43852
rect 230756 43732 230808 43784
rect 621204 43732 621256 43784
rect 230848 43664 230900 43716
rect 621296 43664 621348 43716
rect 230572 43596 230624 43648
rect 621480 43596 621532 43648
rect 230480 43528 230532 43580
rect 621112 43528 621164 43580
rect 230664 43460 230716 43512
rect 621388 43460 621440 43512
rect 226248 43392 226300 43444
rect 622492 43392 622544 43444
rect 223488 43324 223540 43376
rect 622308 43324 622360 43376
rect 209688 43256 209740 43308
rect 631876 43256 631928 43308
rect 52184 42848 52236 42900
rect 215300 42848 215352 42900
rect 455420 42236 455472 42288
rect 530676 42304 530728 42356
rect 531044 42304 531096 42356
rect 574836 42236 574888 42288
rect 510620 42168 510672 42220
rect 530676 42168 530728 42220
rect 531044 42168 531096 42220
rect 579528 42168 579580 42220
rect 502248 41828 502300 41880
rect 518532 41828 518584 41880
rect 416688 41760 416740 41812
rect 420736 41760 420788 41812
rect 471704 41760 471756 41812
rect 475568 41760 475620 41812
rect 514024 41760 514076 41812
rect 514852 41760 514904 41812
rect 529664 41760 529716 41812
rect 530216 41760 530268 41812
rect 141792 41488 141844 41540
rect 207020 41488 207072 41540
rect 209688 41488 209740 41540
rect 505652 38632 505704 38684
rect 510620 38632 510672 38684
rect 420736 38564 420788 38616
rect 455420 38564 455472 38616
rect 475660 38564 475712 38616
rect 514024 38564 514076 38616
rect 475568 38496 475620 38548
rect 505652 38496 505704 38548
rect 213184 24760 213236 24812
rect 213828 24760 213880 24812
rect 224592 22992 224644 23044
rect 226248 22992 226300 23044
rect 221740 22516 221792 22568
rect 223488 22516 223540 22568
rect 229376 6468 229428 6520
rect 233148 6468 233200 6520
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366284 1027806 366496 1027834
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366284 1027752 366312 1027806
rect 366468 1027752 366496 1027806
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366284 1024434 366312 1024488
rect 366468 1024434 366496 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366284 1024406 366496 1024434
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 145196 1007480 145248 1007486
rect 154580 1007480 154632 1007486
rect 145196 1007422 145248 1007428
rect 154578 1007448 154580 1007457
rect 154632 1007448 154634 1007457
rect 144828 1005508 144880 1005514
rect 144828 1005450 144880 1005456
rect 109314 1005408 109370 1005417
rect 92500 1005372 92552 1005378
rect 109314 1005343 109316 1005352
rect 92500 1005314 92552 1005320
rect 109368 1005343 109370 1005352
rect 109316 1005314 109368 1005320
rect 92408 999932 92460 999938
rect 92408 999874 92460 999880
rect 92316 999728 92368 999734
rect 92316 999670 92368 999676
rect 92328 999274 92356 999670
rect 92246 999246 92356 999274
rect 92246 995858 92274 999246
rect 92316 999184 92368 999190
rect 92316 999126 92368 999132
rect 86592 995852 86644 995858
rect 86592 995794 86644 995800
rect 88984 995852 89036 995858
rect 88984 995794 89036 995800
rect 92234 995852 92286 995858
rect 92234 995794 92286 995800
rect 86040 995784 86092 995790
rect 85698 995732 86040 995738
rect 86604 995738 86632 995794
rect 87786 995752 87842 995761
rect 85698 995726 86092 995732
rect 85698 995710 86080 995726
rect 86342 995710 86632 995738
rect 87538 995710 87786 995738
rect 88996 995738 89024 995794
rect 92328 995790 92356 999126
rect 92420 995926 92448 999874
rect 92408 995920 92460 995926
rect 92408 995862 92460 995868
rect 91560 995784 91612 995790
rect 88734 995710 89024 995738
rect 89378 995722 89760 995738
rect 91218 995732 91560 995738
rect 91218 995726 91612 995732
rect 92326 995784 92378 995790
rect 92326 995726 92378 995732
rect 89378 995716 89772 995722
rect 89378 995710 89720 995716
rect 87786 995687 87842 995696
rect 91218 995710 91600 995726
rect 89720 995658 89772 995664
rect 77944 995648 77996 995654
rect 77694 995596 77944 995602
rect 85302 995616 85358 995625
rect 77694 995590 77996 995596
rect 77694 995574 77984 995590
rect 85054 995574 85302 995602
rect 85302 995551 85358 995560
rect 82358 995480 82414 995489
rect 77036 993682 77064 995452
rect 78324 993721 78352 995452
rect 80164 993857 80192 995452
rect 80716 995217 80744 995452
rect 81374 995438 81664 995466
rect 82018 995438 82358 995466
rect 81636 995353 81664 995438
rect 82358 995415 82414 995424
rect 81622 995344 81678 995353
rect 81622 995279 81678 995288
rect 80702 995208 80758 995217
rect 80702 995143 80758 995152
rect 84488 994129 84516 995452
rect 84474 994120 84530 994129
rect 84474 994055 84530 994064
rect 80150 993848 80206 993857
rect 80150 993783 80206 993792
rect 78310 993712 78366 993721
rect 77024 993676 77076 993682
rect 78310 993647 78366 993656
rect 77024 993618 77076 993624
rect 92512 990826 92540 1005314
rect 106464 1005168 106516 1005174
rect 106462 1005136 106464 1005145
rect 125600 1005168 125652 1005174
rect 106516 1005136 106518 1005145
rect 125600 1005110 125652 1005116
rect 143814 1005136 143870 1005145
rect 106462 1005071 106518 1005080
rect 108028 1004896 108080 1004902
rect 108026 1004864 108028 1004873
rect 108080 1004864 108082 1004873
rect 108026 1004799 108082 1004808
rect 108854 1004864 108910 1004873
rect 108854 1004799 108856 1004808
rect 108908 1004799 108910 1004808
rect 108856 1004770 108908 1004776
rect 92960 1004760 93012 1004766
rect 105636 1004760 105688 1004766
rect 92960 1004702 93012 1004708
rect 98274 1004728 98330 1004737
rect 92592 999864 92644 999870
rect 92592 999806 92644 999812
rect 92604 995722 92632 999806
rect 92868 999660 92920 999666
rect 92868 999602 92920 999608
rect 92776 999592 92828 999598
rect 92776 999534 92828 999540
rect 92684 999388 92736 999394
rect 92684 999330 92736 999336
rect 92696 995994 92724 999330
rect 92684 995988 92736 995994
rect 92684 995930 92736 995936
rect 92592 995716 92644 995722
rect 92592 995658 92644 995664
rect 92788 995217 92816 999534
rect 92880 995654 92908 999602
rect 92868 995648 92920 995654
rect 92868 995590 92920 995596
rect 92774 995208 92830 995217
rect 92774 995143 92830 995152
rect 89628 990820 89680 990826
rect 89628 990762 89680 990768
rect 92500 990820 92552 990826
rect 92500 990762 92552 990768
rect 73436 989460 73488 989466
rect 73436 989402 73488 989408
rect 45468 988100 45520 988106
rect 45468 988042 45520 988048
rect 42340 972936 42392 972942
rect 42340 972878 42392 972884
rect 41800 968833 41828 969272
rect 41786 968824 41842 968833
rect 41786 968759 41842 968768
rect 42076 967094 42104 967405
rect 42352 967298 42380 972878
rect 42156 967292 42208 967298
rect 42156 967234 42208 967240
rect 42340 967292 42392 967298
rect 42340 967234 42392 967240
rect 42064 967088 42116 967094
rect 42064 967030 42116 967036
rect 42168 966756 42196 967234
rect 42800 967088 42852 967094
rect 42800 967030 42852 967036
rect 41800 965161 41828 965565
rect 41786 965152 41842 965161
rect 41786 965087 41842 965096
rect 42168 964034 42196 964376
rect 42156 964028 42208 964034
rect 42156 963970 42208 963976
rect 41800 963393 41828 963725
rect 41786 963384 41842 963393
rect 41786 963319 41842 963328
rect 42168 962674 42196 963084
rect 42156 962668 42208 962674
rect 42156 962610 42208 962616
rect 42168 962130 42196 962540
rect 42156 962124 42208 962130
rect 42156 962066 42208 962072
rect 42076 959546 42104 960024
rect 42064 959540 42116 959546
rect 42064 959482 42116 959488
rect 42168 958934 42196 959412
rect 42156 958928 42208 958934
rect 42156 958870 42208 958876
rect 42076 958526 42104 958732
rect 42064 958520 42116 958526
rect 42064 958462 42116 958468
rect 42076 957778 42104 958188
rect 42064 957772 42116 957778
rect 42064 957714 42116 957720
rect 42182 956338 42380 956366
rect 42168 955398 42196 955740
rect 42156 955392 42208 955398
rect 42156 955334 42208 955340
rect 42168 955182 42288 955210
rect 42168 955060 42196 955182
rect 41972 950836 42024 950842
rect 41972 950778 42024 950784
rect 35624 949612 35676 949618
rect 35624 949554 35676 949560
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 35636 934153 35664 949554
rect 35716 949544 35768 949550
rect 35716 949486 35768 949492
rect 35806 949512 35862 949521
rect 35728 934561 35756 949486
rect 35806 949447 35862 949456
rect 41512 949476 41564 949482
rect 35820 934969 35848 949447
rect 41512 949418 41564 949424
rect 41524 943945 41552 949418
rect 41510 943936 41566 943945
rect 41510 943871 41566 943880
rect 41786 943120 41842 943129
rect 41786 943055 41788 943064
rect 41840 943055 41842 943064
rect 41788 943026 41840 943032
rect 41788 942744 41840 942750
rect 41786 942712 41788 942721
rect 41840 942712 41842 942721
rect 41786 942647 41842 942656
rect 41878 942304 41934 942313
rect 41878 942239 41934 942248
rect 41788 941520 41840 941526
rect 41786 941488 41788 941497
rect 41840 941488 41842 941497
rect 41786 941423 41842 941432
rect 41788 941384 41840 941390
rect 41788 941326 41840 941332
rect 41694 940536 41750 940545
rect 41694 940471 41750 940480
rect 41708 936562 41736 940471
rect 41800 936601 41828 941326
rect 41892 941254 41920 942239
rect 41984 941905 42012 950778
rect 41970 941896 42026 941905
rect 41970 941831 42026 941840
rect 41880 941248 41932 941254
rect 41880 941190 41932 941196
rect 41878 941080 41934 941089
rect 41878 941015 41934 941024
rect 41786 936592 41842 936601
rect 41154 936556 41206 936562
rect 41154 936498 41206 936504
rect 41696 936556 41748 936562
rect 41786 936527 41842 936536
rect 41696 936498 41748 936504
rect 35806 934960 35862 934969
rect 35806 934895 35862 934904
rect 35714 934552 35770 934561
rect 35714 934487 35770 934496
rect 35622 934144 35678 934153
rect 35622 934079 35678 934088
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 41166 817018 41194 936498
rect 41892 936442 41920 941015
rect 41970 940264 42026 940273
rect 41970 940199 42026 940208
rect 41984 938505 42012 940199
rect 41970 938496 42026 938505
rect 41970 938431 42026 938440
rect 42260 938233 42288 955182
rect 42352 939049 42380 956338
rect 42708 955392 42760 955398
rect 42708 955334 42760 955340
rect 42720 941390 42748 955334
rect 42708 941384 42760 941390
rect 42708 941326 42760 941332
rect 42708 941248 42760 941254
rect 42708 941190 42760 941196
rect 42338 939040 42394 939049
rect 42338 938975 42394 938984
rect 42246 938224 42302 938233
rect 42246 938159 42302 938168
rect 41708 936414 41920 936442
rect 41708 902534 41736 936414
rect 41786 933328 41842 933337
rect 41786 933263 41842 933272
rect 41800 932113 41828 933263
rect 41786 932104 41842 932113
rect 41786 932039 41788 932048
rect 41840 932039 41842 932048
rect 41788 932010 41840 932016
rect 41800 931979 41828 932010
rect 41524 902506 41736 902534
rect 41524 844574 41552 902506
rect 41524 844546 41736 844574
rect 41154 817012 41206 817018
rect 41154 816954 41206 816960
rect 41708 815833 41736 844546
rect 41786 817728 41842 817737
rect 41786 817663 41788 817672
rect 41840 817663 41842 817672
rect 41788 817634 41840 817640
rect 41788 817352 41840 817358
rect 41786 817320 41788 817329
rect 41840 817320 41842 817329
rect 41786 817255 41842 817264
rect 42720 817086 42748 941190
rect 42812 938641 42840 967030
rect 42984 964028 43036 964034
rect 42984 963970 43036 963976
rect 42892 962668 42944 962674
rect 42892 962610 42944 962616
rect 42904 959682 42932 962610
rect 42892 959676 42944 959682
rect 42892 959618 42944 959624
rect 42892 959540 42944 959546
rect 42892 959482 42944 959488
rect 42904 949550 42932 959482
rect 42892 949544 42944 949550
rect 42892 949486 42944 949492
rect 42996 939978 43024 963970
rect 43076 962124 43128 962130
rect 43076 962066 43128 962072
rect 42904 939950 43024 939978
rect 42798 938632 42854 938641
rect 42798 938567 42854 938576
rect 42904 933745 42932 939950
rect 42982 939856 43038 939865
rect 42982 939791 43038 939800
rect 42890 933736 42946 933745
rect 42890 933671 42946 933680
rect 42798 922040 42854 922049
rect 42798 921975 42854 921984
rect 42708 817080 42760 817086
rect 42708 817022 42760 817028
rect 41788 817012 41840 817018
rect 41788 816954 41840 816960
rect 41694 815824 41750 815833
rect 41694 815759 41750 815768
rect 41800 814473 41828 816954
rect 41878 816504 41934 816513
rect 41878 816439 41934 816448
rect 41786 814464 41842 814473
rect 41786 814399 41842 814408
rect 41788 814292 41840 814298
rect 41788 814234 41840 814240
rect 41800 813657 41828 814234
rect 41892 814201 41920 816439
rect 42720 816105 42748 817022
rect 42706 816096 42762 816105
rect 42706 816031 42762 816040
rect 42338 814872 42394 814881
rect 42338 814807 42394 814816
rect 41878 814192 41934 814201
rect 41878 814127 41934 814136
rect 41786 813648 41842 813657
rect 41786 813583 41842 813592
rect 41786 811608 41842 811617
rect 41786 811543 41842 811552
rect 41800 808722 41828 811543
rect 41878 811200 41934 811209
rect 41878 811135 41934 811144
rect 41788 808716 41840 808722
rect 41788 808658 41840 808664
rect 41786 808344 41842 808353
rect 41786 808279 41788 808288
rect 41840 808279 41842 808288
rect 41788 808250 41840 808256
rect 41786 807936 41842 807945
rect 41786 807871 41842 807880
rect 41800 806070 41828 807871
rect 41788 806064 41840 806070
rect 41788 806006 41840 806012
rect 41892 800222 41920 811135
rect 41970 807528 42026 807537
rect 41970 807463 42026 807472
rect 41984 806313 42012 807463
rect 41970 806304 42026 806313
rect 41970 806239 42026 806248
rect 41984 806002 42012 806239
rect 41972 805996 42024 806002
rect 41972 805938 42024 805944
rect 41880 800216 41932 800222
rect 41880 800158 41932 800164
rect 42352 800086 42380 814807
rect 42616 808308 42668 808314
rect 42616 808250 42668 808256
rect 42340 800080 42392 800086
rect 42340 800022 42392 800028
rect 41880 800012 41932 800018
rect 41880 799954 41932 799960
rect 41892 799445 41920 799954
rect 42156 798176 42208 798182
rect 42156 798118 42208 798124
rect 42168 797605 42196 798118
rect 42628 797910 42656 808250
rect 42708 806064 42760 806070
rect 42708 806006 42760 806012
rect 42616 797904 42668 797910
rect 42616 797846 42668 797852
rect 42432 797632 42484 797638
rect 42432 797574 42484 797580
rect 42156 797292 42208 797298
rect 42156 797234 42208 797240
rect 42168 796960 42196 797234
rect 42156 796340 42208 796346
rect 42156 796282 42208 796288
rect 42168 795765 42196 796282
rect 42156 795048 42208 795054
rect 42156 794990 42208 794996
rect 42168 794580 42196 794990
rect 42156 794300 42208 794306
rect 42156 794242 42208 794248
rect 42168 793900 42196 794242
rect 42444 793830 42472 797574
rect 42720 795054 42748 806006
rect 42708 795048 42760 795054
rect 42708 794990 42760 794996
rect 42156 793824 42208 793830
rect 42156 793766 42208 793772
rect 42432 793824 42484 793830
rect 42432 793766 42484 793772
rect 42168 793288 42196 793766
rect 42156 793008 42208 793014
rect 42156 792950 42208 792956
rect 42168 792744 42196 792950
rect 42156 790696 42208 790702
rect 42156 790638 42208 790644
rect 42168 790228 42196 790638
rect 42156 790152 42208 790158
rect 42156 790094 42208 790100
rect 42168 789616 42196 790094
rect 42156 789472 42208 789478
rect 42156 789414 42208 789420
rect 42168 788936 42196 789414
rect 42156 788860 42208 788866
rect 42156 788802 42208 788808
rect 42168 788392 42196 788802
rect 42156 787024 42208 787030
rect 42156 786966 42208 786972
rect 42168 786556 42196 786966
rect 42064 786276 42116 786282
rect 42064 786218 42116 786224
rect 42076 785944 42104 786218
rect 42156 785664 42208 785670
rect 42156 785606 42208 785612
rect 42168 785264 42196 785606
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 41512 774784 41564 774790
rect 41510 774752 41512 774761
rect 41564 774752 41566 774761
rect 41510 774687 41566 774696
rect 41512 774444 41564 774450
rect 41512 774386 41564 774392
rect 41524 774353 41552 774386
rect 41510 774344 41566 774353
rect 41510 774279 41566 774288
rect 41512 773968 41564 773974
rect 41510 773936 41512 773945
rect 41564 773936 41566 773945
rect 41510 773871 41566 773880
rect 42062 773256 42118 773265
rect 42062 773191 42118 773200
rect 42076 772818 42104 773191
rect 42064 772812 42116 772818
rect 42064 772754 42116 772760
rect 41878 767952 41934 767961
rect 41878 767887 41934 767896
rect 41510 764144 41566 764153
rect 41510 764079 41566 764088
rect 41524 762929 41552 764079
rect 41510 762920 41566 762929
rect 41510 762855 41512 762864
rect 41564 762855 41566 762864
rect 41512 762826 41564 762832
rect 41788 760572 41840 760578
rect 41788 760514 41840 760520
rect 41800 757081 41828 760514
rect 41786 757072 41842 757081
rect 41892 757042 41920 767887
rect 41970 766728 42026 766737
rect 41970 766663 42026 766672
rect 41984 757081 42012 766663
rect 42076 757654 42104 772754
rect 42154 772032 42210 772041
rect 42154 771967 42210 771976
rect 42064 757648 42116 757654
rect 42064 757590 42116 757596
rect 42168 757450 42196 771967
rect 42430 769584 42486 769593
rect 42430 769519 42486 769528
rect 42156 757444 42208 757450
rect 42156 757386 42208 757392
rect 41970 757072 42026 757081
rect 41786 757007 41842 757016
rect 41880 757036 41932 757042
rect 41970 757007 42026 757016
rect 41880 756978 41932 756984
rect 41880 756764 41932 756770
rect 41880 756706 41932 756712
rect 41892 756228 41920 756706
rect 42444 755546 42472 769519
rect 42706 767136 42762 767145
rect 42706 767071 42762 767080
rect 42720 757382 42748 767071
rect 42708 757376 42760 757382
rect 42708 757318 42760 757324
rect 42432 755540 42484 755546
rect 42432 755482 42484 755488
rect 42156 755472 42208 755478
rect 42156 755414 42208 755420
rect 42168 755206 42196 755414
rect 42614 755304 42670 755313
rect 42614 755239 42670 755248
rect 42156 755200 42208 755206
rect 42156 755142 42208 755148
rect 42156 754928 42208 754934
rect 42156 754870 42208 754876
rect 42168 754392 42196 754870
rect 41878 754080 41934 754089
rect 41878 754015 41934 754024
rect 41892 753780 41920 754015
rect 42156 753092 42208 753098
rect 42156 753034 42208 753040
rect 42168 752556 42196 753034
rect 42156 751800 42208 751806
rect 42156 751742 42208 751748
rect 42168 751369 42196 751742
rect 42156 751120 42208 751126
rect 42156 751062 42208 751068
rect 42168 750720 42196 751062
rect 42064 750644 42116 750650
rect 42064 750586 42116 750592
rect 42076 750108 42104 750586
rect 42156 749828 42208 749834
rect 42156 749770 42208 749776
rect 42168 749529 42196 749770
rect 42628 749698 42656 755239
rect 42616 749692 42668 749698
rect 42616 749634 42668 749640
rect 42168 746978 42196 747048
rect 42156 746972 42208 746978
rect 42156 746914 42208 746920
rect 42156 746768 42208 746774
rect 42156 746710 42208 746716
rect 42168 746401 42196 746710
rect 42156 746292 42208 746298
rect 42156 746234 42208 746240
rect 42168 745756 42196 746234
rect 42156 745476 42208 745482
rect 42156 745418 42208 745424
rect 42168 745212 42196 745418
rect 42156 743776 42208 743782
rect 42156 743718 42208 743724
rect 42168 743376 42196 743718
rect 42156 743096 42208 743102
rect 42156 743038 42208 743044
rect 42168 742696 42196 743038
rect 42156 742620 42208 742626
rect 42156 742562 42208 742568
rect 42168 742084 42196 742562
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 39762 731096 39818 731105
rect 39762 731031 39818 731040
rect 39776 730289 39804 731031
rect 39762 730280 39818 730289
rect 39762 730215 39818 730224
rect 39776 728249 39804 730215
rect 42812 730153 42840 921975
rect 42996 902534 43024 939791
rect 43088 937417 43116 962066
rect 43628 959676 43680 959682
rect 43628 959618 43680 959624
rect 43260 958928 43312 958934
rect 43260 958870 43312 958876
rect 43168 957772 43220 957778
rect 43168 957714 43220 957720
rect 43180 937825 43208 957714
rect 43166 937816 43222 937825
rect 43166 937751 43222 937760
rect 43074 937408 43130 937417
rect 43074 937343 43130 937352
rect 43272 935785 43300 958870
rect 43352 958520 43404 958526
rect 43352 958462 43404 958468
rect 43364 936193 43392 958462
rect 43640 949618 43668 959618
rect 43628 949612 43680 949618
rect 43628 949554 43680 949560
rect 43350 936184 43406 936193
rect 43350 936119 43406 936128
rect 43258 935776 43314 935785
rect 43258 935711 43314 935720
rect 43810 927208 43866 927217
rect 43810 927143 43866 927152
rect 42904 902506 43024 902534
rect 42904 814298 42932 902506
rect 43718 815280 43774 815289
rect 43718 815215 43774 815224
rect 42892 814292 42944 814298
rect 42892 814234 42944 814240
rect 43350 814056 43406 814065
rect 43350 813991 43406 814000
rect 42982 813240 43038 813249
rect 42982 813175 43038 813184
rect 42890 812832 42946 812841
rect 42890 812767 42946 812776
rect 42904 798182 42932 812767
rect 42892 798176 42944 798182
rect 42892 798118 42944 798124
rect 42892 798040 42944 798046
rect 42892 797982 42944 797988
rect 42904 772886 42932 797982
rect 42996 787030 43024 813175
rect 43166 810384 43222 810393
rect 43166 810319 43222 810328
rect 43074 809568 43130 809577
rect 43074 809503 43130 809512
rect 43088 796346 43116 809503
rect 43076 796340 43128 796346
rect 43076 796282 43128 796288
rect 43076 796204 43128 796210
rect 43076 796146 43128 796152
rect 42984 787024 43036 787030
rect 42984 786966 43036 786972
rect 43088 786282 43116 796146
rect 43180 789478 43208 810319
rect 43258 809160 43314 809169
rect 43258 809095 43314 809104
rect 43272 794306 43300 809095
rect 43364 798046 43392 813991
rect 43442 812424 43498 812433
rect 43442 812359 43498 812368
rect 43352 798040 43404 798046
rect 43352 797982 43404 797988
rect 43352 797904 43404 797910
rect 43352 797846 43404 797852
rect 43260 794300 43312 794306
rect 43260 794242 43312 794248
rect 43168 789472 43220 789478
rect 43168 789414 43220 789420
rect 43076 786276 43128 786282
rect 43076 786218 43128 786224
rect 42892 772880 42944 772886
rect 42892 772822 42944 772828
rect 42904 770409 42932 772822
rect 43364 772449 43392 797846
rect 43456 785670 43484 812359
rect 43534 812016 43590 812025
rect 43534 811951 43590 811960
rect 43548 788866 43576 811951
rect 43626 808752 43682 808761
rect 43626 808687 43682 808696
rect 43640 790702 43668 808687
rect 43732 797910 43760 815215
rect 43720 797904 43772 797910
rect 43720 797846 43772 797852
rect 43720 797768 43772 797774
rect 43720 797710 43772 797716
rect 43628 790696 43680 790702
rect 43628 790638 43680 790644
rect 43536 788860 43588 788866
rect 43536 788802 43588 788808
rect 43444 785664 43496 785670
rect 43444 785606 43496 785612
rect 43350 772440 43406 772449
rect 43350 772375 43406 772384
rect 43732 771225 43760 797710
rect 43718 771216 43774 771225
rect 43718 771151 43774 771160
rect 42890 770400 42946 770409
rect 42890 770335 42946 770344
rect 43258 769176 43314 769185
rect 43258 769111 43314 769120
rect 43166 768360 43222 768369
rect 43166 768295 43222 768304
rect 43074 766320 43130 766329
rect 43074 766255 43130 766264
rect 42890 764688 42946 764697
rect 42890 764623 42946 764632
rect 42904 751806 42932 764623
rect 42984 757648 43036 757654
rect 42984 757590 43036 757596
rect 42892 751800 42944 751806
rect 42892 751742 42944 751748
rect 42798 730144 42854 730153
rect 42798 730079 42854 730088
rect 42996 729745 43024 757590
rect 43088 753098 43116 766255
rect 43180 766034 43208 768295
rect 43272 766154 43300 769111
rect 43442 768768 43498 768777
rect 43442 768703 43498 768712
rect 43260 766148 43312 766154
rect 43260 766090 43312 766096
rect 43180 766006 43392 766034
rect 43258 765912 43314 765921
rect 43258 765847 43314 765856
rect 43166 765096 43222 765105
rect 43166 765031 43222 765040
rect 43076 753092 43128 753098
rect 43076 753034 43128 753040
rect 43074 752992 43130 753001
rect 43074 752927 43130 752936
rect 42982 729736 43038 729745
rect 41512 729700 41564 729706
rect 42982 729671 43038 729680
rect 41512 729642 41564 729648
rect 41524 729473 41552 729642
rect 43088 729570 43116 752927
rect 43180 750650 43208 765031
rect 43272 751126 43300 765847
rect 43260 751120 43312 751126
rect 43260 751062 43312 751068
rect 43260 750984 43312 750990
rect 43260 750926 43312 750932
rect 43168 750644 43220 750650
rect 43168 750586 43220 750592
rect 43168 750508 43220 750514
rect 43168 750450 43220 750456
rect 43180 746298 43208 750450
rect 43272 746978 43300 750926
rect 43364 749834 43392 766006
rect 43456 757602 43484 768703
rect 43626 767544 43682 767553
rect 43626 767479 43682 767488
rect 43640 766426 43668 767479
rect 43824 767294 43852 927143
rect 43902 810792 43958 810801
rect 43902 810727 43958 810736
rect 43916 800222 43944 810727
rect 43994 809976 44050 809985
rect 43994 809911 44050 809920
rect 43904 800216 43956 800222
rect 43904 800158 43956 800164
rect 43904 800080 43956 800086
rect 43904 800022 43956 800028
rect 43916 798182 43944 800022
rect 43904 798176 43956 798182
rect 43904 798118 43956 798124
rect 43904 798040 43956 798046
rect 43904 797982 43956 797988
rect 43916 793014 43944 797982
rect 43904 793008 43956 793014
rect 43904 792950 43956 792956
rect 44008 790158 44036 809911
rect 44088 808716 44140 808722
rect 44088 808658 44140 808664
rect 44100 800306 44128 808658
rect 44272 800488 44324 800494
rect 44272 800430 44324 800436
rect 44100 800278 44220 800306
rect 44088 800216 44140 800222
rect 44088 800158 44140 800164
rect 44100 796210 44128 800158
rect 44192 798046 44220 800278
rect 44180 798040 44232 798046
rect 44180 797982 44232 797988
rect 44284 797298 44312 800430
rect 44272 797292 44324 797298
rect 44272 797234 44324 797240
rect 44088 796204 44140 796210
rect 44088 796146 44140 796152
rect 43996 790152 44048 790158
rect 43996 790094 44048 790100
rect 44086 770808 44142 770817
rect 44086 770743 44142 770752
rect 43994 769992 44050 770001
rect 43994 769927 44050 769936
rect 43732 767266 43852 767294
rect 43628 766420 43680 766426
rect 43628 766362 43680 766368
rect 43628 766284 43680 766290
rect 43628 766226 43680 766232
rect 43640 757761 43668 766226
rect 43732 765626 43760 767266
rect 43904 766420 43956 766426
rect 43904 766362 43956 766368
rect 43732 765598 43852 765626
rect 43718 765504 43774 765513
rect 43718 765439 43774 765448
rect 43626 757752 43682 757761
rect 43626 757687 43682 757696
rect 43456 757574 43668 757602
rect 43444 757512 43496 757518
rect 43444 757454 43496 757460
rect 43352 749828 43404 749834
rect 43352 749770 43404 749776
rect 43352 749692 43404 749698
rect 43352 749634 43404 749640
rect 43260 746972 43312 746978
rect 43260 746914 43312 746920
rect 43364 746774 43392 749634
rect 43352 746768 43404 746774
rect 43352 746710 43404 746716
rect 43168 746292 43220 746298
rect 43168 746234 43220 746240
rect 43456 743782 43484 757454
rect 43536 757444 43588 757450
rect 43536 757386 43588 757392
rect 43444 743776 43496 743782
rect 43444 743718 43496 743724
rect 43548 729706 43576 757386
rect 43640 745482 43668 757574
rect 43732 750990 43760 765439
rect 43720 750984 43772 750990
rect 43720 750926 43772 750932
rect 43628 745476 43680 745482
rect 43628 745418 43680 745424
rect 43536 729700 43588 729706
rect 43536 729642 43588 729648
rect 42524 729564 42576 729570
rect 42524 729506 42576 729512
rect 43076 729564 43128 729570
rect 43076 729506 43128 729512
rect 41510 729464 41566 729473
rect 41510 729399 41566 729408
rect 41786 728920 41842 728929
rect 41786 728855 41788 728864
rect 41840 728855 41842 728864
rect 41788 728826 41840 728832
rect 42536 728754 42564 729506
rect 42524 728748 42576 728754
rect 42524 728690 42576 728696
rect 39762 728240 39818 728249
rect 39762 728175 39818 728184
rect 42536 727297 42564 728690
rect 43824 728654 43852 765598
rect 43916 743102 43944 766362
rect 44008 757518 44036 769927
rect 44100 766290 44128 770743
rect 44088 766284 44140 766290
rect 44088 766226 44140 766232
rect 44088 766148 44140 766154
rect 44088 766090 44140 766096
rect 43996 757512 44048 757518
rect 43996 757454 44048 757460
rect 43996 757376 44048 757382
rect 43996 757318 44048 757324
rect 44008 750514 44036 757318
rect 43996 750508 44048 750514
rect 43996 750450 44048 750456
rect 44100 747974 44128 766090
rect 44008 747946 44128 747974
rect 43904 743096 43956 743102
rect 43904 743038 43956 743044
rect 44008 742626 44036 747946
rect 43996 742620 44048 742626
rect 43996 742562 44048 742568
rect 44178 730144 44234 730153
rect 44178 730079 44234 730088
rect 43640 728626 43852 728654
rect 43640 728521 43668 728626
rect 43626 728512 43682 728521
rect 43626 728447 43682 728456
rect 42522 727288 42578 727297
rect 42522 727223 42578 727232
rect 43534 726880 43590 726889
rect 43534 726815 43590 726824
rect 42890 726472 42946 726481
rect 42890 726407 42946 726416
rect 41878 724840 41934 724849
rect 41878 724775 41934 724784
rect 41326 723752 41382 723761
rect 41326 723687 41382 723696
rect 41340 717602 41368 723687
rect 41510 720896 41566 720905
rect 41510 720831 41566 720840
rect 41524 719681 41552 720831
rect 41510 719672 41566 719681
rect 41510 719607 41512 719616
rect 41564 719607 41566 719616
rect 41512 719578 41564 719584
rect 41328 717596 41380 717602
rect 41328 717538 41380 717544
rect 41892 713862 41920 724775
rect 42798 723208 42854 723217
rect 42798 723143 42854 723152
rect 42524 716644 42576 716650
rect 42524 716586 42576 716592
rect 41880 713856 41932 713862
rect 41880 713798 41932 713804
rect 41880 713584 41932 713590
rect 41880 713526 41932 713532
rect 41892 713048 41920 713526
rect 42156 711680 42208 711686
rect 42156 711622 42208 711628
rect 42168 711212 42196 711622
rect 42536 711142 42564 716586
rect 42156 711136 42208 711142
rect 42156 711078 42208 711084
rect 42524 711136 42576 711142
rect 42524 711078 42576 711084
rect 42168 710561 42196 711078
rect 42812 709918 42840 723143
rect 42904 711686 42932 726407
rect 43258 726064 43314 726073
rect 43258 725999 43314 726008
rect 42982 724432 43038 724441
rect 42982 724367 43038 724376
rect 42892 711680 42944 711686
rect 42892 711622 42944 711628
rect 42996 711498 43024 724367
rect 43074 723616 43130 723625
rect 43074 723551 43130 723560
rect 42904 711470 43024 711498
rect 42156 709912 42208 709918
rect 42156 709854 42208 709860
rect 42800 709912 42852 709918
rect 42800 709854 42852 709860
rect 42168 709376 42196 709854
rect 42800 709776 42852 709782
rect 42800 709718 42852 709724
rect 42156 708620 42208 708626
rect 42156 708562 42208 708568
rect 42168 708152 42196 708562
rect 42156 708076 42208 708082
rect 42156 708018 42208 708024
rect 42168 707540 42196 708018
rect 42156 707396 42208 707402
rect 42156 707338 42208 707344
rect 42168 706860 42196 707338
rect 42156 706784 42208 706790
rect 42156 706726 42208 706732
rect 42168 706316 42196 706726
rect 42248 704880 42300 704886
rect 42248 704822 42300 704828
rect 42064 704268 42116 704274
rect 42064 704210 42116 704216
rect 42076 703868 42104 704210
rect 42260 703202 42288 704822
rect 42182 703174 42288 703202
rect 42064 702908 42116 702914
rect 42064 702850 42116 702856
rect 42076 702576 42104 702850
rect 42064 702432 42116 702438
rect 42064 702374 42116 702380
rect 42076 702032 42104 702374
rect 42156 700460 42208 700466
rect 42156 700402 42208 700408
rect 42168 700165 42196 700402
rect 42156 700052 42208 700058
rect 42156 699994 42208 700000
rect 42168 699516 42196 699994
rect 42812 699446 42840 709718
rect 42904 700058 42932 711470
rect 42984 711408 43036 711414
rect 42984 711350 43036 711356
rect 42892 700052 42944 700058
rect 42892 699994 42944 700000
rect 42064 699440 42116 699446
rect 42064 699382 42116 699388
rect 42800 699440 42852 699446
rect 42800 699382 42852 699388
rect 42076 698904 42104 699382
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 41512 688424 41564 688430
rect 41510 688392 41512 688401
rect 41564 688392 41566 688401
rect 41510 688327 41566 688336
rect 41696 688084 41748 688090
rect 41696 688026 41748 688032
rect 41708 687585 41736 688026
rect 41788 687744 41840 687750
rect 41786 687712 41788 687721
rect 41840 687712 41842 687721
rect 41786 687647 41842 687656
rect 41694 687576 41750 687585
rect 41694 687511 41750 687520
rect 42996 684865 43024 711350
rect 43088 704886 43116 723551
rect 43166 721576 43222 721585
rect 43166 721511 43222 721520
rect 43180 708626 43208 721511
rect 43272 709782 43300 725999
rect 43442 725656 43498 725665
rect 43442 725591 43498 725600
rect 43350 725248 43406 725257
rect 43350 725183 43406 725192
rect 43260 709776 43312 709782
rect 43260 709718 43312 709724
rect 43364 709334 43392 725183
rect 43272 709306 43392 709334
rect 43168 708620 43220 708626
rect 43168 708562 43220 708568
rect 43272 706790 43300 709306
rect 43260 706784 43312 706790
rect 43260 706726 43312 706732
rect 43076 704880 43128 704886
rect 43076 704822 43128 704828
rect 43456 702438 43484 725591
rect 43444 702432 43496 702438
rect 43444 702374 43496 702380
rect 43548 700466 43576 726815
rect 43640 711414 43668 728447
rect 43902 722800 43958 722809
rect 43902 722735 43958 722744
rect 43810 721984 43866 721993
rect 43810 721919 43866 721928
rect 43720 717596 43772 717602
rect 43720 717538 43772 717544
rect 43628 711408 43680 711414
rect 43628 711350 43680 711356
rect 43732 702914 43760 717538
rect 43824 707402 43852 721919
rect 43916 708082 43944 722735
rect 43994 722392 44050 722401
rect 43994 722327 44050 722336
rect 43904 708076 43956 708082
rect 43904 708018 43956 708024
rect 43812 707396 43864 707402
rect 43812 707338 43864 707344
rect 44008 704274 44036 722327
rect 43996 704268 44048 704274
rect 43996 704210 44048 704216
rect 43720 702908 43772 702914
rect 43720 702850 43772 702856
rect 43536 700460 43588 700466
rect 43536 700402 43588 700408
rect 44192 686497 44220 730079
rect 44364 728884 44416 728890
rect 44364 728826 44416 728832
rect 44270 727696 44326 727705
rect 44270 727631 44326 727640
rect 44178 686488 44234 686497
rect 44178 686423 44234 686432
rect 43166 685672 43222 685681
rect 43166 685607 43222 685616
rect 42982 684856 43038 684865
rect 42982 684791 43038 684800
rect 42798 684448 42854 684457
rect 42798 684383 42854 684392
rect 41694 681864 41750 681873
rect 41340 681822 41694 681850
rect 41340 673470 41368 681822
rect 41694 681799 41750 681808
rect 42812 681698 42840 684383
rect 43074 682816 43130 682825
rect 43074 682751 43130 682760
rect 42982 682408 43038 682417
rect 42982 682343 43038 682352
rect 42800 681692 42852 681698
rect 42800 681634 42852 681640
rect 41878 681592 41934 681601
rect 41878 681527 41934 681536
rect 41786 678736 41842 678745
rect 41786 678671 41842 678680
rect 41800 678366 41828 678671
rect 41788 678360 41840 678366
rect 41788 678302 41840 678308
rect 41786 677920 41842 677929
rect 41786 677855 41842 677864
rect 41800 676705 41828 677855
rect 41786 676696 41842 676705
rect 41786 676631 41788 676640
rect 41840 676631 41842 676640
rect 41788 676602 41840 676608
rect 41328 673464 41380 673470
rect 41328 673406 41380 673412
rect 41892 670614 41920 681527
rect 41970 678328 42026 678337
rect 41970 678263 42026 678272
rect 41984 670614 42012 678263
rect 41880 670608 41932 670614
rect 41880 670550 41932 670556
rect 41972 670608 42024 670614
rect 41972 670550 42024 670556
rect 42708 670608 42760 670614
rect 42708 670550 42760 670556
rect 41880 670404 41932 670410
rect 41880 670346 41932 670352
rect 41892 669868 41920 670346
rect 42064 668500 42116 668506
rect 42064 668442 42116 668448
rect 42076 668032 42104 668442
rect 42156 667752 42208 667758
rect 42156 667694 42208 667700
rect 42168 667352 42196 667694
rect 42156 666732 42208 666738
rect 42156 666674 42208 666680
rect 42168 666165 42196 666674
rect 42720 665446 42748 670550
rect 42156 665440 42208 665446
rect 42156 665382 42208 665388
rect 42708 665440 42760 665446
rect 42708 665382 42760 665388
rect 42168 664972 42196 665382
rect 42156 664692 42208 664698
rect 42156 664634 42208 664640
rect 42168 664325 42196 664634
rect 42156 664012 42208 664018
rect 42156 663954 42208 663960
rect 42168 663680 42196 663954
rect 42156 663604 42208 663610
rect 42156 663546 42208 663552
rect 42168 663136 42196 663546
rect 42156 661088 42208 661094
rect 42156 661030 42208 661036
rect 42168 660620 42196 661030
rect 42156 660544 42208 660550
rect 42156 660486 42208 660492
rect 42168 660008 42196 660486
rect 42156 659932 42208 659938
rect 42156 659874 42208 659880
rect 42168 659357 42196 659874
rect 42156 659252 42208 659258
rect 42156 659194 42208 659200
rect 42168 658784 42196 659194
rect 42156 657280 42208 657286
rect 42156 657222 42208 657228
rect 42168 656948 42196 657222
rect 42156 656872 42208 656878
rect 42156 656814 42208 656820
rect 42168 656336 42196 656814
rect 42156 656192 42208 656198
rect 42156 656134 42208 656140
rect 42168 655656 42196 656134
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 41512 645176 41564 645182
rect 41510 645144 41512 645153
rect 41564 645144 41566 645153
rect 41510 645079 41566 645088
rect 41512 644836 41564 644842
rect 41512 644778 41564 644784
rect 41524 644337 41552 644778
rect 41788 644564 41840 644570
rect 41786 644532 41788 644541
rect 41840 644532 41842 644541
rect 41786 644467 41842 644476
rect 41510 644328 41566 644337
rect 41510 644263 41566 644272
rect 42812 641073 42840 681634
rect 42892 673464 42944 673470
rect 42892 673406 42944 673412
rect 42904 663610 42932 673406
rect 42892 663604 42944 663610
rect 42892 663546 42944 663552
rect 42996 659258 43024 682343
rect 42984 659252 43036 659258
rect 42984 659194 43036 659200
rect 43088 656198 43116 682751
rect 43076 656192 43128 656198
rect 43076 656134 43128 656140
rect 43180 643113 43208 685607
rect 43350 685264 43406 685273
rect 43350 685199 43406 685208
rect 43258 680776 43314 680785
rect 43258 680711 43314 680720
rect 43272 659938 43300 680711
rect 43260 659932 43312 659938
rect 43260 659874 43312 659880
rect 43166 643104 43222 643113
rect 43166 643039 43222 643048
rect 43364 641889 43392 685199
rect 44284 684049 44312 727631
rect 44376 686089 44404 728826
rect 44362 686080 44418 686089
rect 44362 686015 44418 686024
rect 44270 684040 44326 684049
rect 44270 683975 44326 683984
rect 43626 683632 43682 683641
rect 43626 683567 43682 683576
rect 43442 680368 43498 680377
rect 43442 680303 43498 680312
rect 43456 660550 43484 680303
rect 43534 679552 43590 679561
rect 43534 679487 43590 679496
rect 43548 664698 43576 679487
rect 43536 664692 43588 664698
rect 43536 664634 43588 664640
rect 43444 660544 43496 660550
rect 43444 660486 43496 660492
rect 43640 657286 43668 683567
rect 43902 683224 43958 683233
rect 43902 683159 43958 683168
rect 43810 681184 43866 681193
rect 43810 681119 43866 681128
rect 43718 679960 43774 679969
rect 43718 679895 43774 679904
rect 43732 666738 43760 679895
rect 43824 670682 43852 681119
rect 43812 670676 43864 670682
rect 43812 670618 43864 670624
rect 43812 670472 43864 670478
rect 43812 670414 43864 670420
rect 43720 666732 43772 666738
rect 43720 666674 43772 666680
rect 43824 661094 43852 670414
rect 43916 668506 43944 683159
rect 43994 679144 44050 679153
rect 43994 679079 44050 679088
rect 44008 670682 44036 679079
rect 44088 678360 44140 678366
rect 44088 678302 44140 678308
rect 44100 670682 44128 678302
rect 44180 670744 44232 670750
rect 44180 670686 44232 670692
rect 43996 670676 44048 670682
rect 43996 670618 44048 670624
rect 44088 670676 44140 670682
rect 44088 670618 44140 670624
rect 43996 670472 44048 670478
rect 43996 670414 44048 670420
rect 43904 668500 43956 668506
rect 43904 668442 43956 668448
rect 44008 664018 44036 670414
rect 44192 670290 44220 670686
rect 44100 670262 44220 670290
rect 44100 667758 44128 670262
rect 44180 670200 44232 670206
rect 44180 670142 44232 670148
rect 44088 667752 44140 667758
rect 44088 667694 44140 667700
rect 44192 667570 44220 670142
rect 44100 667542 44220 667570
rect 43996 664012 44048 664018
rect 43996 663954 44048 663960
rect 43812 661088 43864 661094
rect 43812 661030 43864 661036
rect 43628 657280 43680 657286
rect 43628 657222 43680 657228
rect 44100 656878 44128 667542
rect 44088 656872 44140 656878
rect 44088 656814 44140 656820
rect 44086 643512 44142 643521
rect 44142 643470 44220 643498
rect 44086 643447 44142 643456
rect 43350 641880 43406 641889
rect 43350 641815 43406 641824
rect 42798 641064 42854 641073
rect 42798 640999 42854 641008
rect 43350 640384 43406 640393
rect 43350 640319 43406 640328
rect 42798 639432 42854 639441
rect 42798 639367 42854 639376
rect 41786 638412 41842 638421
rect 41786 638347 41842 638356
rect 30286 634944 30342 634953
rect 30286 634879 30342 634888
rect 30300 627910 30328 634879
rect 41510 634536 41566 634545
rect 41510 634471 41566 634480
rect 41524 633321 41552 634471
rect 41510 633312 41566 633321
rect 41510 633247 41512 633256
rect 41564 633247 41566 633256
rect 41512 633218 41564 633224
rect 30288 627904 30340 627910
rect 30288 627846 30340 627852
rect 41800 627434 41828 638347
rect 42524 627904 42576 627910
rect 42524 627846 42576 627852
rect 41788 627428 41840 627434
rect 41788 627370 41840 627376
rect 41788 627088 41840 627094
rect 41788 627030 41840 627036
rect 41800 626620 41828 627030
rect 42156 625320 42208 625326
rect 42156 625262 42208 625268
rect 42168 624784 42196 625262
rect 42156 624708 42208 624714
rect 42156 624650 42208 624656
rect 42168 624172 42196 624650
rect 42156 623484 42208 623490
rect 42156 623426 42208 623432
rect 42168 622948 42196 623426
rect 42536 622198 42564 627846
rect 42064 622192 42116 622198
rect 42064 622134 42116 622140
rect 42524 622192 42576 622198
rect 42524 622134 42576 622140
rect 42076 621792 42104 622134
rect 42156 621512 42208 621518
rect 42156 621454 42208 621460
rect 42168 621112 42196 621454
rect 42064 621036 42116 621042
rect 42064 620978 42116 620984
rect 42076 620500 42104 620978
rect 42064 620220 42116 620226
rect 42064 620162 42116 620168
rect 42076 619956 42104 620162
rect 42248 619064 42300 619070
rect 42248 619006 42300 619012
rect 42156 617908 42208 617914
rect 42156 617850 42208 617856
rect 42168 617440 42196 617850
rect 42064 617364 42116 617370
rect 42064 617306 42116 617312
rect 42076 616828 42104 617306
rect 42260 616162 42288 619006
rect 42182 616134 42288 616162
rect 42248 616072 42300 616078
rect 42248 616014 42300 616020
rect 42260 615618 42288 616014
rect 42182 615590 42288 615618
rect 42156 614236 42208 614242
rect 42156 614178 42208 614184
rect 42168 613768 42196 614178
rect 42156 613692 42208 613698
rect 42156 613634 42208 613640
rect 42168 613121 42196 613634
rect 42812 613018 42840 639367
rect 42982 637800 43038 637809
rect 42982 637735 43038 637744
rect 42890 637664 42946 637673
rect 42890 637599 42946 637608
rect 42904 619070 42932 637599
rect 42892 619064 42944 619070
rect 42892 619006 42944 619012
rect 42996 613698 43024 637735
rect 43074 636576 43130 636585
rect 43074 636511 43130 636520
rect 43088 623490 43116 636511
rect 43258 636168 43314 636177
rect 43258 636103 43314 636112
rect 43166 635352 43222 635361
rect 43166 635287 43222 635296
rect 43076 623484 43128 623490
rect 43076 623426 43128 623432
rect 43180 621042 43208 635287
rect 43272 621518 43300 636103
rect 43260 621512 43312 621518
rect 43260 621454 43312 621460
rect 43168 621036 43220 621042
rect 43168 620978 43220 620984
rect 43364 614242 43392 640319
rect 43718 639840 43774 639849
rect 43718 639775 43774 639784
rect 43534 639024 43590 639033
rect 43534 638959 43590 638968
rect 43442 636984 43498 636993
rect 43442 636919 43498 636928
rect 43456 617370 43484 636919
rect 43444 617364 43496 617370
rect 43444 617306 43496 617312
rect 43548 616078 43576 638959
rect 43628 629332 43680 629338
rect 43628 629274 43680 629280
rect 43640 624714 43668 629274
rect 43732 625326 43760 639775
rect 43902 638616 43958 638625
rect 43902 638551 43958 638560
rect 43810 635760 43866 635769
rect 43810 635695 43866 635704
rect 43720 625320 43772 625326
rect 43720 625262 43772 625268
rect 43628 624708 43680 624714
rect 43628 624650 43680 624656
rect 43824 617914 43852 635695
rect 43916 620226 43944 638551
rect 43904 620220 43956 620226
rect 43904 620162 43956 620168
rect 43812 617908 43864 617914
rect 43812 617850 43864 617856
rect 43536 616072 43588 616078
rect 43536 616014 43588 616020
rect 43352 614236 43404 614242
rect 43352 614178 43404 614184
rect 42984 613692 43036 613698
rect 42984 613634 43036 613640
rect 42156 613012 42208 613018
rect 42156 612954 42208 612960
rect 42800 613012 42852 613018
rect 42800 612954 42852 612960
rect 42168 612476 42196 612954
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 41512 601928 41564 601934
rect 41510 601896 41512 601905
rect 41564 601896 41566 601905
rect 41510 601831 41566 601840
rect 42430 600536 42486 600545
rect 42430 600471 42486 600480
rect 42444 598942 42472 600471
rect 44192 600137 44220 643470
rect 44822 642288 44878 642297
rect 44822 642223 44878 642232
rect 44362 642016 44418 642025
rect 44362 641951 44418 641960
rect 44178 600128 44234 600137
rect 44178 600063 44234 600072
rect 43442 599312 43498 599321
rect 43442 599247 43498 599256
rect 42432 598936 42484 598942
rect 42432 598878 42484 598884
rect 41878 595232 41934 595241
rect 41878 595167 41934 595176
rect 41142 594144 41198 594153
rect 41142 594079 41198 594088
rect 41156 585206 41184 594079
rect 41510 591288 41566 591297
rect 41510 591223 41566 591232
rect 41524 590073 41552 591223
rect 41510 590064 41566 590073
rect 41510 589999 41512 590008
rect 41564 589999 41566 590008
rect 41512 589970 41564 589976
rect 41144 585200 41196 585206
rect 41144 585142 41196 585148
rect 41892 584254 41920 595167
rect 41880 584248 41932 584254
rect 41880 584190 41932 584196
rect 41880 583976 41932 583982
rect 41880 583918 41932 583924
rect 41892 583440 41920 583918
rect 42444 583778 42472 598878
rect 43258 597272 43314 597281
rect 43258 597207 43314 597216
rect 42890 596864 42946 596873
rect 42890 596799 42946 596808
rect 42798 593600 42854 593609
rect 42798 593535 42854 593544
rect 42812 586634 42840 593535
rect 42800 586628 42852 586634
rect 42800 586570 42852 586576
rect 42904 583930 42932 596799
rect 43074 596456 43130 596465
rect 43074 596391 43130 596400
rect 42982 594824 43038 594833
rect 42982 594759 43038 594768
rect 42720 583902 42932 583930
rect 42432 583772 42484 583778
rect 42432 583714 42484 583720
rect 42720 582146 42748 583902
rect 42800 583772 42852 583778
rect 42800 583714 42852 583720
rect 42892 583772 42944 583778
rect 42892 583714 42944 583720
rect 42156 582140 42208 582146
rect 42156 582082 42208 582088
rect 42708 582140 42760 582146
rect 42708 582082 42760 582088
rect 42168 581604 42196 582082
rect 42156 581324 42208 581330
rect 42156 581266 42208 581272
rect 42168 580961 42196 581266
rect 42156 580304 42208 580310
rect 42156 580246 42208 580252
rect 42168 579768 42196 580246
rect 42156 579012 42208 579018
rect 42156 578954 42208 578960
rect 42168 578544 42196 578954
rect 42156 578468 42208 578474
rect 42156 578410 42208 578416
rect 42168 577932 42196 578410
rect 42156 577856 42208 577862
rect 42156 577798 42208 577804
rect 42168 577281 42196 577798
rect 42156 576972 42208 576978
rect 42156 576914 42208 576920
rect 42168 576708 42196 576914
rect 42156 574728 42208 574734
rect 42156 574670 42208 574676
rect 42168 574260 42196 574670
rect 42156 573844 42208 573850
rect 42156 573786 42208 573792
rect 42168 573580 42196 573786
rect 42156 573504 42208 573510
rect 42156 573446 42208 573452
rect 42168 572968 42196 573446
rect 42064 572688 42116 572694
rect 42064 572630 42116 572636
rect 42076 572424 42104 572630
rect 42064 570920 42116 570926
rect 42064 570862 42116 570868
rect 42076 570588 42104 570862
rect 42156 570308 42208 570314
rect 42156 570250 42208 570256
rect 42168 569908 42196 570250
rect 42064 569628 42116 569634
rect 42064 569570 42116 569576
rect 42076 569296 42104 569570
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 41512 558816 41564 558822
rect 41510 558784 41512 558793
rect 41564 558784 41566 558793
rect 41510 558719 41566 558728
rect 41420 558544 41472 558550
rect 41420 558486 41472 558492
rect 41432 557977 41460 558486
rect 41512 558476 41564 558482
rect 41512 558418 41564 558424
rect 41524 558385 41552 558418
rect 41510 558376 41566 558385
rect 41510 558311 41566 558320
rect 41418 557968 41474 557977
rect 41418 557903 41474 557912
rect 42812 556889 42840 583714
rect 42904 569634 42932 583714
rect 42996 570314 43024 594759
rect 43088 583778 43116 596391
rect 43166 594008 43222 594017
rect 43166 593943 43222 593952
rect 43076 583772 43128 583778
rect 43076 583714 43128 583720
rect 43076 583636 43128 583642
rect 43076 583578 43128 583584
rect 43088 570926 43116 583578
rect 43180 573850 43208 593943
rect 43272 583642 43300 597207
rect 43350 595640 43406 595649
rect 43350 595575 43406 595584
rect 43364 586770 43392 595575
rect 43352 586764 43404 586770
rect 43352 586706 43404 586712
rect 43352 586628 43404 586634
rect 43352 586570 43404 586576
rect 43260 583636 43312 583642
rect 43260 583578 43312 583584
rect 43260 583500 43312 583506
rect 43260 583442 43312 583448
rect 43168 573844 43220 573850
rect 43168 573786 43220 573792
rect 43076 570920 43128 570926
rect 43076 570862 43128 570868
rect 42984 570308 43036 570314
rect 42984 570250 43036 570256
rect 42892 569628 42944 569634
rect 42892 569570 42944 569576
rect 42798 556880 42854 556889
rect 42798 556815 42854 556824
rect 43272 554441 43300 583442
rect 43364 580310 43392 586570
rect 43352 580304 43404 580310
rect 43352 580246 43404 580252
rect 43456 556481 43484 599247
rect 44376 598505 44404 641951
rect 44638 641200 44694 641209
rect 44638 641135 44694 641144
rect 44362 598496 44418 598505
rect 44362 598431 44418 598440
rect 43994 598088 44050 598097
rect 43994 598023 44050 598032
rect 43810 596048 43866 596057
rect 43810 595983 43866 595992
rect 43718 593192 43774 593201
rect 43718 593127 43774 593136
rect 43626 592376 43682 592385
rect 43626 592311 43682 592320
rect 43534 591968 43590 591977
rect 43534 591903 43590 591912
rect 43548 579018 43576 591903
rect 43536 579012 43588 579018
rect 43536 578954 43588 578960
rect 43640 577862 43668 592311
rect 43732 578474 43760 593127
rect 43720 578468 43772 578474
rect 43720 578410 43772 578416
rect 43628 577856 43680 577862
rect 43628 577798 43680 577804
rect 43628 577720 43680 577726
rect 43628 577662 43680 577668
rect 43640 573510 43668 577662
rect 43628 573504 43680 573510
rect 43628 573446 43680 573452
rect 43824 572694 43852 595983
rect 43902 592784 43958 592793
rect 43902 592719 43958 592728
rect 43916 574734 43944 592719
rect 44008 583506 44036 598023
rect 44652 597689 44680 641135
rect 44836 599729 44864 642223
rect 44822 599720 44878 599729
rect 44822 599655 44878 599664
rect 44638 597680 44694 597689
rect 44638 597615 44694 597624
rect 44088 586764 44140 586770
rect 44088 586706 44140 586712
rect 44100 583506 44128 586706
rect 44180 585200 44232 585206
rect 44180 585142 44232 585148
rect 44272 585200 44324 585206
rect 44272 585142 44324 585148
rect 43996 583500 44048 583506
rect 43996 583442 44048 583448
rect 44088 583500 44140 583506
rect 44088 583442 44140 583448
rect 44192 583386 44220 585142
rect 44008 583358 44220 583386
rect 44008 577726 44036 583358
rect 44088 583160 44140 583166
rect 44088 583102 44140 583108
rect 43996 577720 44048 577726
rect 43996 577662 44048 577668
rect 44100 576978 44128 583102
rect 44284 581330 44312 585142
rect 44272 581324 44324 581330
rect 44272 581266 44324 581272
rect 44088 576972 44140 576978
rect 44088 576914 44140 576920
rect 43904 574728 43956 574734
rect 43904 574670 43956 574676
rect 43812 572688 43864 572694
rect 43812 572630 43864 572636
rect 43442 556472 43498 556481
rect 43442 556407 43498 556416
rect 43258 554432 43314 554441
rect 43258 554367 43314 554376
rect 43810 554024 43866 554033
rect 43810 553959 43866 553968
rect 42706 553616 42762 553625
rect 42706 553551 42762 553560
rect 41786 551984 41842 551993
rect 41786 551919 41842 551928
rect 41510 548992 41566 549001
rect 41510 548927 41566 548936
rect 41524 548690 41552 548927
rect 41512 548684 41564 548690
rect 41512 548626 41564 548632
rect 41510 548584 41566 548593
rect 41510 548519 41566 548528
rect 41524 546786 41552 548519
rect 41602 548176 41658 548185
rect 41602 548111 41658 548120
rect 41616 546961 41644 548111
rect 41602 546952 41658 546961
rect 41602 546887 41604 546896
rect 41656 546887 41658 546896
rect 41604 546858 41656 546864
rect 41512 546780 41564 546786
rect 41512 546722 41564 546728
rect 41800 541074 41828 551919
rect 41788 541068 41840 541074
rect 41788 541010 41840 541016
rect 41788 540796 41840 540802
rect 41788 540738 41840 540744
rect 41800 540260 41828 540738
rect 42720 538966 42748 553551
rect 43166 553208 43222 553217
rect 43166 553143 43222 553152
rect 43074 551168 43130 551177
rect 43074 551103 43130 551112
rect 42982 550352 43038 550361
rect 42982 550287 43038 550296
rect 42800 546780 42852 546786
rect 42800 546722 42852 546728
rect 42064 538960 42116 538966
rect 42064 538902 42116 538908
rect 42708 538960 42760 538966
rect 42708 538902 42760 538908
rect 42076 538424 42104 538902
rect 42156 538144 42208 538150
rect 42156 538086 42208 538092
rect 42168 537744 42196 538086
rect 42064 537124 42116 537130
rect 42064 537066 42116 537072
rect 42076 536588 42104 537066
rect 42812 535838 42840 546722
rect 42890 540968 42946 540977
rect 42890 540903 42946 540912
rect 42156 535832 42208 535838
rect 42156 535774 42208 535780
rect 42800 535832 42852 535838
rect 42800 535774 42852 535780
rect 42168 535364 42196 535774
rect 42064 535084 42116 535090
rect 42064 535026 42116 535032
rect 42076 534752 42104 535026
rect 42156 534472 42208 534478
rect 42156 534414 42208 534420
rect 42168 534072 42196 534414
rect 42156 533996 42208 534002
rect 42156 533938 42208 533944
rect 42168 533528 42196 533938
rect 42156 531480 42208 531486
rect 42156 531422 42208 531428
rect 42168 531045 42196 531422
rect 42156 530732 42208 530738
rect 42156 530674 42208 530680
rect 42168 530400 42196 530674
rect 42156 530324 42208 530330
rect 42156 530266 42208 530272
rect 42168 529757 42196 530266
rect 42156 529508 42208 529514
rect 42156 529450 42208 529456
rect 42168 529205 42196 529450
rect 42076 527202 42104 527340
rect 42156 527264 42208 527270
rect 42156 527206 42208 527212
rect 42064 527196 42116 527202
rect 42064 527138 42116 527144
rect 42168 526728 42196 527206
rect 42156 526652 42208 526658
rect 42156 526594 42208 526600
rect 42168 526077 42196 526594
rect 42904 450809 42932 540903
rect 42996 537130 43024 550287
rect 42984 537124 43036 537130
rect 42984 537066 43036 537072
rect 42984 536988 43036 536994
rect 42984 536930 43036 536936
rect 42996 526658 43024 536930
rect 43088 530330 43116 551103
rect 43180 536994 43208 553143
rect 43350 552800 43406 552809
rect 43350 552735 43406 552744
rect 43258 549944 43314 549953
rect 43258 549879 43314 549888
rect 43168 536988 43220 536994
rect 43168 536930 43220 536936
rect 43168 536852 43220 536858
rect 43168 536794 43220 536800
rect 43076 530324 43128 530330
rect 43076 530266 43128 530272
rect 43180 529514 43208 536794
rect 43272 535090 43300 549879
rect 43364 536858 43392 552735
rect 43626 552392 43682 552401
rect 43626 552327 43682 552336
rect 43442 551576 43498 551585
rect 43442 551511 43498 551520
rect 43352 536852 43404 536858
rect 43352 536794 43404 536800
rect 43352 536716 43404 536722
rect 43352 536658 43404 536664
rect 43260 535084 43312 535090
rect 43260 535026 43312 535032
rect 43364 534002 43392 536658
rect 43352 533996 43404 534002
rect 43352 533938 43404 533944
rect 43168 529508 43220 529514
rect 43168 529450 43220 529456
rect 43456 527270 43484 551511
rect 43536 548684 43588 548690
rect 43536 548626 43588 548632
rect 43548 534478 43576 548626
rect 43640 536722 43668 552327
rect 43720 541748 43772 541754
rect 43720 541690 43772 541696
rect 43732 538150 43760 541690
rect 43720 538144 43772 538150
rect 43720 538086 43772 538092
rect 43628 536716 43680 536722
rect 43628 536658 43680 536664
rect 43536 534472 43588 534478
rect 43536 534414 43588 534420
rect 43444 527264 43496 527270
rect 43444 527206 43496 527212
rect 43824 527202 43852 553959
rect 43994 550760 44050 550769
rect 43994 550695 44050 550704
rect 43902 549536 43958 549545
rect 43902 549471 43958 549480
rect 43916 531486 43944 549471
rect 43904 531480 43956 531486
rect 43904 531422 43956 531428
rect 44008 530738 44036 550695
rect 44086 540832 44142 540841
rect 44086 540767 44142 540776
rect 43996 530732 44048 530738
rect 43996 530674 44048 530680
rect 43812 527196 43864 527202
rect 43812 527138 43864 527144
rect 42984 526652 43036 526658
rect 42984 526594 43036 526600
rect 42890 450800 42946 450809
rect 42890 450735 42946 450744
rect 8588 431596 8616 431732
rect 9048 431596 9076 431732
rect 9508 431596 9536 431732
rect 9968 431596 9996 431732
rect 10428 431596 10456 431732
rect 10888 431596 10916 431732
rect 11348 431596 11376 431732
rect 11808 431596 11836 431732
rect 12268 431596 12296 431732
rect 12728 431596 12756 431732
rect 13188 431596 13216 431732
rect 13648 431596 13676 431732
rect 14108 431596 14136 431732
rect 41786 430944 41842 430953
rect 41786 430879 41842 430888
rect 41800 430846 41828 430879
rect 41788 430840 41840 430846
rect 41788 430782 41840 430788
rect 43074 430672 43130 430681
rect 43074 430607 43130 430616
rect 43088 429321 43116 430607
rect 43626 429720 43682 429729
rect 43626 429655 43682 429664
rect 43074 429312 43130 429321
rect 43074 429247 43130 429256
rect 41788 427848 41840 427854
rect 41788 427790 41840 427796
rect 41800 426873 41828 427790
rect 41786 426864 41842 426873
rect 41786 426799 41842 426808
rect 42890 426456 42946 426465
rect 42890 426391 42946 426400
rect 42798 426048 42854 426057
rect 42798 425983 42854 425992
rect 42338 424416 42394 424425
rect 42338 424351 42394 424360
rect 41878 421560 41934 421569
rect 41878 421495 41934 421504
rect 41786 420744 41842 420753
rect 41786 420679 41842 420688
rect 41800 419529 41828 420679
rect 41786 419520 41842 419529
rect 41786 419455 41788 419464
rect 41840 419455 41842 419464
rect 41788 419426 41840 419432
rect 41892 416362 41920 421495
rect 41880 416356 41932 416362
rect 41880 416298 41932 416304
rect 42352 413166 42380 424351
rect 42522 421152 42578 421161
rect 42522 421087 42578 421096
rect 42156 413160 42208 413166
rect 42156 413102 42208 413108
rect 42340 413160 42392 413166
rect 42340 413102 42392 413108
rect 42168 412624 42196 413102
rect 42156 411324 42208 411330
rect 42156 411266 42208 411272
rect 42168 410788 42196 411266
rect 42156 410712 42208 410718
rect 42156 410654 42208 410660
rect 42168 410176 42196 410654
rect 42156 409488 42208 409494
rect 42156 409430 42208 409436
rect 42168 408952 42196 409430
rect 42536 408202 42564 421087
rect 42812 411398 42840 425983
rect 42800 411392 42852 411398
rect 42800 411334 42852 411340
rect 42798 411268 42854 411277
rect 42798 411203 42854 411212
rect 42064 408196 42116 408202
rect 42064 408138 42116 408144
rect 42524 408196 42576 408202
rect 42524 408138 42576 408144
rect 42076 407796 42104 408138
rect 42156 407516 42208 407522
rect 42156 407458 42208 407464
rect 42168 407116 42196 407458
rect 42064 407040 42116 407046
rect 42064 406982 42116 406988
rect 42076 406504 42104 406982
rect 42156 406224 42208 406230
rect 42156 406166 42208 406172
rect 42168 405929 42196 406166
rect 42156 403912 42208 403918
rect 42156 403854 42208 403860
rect 42168 403444 42196 403854
rect 42156 403368 42208 403374
rect 42156 403310 42208 403316
rect 42168 402801 42196 403310
rect 42156 402552 42208 402558
rect 42156 402494 42208 402500
rect 42168 402152 42196 402494
rect 42156 402076 42208 402082
rect 42156 402018 42208 402024
rect 42168 401608 42196 402018
rect 42156 400036 42208 400042
rect 42156 399978 42208 399984
rect 42168 399772 42196 399978
rect 42156 399492 42208 399498
rect 42156 399434 42208 399440
rect 42168 399121 42196 399434
rect 42156 398812 42208 398818
rect 42156 398754 42208 398760
rect 42168 398480 42196 398754
rect 41142 389056 41198 389065
rect 41142 388991 41198 389000
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41156 386753 41184 388991
rect 41512 388000 41564 388006
rect 41510 387968 41512 387977
rect 41564 387968 41566 387977
rect 41510 387903 41566 387912
rect 41512 387660 41564 387666
rect 41512 387602 41564 387608
rect 41524 387569 41552 387602
rect 41510 387560 41566 387569
rect 41510 387495 41566 387504
rect 41512 387184 41564 387190
rect 41510 387152 41512 387161
rect 41564 387152 41566 387161
rect 41510 387087 41566 387096
rect 41142 386744 41198 386753
rect 41142 386679 41198 386688
rect 41156 384713 41184 386679
rect 42812 386442 42840 411203
rect 42904 400042 42932 426391
rect 43258 425640 43314 425649
rect 43258 425575 43314 425584
rect 42982 422784 43038 422793
rect 42982 422719 43038 422728
rect 42996 409494 43024 422719
rect 43166 422376 43222 422385
rect 43166 422311 43222 422320
rect 43076 416356 43128 416362
rect 43076 416298 43128 416304
rect 42984 409488 43036 409494
rect 42984 409430 43036 409436
rect 43088 407046 43116 416298
rect 43180 407522 43208 422311
rect 43168 407516 43220 407522
rect 43168 407458 43220 407464
rect 43076 407040 43128 407046
rect 43076 406982 43128 406988
rect 42892 400036 42944 400042
rect 42892 399978 42944 399984
rect 43272 398818 43300 425575
rect 43350 425232 43406 425241
rect 43350 425167 43406 425176
rect 43364 402082 43392 425167
rect 43442 424824 43498 424833
rect 43442 424759 43498 424768
rect 43456 406230 43484 424759
rect 43534 423192 43590 423201
rect 43534 423127 43590 423136
rect 43444 406224 43496 406230
rect 43444 406166 43496 406172
rect 43548 403374 43576 423127
rect 43640 411505 43668 429655
rect 43810 428496 43866 428505
rect 43810 428431 43866 428440
rect 43718 423600 43774 423609
rect 43718 423535 43774 423544
rect 43626 411496 43682 411505
rect 43626 411431 43682 411440
rect 43536 403368 43588 403374
rect 43536 403310 43588 403316
rect 43732 402558 43760 423535
rect 43720 402552 43772 402558
rect 43720 402494 43772 402500
rect 43824 402490 43852 428431
rect 44100 427854 44128 540767
rect 44088 427848 44140 427854
rect 44088 427790 44140 427796
rect 43902 424008 43958 424017
rect 43902 423943 43958 423952
rect 43812 402484 43864 402490
rect 43812 402426 43864 402432
rect 43916 402370 43944 423943
rect 43994 421968 44050 421977
rect 43994 421903 44050 421912
rect 44008 403918 44036 421903
rect 43996 403912 44048 403918
rect 43996 403854 44048 403860
rect 43732 402342 43944 402370
rect 43352 402076 43404 402082
rect 43352 402018 43404 402024
rect 43732 399498 43760 402342
rect 43812 402280 43864 402286
rect 43812 402222 43864 402228
rect 43720 399492 43772 399498
rect 43720 399434 43772 399440
rect 43260 398812 43312 398818
rect 43260 398754 43312 398760
rect 42800 386436 42852 386442
rect 42800 386378 42852 386384
rect 42812 386073 42840 386378
rect 42798 386064 42854 386073
rect 42798 385999 42854 386008
rect 43824 385665 43852 402222
rect 43810 385656 43866 385665
rect 43810 385591 43866 385600
rect 43534 385248 43590 385257
rect 43534 385183 43590 385192
rect 41142 384704 41198 384713
rect 41142 384639 41198 384648
rect 43350 383208 43406 383217
rect 43350 383143 43406 383152
rect 42798 382800 42854 382809
rect 42798 382735 42854 382744
rect 42338 381168 42394 381177
rect 42338 381103 42394 381112
rect 41510 377768 41566 377777
rect 41510 377703 41566 377712
rect 41524 371482 41552 377703
rect 41602 377360 41658 377369
rect 41602 377295 41658 377304
rect 41616 376145 41644 377295
rect 41602 376136 41658 376145
rect 41602 376071 41604 376080
rect 41656 376071 41658 376080
rect 41604 376042 41656 376048
rect 41512 371476 41564 371482
rect 41512 371418 41564 371424
rect 42352 369986 42380 381103
rect 42708 371476 42760 371482
rect 42708 371418 42760 371424
rect 42156 369980 42208 369986
rect 42156 369922 42208 369928
rect 42340 369980 42392 369986
rect 42340 369922 42392 369928
rect 42168 369444 42196 369922
rect 42156 368144 42208 368150
rect 42156 368086 42208 368092
rect 42168 367608 42196 368086
rect 42168 366858 42196 366961
rect 42156 366852 42208 366858
rect 42156 366794 42208 366800
rect 42156 366308 42208 366314
rect 42156 366250 42208 366256
rect 42168 365772 42196 366250
rect 42720 365022 42748 371418
rect 42812 368150 42840 382735
rect 42982 381984 43038 381993
rect 42982 381919 43038 381928
rect 42890 379536 42946 379545
rect 42890 379471 42946 379480
rect 42800 368144 42852 368150
rect 42800 368086 42852 368092
rect 42904 366314 42932 379471
rect 42892 366308 42944 366314
rect 42892 366250 42944 366256
rect 42892 366172 42944 366178
rect 42892 366114 42944 366120
rect 42156 365016 42208 365022
rect 42156 364958 42208 364964
rect 42708 365016 42760 365022
rect 42708 364958 42760 364964
rect 42168 364548 42196 364958
rect 42156 364472 42208 364478
rect 42156 364414 42208 364420
rect 42168 363936 42196 364414
rect 42156 363860 42208 363866
rect 42156 363802 42208 363808
rect 42168 363256 42196 363802
rect 42156 363180 42208 363186
rect 42156 363122 42208 363128
rect 42168 362712 42196 363122
rect 42064 360732 42116 360738
rect 42064 360674 42116 360680
rect 42076 360264 42104 360674
rect 42156 359984 42208 359990
rect 42156 359926 42208 359932
rect 42168 359584 42196 359926
rect 42156 359508 42208 359514
rect 42156 359450 42208 359456
rect 42168 358972 42196 359450
rect 42064 358692 42116 358698
rect 42064 358634 42116 358640
rect 42076 358428 42104 358634
rect 42064 356992 42116 356998
rect 42064 356934 42116 356940
rect 42076 356592 42104 356934
rect 42904 356454 42932 366114
rect 42996 358698 43024 381919
rect 43166 379128 43222 379137
rect 43166 379063 43222 379072
rect 43074 378312 43130 378321
rect 43074 378247 43130 378256
rect 43088 363866 43116 378247
rect 43180 364478 43208 379063
rect 43258 378720 43314 378729
rect 43258 378655 43314 378664
rect 43168 364472 43220 364478
rect 43168 364414 43220 364420
rect 43076 363860 43128 363866
rect 43076 363802 43128 363808
rect 43076 363724 43128 363730
rect 43076 363666 43128 363672
rect 43088 359514 43116 363666
rect 43272 360738 43300 378655
rect 43260 360732 43312 360738
rect 43260 360674 43312 360680
rect 43076 359508 43128 359514
rect 43076 359450 43128 359456
rect 42984 358692 43036 358698
rect 42984 358634 43036 358640
rect 43364 356998 43392 383143
rect 43442 380760 43498 380769
rect 43442 380695 43498 380704
rect 43456 366178 43484 380695
rect 43444 366172 43496 366178
rect 43444 366114 43496 366120
rect 43352 356992 43404 356998
rect 43352 356934 43404 356940
rect 42156 356448 42208 356454
rect 42156 356390 42208 356396
rect 42892 356448 42944 356454
rect 42892 356390 42944 356396
rect 42168 355912 42196 356390
rect 41786 355736 41842 355745
rect 41786 355671 41842 355680
rect 41800 355300 41828 355671
rect 33046 351928 33102 351937
rect 33046 351863 33102 351872
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 33060 343097 33088 351863
rect 43548 344758 43576 385183
rect 43902 381576 43958 381585
rect 43902 381511 43958 381520
rect 43626 380352 43682 380361
rect 43626 380287 43682 380296
rect 43640 363730 43668 380287
rect 43718 379944 43774 379953
rect 43718 379879 43774 379888
rect 43628 363724 43680 363730
rect 43628 363666 43680 363672
rect 43732 361574 43760 379879
rect 43916 363186 43944 381511
rect 43904 363180 43956 363186
rect 43904 363122 43956 363128
rect 43640 361546 43760 361574
rect 43640 359990 43668 361546
rect 43628 359984 43680 359990
rect 43628 359926 43680 359932
rect 44180 345024 44232 345030
rect 44180 344966 44232 344972
rect 41512 344752 41564 344758
rect 41512 344694 41564 344700
rect 43536 344752 43588 344758
rect 43536 344694 43588 344700
rect 33046 343088 33102 343097
rect 33046 343023 33102 343032
rect 41524 342689 41552 344694
rect 41786 344584 41842 344593
rect 41786 344519 41842 344528
rect 41800 344486 41828 344519
rect 41788 344480 41840 344486
rect 41788 344422 41840 344428
rect 41604 344344 41656 344350
rect 41602 344312 41604 344321
rect 41656 344312 41658 344321
rect 41602 344247 41658 344256
rect 41604 343936 41656 343942
rect 41602 343904 41604 343913
rect 41656 343904 41658 343913
rect 41602 343839 41658 343848
rect 44192 343398 44220 344966
rect 41788 343392 41840 343398
rect 41786 343360 41788 343369
rect 44180 343392 44232 343398
rect 41840 343360 41842 343369
rect 44180 343334 44232 343340
rect 41786 343295 41842 343304
rect 41510 342680 41566 342689
rect 41510 342615 41566 342624
rect 43258 342136 43314 342145
rect 43258 342071 43314 342080
rect 32678 339824 32734 339833
rect 32678 339759 32734 339768
rect 32692 329866 32720 339759
rect 32770 338192 32826 338201
rect 32770 338127 32826 338136
rect 32680 329860 32732 329866
rect 32680 329802 32732 329808
rect 32784 329769 32812 338127
rect 33046 337784 33102 337793
rect 33046 337719 33102 337728
rect 32862 336152 32918 336161
rect 32862 336087 32918 336096
rect 32876 330002 32904 336087
rect 32954 335744 33010 335753
rect 32954 335679 33010 335688
rect 32864 329996 32916 330002
rect 32864 329938 32916 329944
rect 32968 329934 32996 335679
rect 33060 330138 33088 337719
rect 43074 335608 43130 335617
rect 43074 335543 43130 335552
rect 42982 335200 43038 335209
rect 42982 335135 43038 335144
rect 41510 334112 41566 334121
rect 41510 334047 41566 334056
rect 41524 332897 41552 334047
rect 41510 332888 41566 332897
rect 41510 332823 41512 332832
rect 41564 332823 41566 332832
rect 41512 332794 41564 332800
rect 33048 330132 33100 330138
rect 33048 330074 33100 330080
rect 41880 330132 41932 330138
rect 41880 330074 41932 330080
rect 32956 329928 33008 329934
rect 32956 329870 33008 329876
rect 32770 329760 32826 329769
rect 32770 329695 32826 329704
rect 41892 327010 41920 330074
rect 42892 329996 42944 330002
rect 42892 329938 42944 329944
rect 42800 329860 42852 329866
rect 42800 329802 42852 329808
rect 41880 327004 41932 327010
rect 41880 326946 41932 326952
rect 41880 326800 41932 326806
rect 41880 326742 41932 326748
rect 41892 326264 41920 326742
rect 42812 324970 42840 329802
rect 42064 324964 42116 324970
rect 42064 324906 42116 324912
rect 42800 324964 42852 324970
rect 42800 324906 42852 324912
rect 42076 324428 42104 324906
rect 42800 324828 42852 324834
rect 42800 324770 42852 324776
rect 42168 323338 42196 323748
rect 42156 323332 42208 323338
rect 42156 323274 42208 323280
rect 42616 323332 42668 323338
rect 42616 323274 42668 323280
rect 42064 323128 42116 323134
rect 42064 323070 42116 323076
rect 42076 322592 42104 323070
rect 42156 321836 42208 321842
rect 42156 321778 42208 321784
rect 42168 321368 42196 321778
rect 42156 321088 42208 321094
rect 42156 321030 42208 321036
rect 42168 320725 42196 321030
rect 42156 320612 42208 320618
rect 42156 320554 42208 320560
rect 42168 320076 42196 320554
rect 42628 320142 42656 323274
rect 42616 320136 42668 320142
rect 42616 320078 42668 320084
rect 41786 319968 41842 319977
rect 41786 319903 41842 319912
rect 41800 319532 41828 319903
rect 42812 317490 42840 324770
rect 42904 323134 42932 329938
rect 42892 323128 42944 323134
rect 42892 323070 42944 323076
rect 42996 320618 43024 335135
rect 43088 324834 43116 335543
rect 43166 334792 43222 334801
rect 43166 334727 43222 334736
rect 43180 324834 43208 334727
rect 43076 324828 43128 324834
rect 43076 324770 43128 324776
rect 43168 324828 43220 324834
rect 43168 324770 43220 324776
rect 43272 324714 43300 342071
rect 43352 329928 43404 329934
rect 43352 329870 43404 329876
rect 43088 324686 43300 324714
rect 42984 320612 43036 320618
rect 42984 320554 43036 320560
rect 42156 317484 42208 317490
rect 42156 317426 42208 317432
rect 42800 317484 42852 317490
rect 42800 317426 42852 317432
rect 42168 317045 42196 317426
rect 42154 316976 42210 316985
rect 42154 316911 42210 316920
rect 42168 316404 42196 316911
rect 42154 316296 42210 316305
rect 42154 316231 42210 316240
rect 42168 315757 42196 316231
rect 41970 315616 42026 315625
rect 41970 315551 42026 315560
rect 41984 315180 42012 315551
rect 41878 313848 41934 313857
rect 41878 313783 41934 313792
rect 41892 313344 41920 313783
rect 41786 313032 41842 313041
rect 41786 312967 41842 312976
rect 41800 312732 41828 312967
rect 42154 312352 42210 312361
rect 42154 312287 42210 312296
rect 42168 312052 42196 312287
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41512 301640 41564 301646
rect 41510 301608 41512 301617
rect 41564 301608 41566 301617
rect 41510 301543 41566 301552
rect 41788 300960 41840 300966
rect 41786 300928 41788 300937
rect 41840 300928 41842 300937
rect 41786 300863 41842 300872
rect 43088 299305 43116 324686
rect 43168 324624 43220 324630
rect 43168 324566 43220 324572
rect 43180 321842 43208 324566
rect 43168 321836 43220 321842
rect 43168 321778 43220 321784
rect 43364 321094 43392 329870
rect 43352 321088 43404 321094
rect 43352 321030 43404 321036
rect 44192 299713 44220 343334
rect 44270 341728 44326 341737
rect 44270 341663 44326 341672
rect 44284 339969 44312 341663
rect 44362 340912 44418 340921
rect 44362 340847 44418 340856
rect 44270 339960 44326 339969
rect 44270 339895 44326 339904
rect 44178 299704 44234 299713
rect 44178 299639 44234 299648
rect 43074 299296 43130 299305
rect 43074 299231 43130 299240
rect 43442 298888 43498 298897
rect 43442 298823 43498 298832
rect 32586 296848 32642 296857
rect 32586 296783 32642 296792
rect 32600 285705 32628 296783
rect 32678 296440 32734 296449
rect 32678 296375 32734 296384
rect 32692 285802 32720 296375
rect 32954 296032 33010 296041
rect 32954 295967 33010 295976
rect 32862 295216 32918 295225
rect 32862 295151 32918 295160
rect 32770 292360 32826 292369
rect 32770 292295 32826 292304
rect 32680 285796 32732 285802
rect 32680 285738 32732 285744
rect 32586 285696 32642 285705
rect 32784 285666 32812 292295
rect 32876 285734 32904 295151
rect 32968 285841 32996 295967
rect 41878 294808 41934 294817
rect 41878 294743 41934 294752
rect 33046 294400 33102 294409
rect 33046 294335 33102 294344
rect 33060 285977 33088 294335
rect 41786 293992 41842 294001
rect 41786 293927 41842 293936
rect 41800 292058 41828 293927
rect 41788 292052 41840 292058
rect 41788 291994 41840 292000
rect 41786 291952 41842 291961
rect 41786 291887 41842 291896
rect 41800 291650 41828 291887
rect 41788 291644 41840 291650
rect 41788 291586 41840 291592
rect 41786 291544 41842 291553
rect 41786 291479 41842 291488
rect 41800 289882 41828 291479
rect 41892 291174 41920 294743
rect 42430 293584 42486 293593
rect 42430 293519 42486 293528
rect 41880 291168 41932 291174
rect 41880 291110 41932 291116
rect 41788 289876 41840 289882
rect 41788 289818 41840 289824
rect 33046 285968 33102 285977
rect 33046 285903 33102 285912
rect 32954 285832 33010 285841
rect 32954 285767 33010 285776
rect 32864 285728 32916 285734
rect 32864 285670 32916 285676
rect 32586 285631 32642 285640
rect 32772 285660 32824 285666
rect 32772 285602 32824 285608
rect 42156 283620 42208 283626
rect 42156 283562 42208 283568
rect 42168 283045 42196 283562
rect 42444 283354 42472 293519
rect 43074 293176 43130 293185
rect 43074 293111 43130 293120
rect 42708 291168 42760 291174
rect 42708 291110 42760 291116
rect 42720 283626 42748 291110
rect 42800 285796 42852 285802
rect 42800 285738 42852 285744
rect 42708 283620 42760 283626
rect 42708 283562 42760 283568
rect 42432 283348 42484 283354
rect 42432 283290 42484 283296
rect 42708 283348 42760 283354
rect 42708 283290 42760 283296
rect 42156 281784 42208 281790
rect 42156 281726 42208 281732
rect 42168 281180 42196 281726
rect 42156 281104 42208 281110
rect 42156 281046 42208 281052
rect 42168 280568 42196 281046
rect 42156 279880 42208 279886
rect 42156 279822 42208 279828
rect 42168 279344 42196 279822
rect 42064 278656 42116 278662
rect 42064 278598 42116 278604
rect 42076 278188 42104 278598
rect 42156 277908 42208 277914
rect 42156 277850 42208 277856
rect 42168 277508 42196 277850
rect 42156 277432 42208 277438
rect 42156 277374 42208 277380
rect 42168 276896 42196 277374
rect 42064 276752 42116 276758
rect 42064 276694 42116 276700
rect 42076 276352 42104 276694
rect 42156 274304 42208 274310
rect 42156 274246 42208 274252
rect 42168 273836 42196 274246
rect 42720 273766 42748 283290
rect 42812 281790 42840 285738
rect 42984 285728 43036 285734
rect 42984 285670 43036 285676
rect 42892 285660 42944 285666
rect 42892 285602 42944 285608
rect 42800 281784 42852 281790
rect 42800 281726 42852 281732
rect 42904 274310 42932 285602
rect 42996 276758 43024 285670
rect 43088 279886 43116 293111
rect 43258 292768 43314 292777
rect 43258 292703 43314 292712
rect 43168 289876 43220 289882
rect 43168 289818 43220 289824
rect 43076 279880 43128 279886
rect 43076 279822 43128 279828
rect 43180 278662 43208 289818
rect 43168 278656 43220 278662
rect 43168 278598 43220 278604
rect 43272 277914 43300 292703
rect 43352 292052 43404 292058
rect 43352 291994 43404 292000
rect 43260 277908 43312 277914
rect 43260 277850 43312 277856
rect 42984 276752 43036 276758
rect 42984 276694 43036 276700
rect 42892 274304 42944 274310
rect 42892 274246 42944 274252
rect 42064 273760 42116 273766
rect 42064 273702 42116 273708
rect 42708 273760 42760 273766
rect 42708 273702 42760 273708
rect 42076 273224 42104 273702
rect 43364 272950 43392 291994
rect 42156 272944 42208 272950
rect 42156 272886 42208 272892
rect 43352 272944 43404 272950
rect 43352 272886 43404 272892
rect 42168 272544 42196 272886
rect 41970 272368 42026 272377
rect 41970 272303 42026 272312
rect 41984 272000 42012 272303
rect 42154 270464 42210 270473
rect 42154 270399 42210 270408
rect 42168 270164 42196 270399
rect 42154 270056 42210 270065
rect 42154 269991 42210 270000
rect 42168 269521 42196 269991
rect 42154 269376 42210 269385
rect 42154 269311 42210 269320
rect 42168 268872 42196 269311
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 41512 258392 41564 258398
rect 41510 258360 41512 258369
rect 41564 258360 41566 258369
rect 41510 258295 41566 258304
rect 41512 258052 41564 258058
rect 41512 257994 41564 258000
rect 41524 257961 41552 257994
rect 41510 257952 41566 257961
rect 41510 257887 41566 257896
rect 41512 257576 41564 257582
rect 41510 257544 41512 257553
rect 41564 257544 41566 257553
rect 41510 257479 41566 257488
rect 41788 256896 41840 256902
rect 41786 256864 41788 256873
rect 41840 256864 41842 256873
rect 41786 256799 41842 256808
rect 43456 256057 43484 298823
rect 44284 298081 44312 339895
rect 44376 339561 44404 340847
rect 44362 339552 44418 339561
rect 44362 339487 44418 339496
rect 44270 298072 44326 298081
rect 44270 298007 44326 298016
rect 44376 297265 44404 339487
rect 44362 297256 44418 297265
rect 44362 297191 44418 297200
rect 43536 291644 43588 291650
rect 43536 291586 43588 291592
rect 43548 277438 43576 291586
rect 45374 289912 45430 289921
rect 45374 289847 45430 289856
rect 43536 277432 43588 277438
rect 43536 277374 43588 277380
rect 43442 256048 43498 256057
rect 43442 255983 43498 255992
rect 43442 255640 43498 255649
rect 43442 255575 43498 255584
rect 42706 253600 42762 253609
rect 42706 253535 42762 253544
rect 31666 253056 31722 253065
rect 31666 252991 31722 253000
rect 31680 244322 31708 252991
rect 33046 251832 33102 251841
rect 33046 251767 33102 251776
rect 32770 250608 32826 250617
rect 32770 250543 32826 250552
rect 32784 245654 32812 250543
rect 32862 250200 32918 250209
rect 32862 250135 32918 250144
rect 32876 247602 32904 250135
rect 33060 249830 33088 251767
rect 33048 249824 33100 249830
rect 32954 249792 33010 249801
rect 33048 249766 33100 249772
rect 32954 249727 33010 249736
rect 32968 247738 32996 249727
rect 38290 248160 38346 248169
rect 38290 248095 38346 248104
rect 32968 247710 33088 247738
rect 32876 247574 32996 247602
rect 32784 245626 32904 245654
rect 31668 244316 31720 244322
rect 31668 244258 31720 244264
rect 32876 244254 32904 245626
rect 32968 244458 32996 247574
rect 32956 244452 33008 244458
rect 32956 244394 33008 244400
rect 33060 244390 33088 247710
rect 33048 244384 33100 244390
rect 33048 244326 33100 244332
rect 32864 244248 32916 244254
rect 32864 244190 32916 244196
rect 38304 242894 38332 248095
rect 41510 247752 41566 247761
rect 41510 247687 41512 247696
rect 41564 247687 41566 247696
rect 41512 247658 41564 247664
rect 41510 247344 41566 247353
rect 41510 247279 41512 247288
rect 41564 247279 41566 247288
rect 41512 247250 41564 247256
rect 41510 246528 41566 246537
rect 41510 246463 41512 246472
rect 41564 246463 41566 246472
rect 41512 246434 41564 246440
rect 42720 244526 42748 253535
rect 42798 252376 42854 252385
rect 42798 252311 42854 252320
rect 42708 244520 42760 244526
rect 42708 244462 42760 244468
rect 42708 244316 42760 244322
rect 42708 244258 42760 244264
rect 42432 243364 42484 243370
rect 42432 243306 42484 243312
rect 38292 242888 38344 242894
rect 38292 242830 38344 242836
rect 42444 240378 42472 243306
rect 42156 240372 42208 240378
rect 42156 240314 42208 240320
rect 42432 240372 42484 240378
rect 42432 240314 42484 240320
rect 42168 239836 42196 240314
rect 42720 238474 42748 244258
rect 42812 243030 42840 252311
rect 43258 249520 43314 249529
rect 43258 249455 43314 249464
rect 43166 248704 43222 248713
rect 43166 248639 43222 248648
rect 43076 244452 43128 244458
rect 43076 244394 43128 244400
rect 42892 244384 42944 244390
rect 42892 244326 42944 244332
rect 42800 243024 42852 243030
rect 42800 242966 42852 242972
rect 42800 242888 42852 242894
rect 42800 242830 42852 242836
rect 42156 238468 42208 238474
rect 42156 238410 42208 238416
rect 42708 238468 42760 238474
rect 42708 238410 42760 238416
rect 42168 238000 42196 238410
rect 42156 236700 42208 236706
rect 42156 236642 42208 236648
rect 42168 236164 42196 236642
rect 42812 235414 42840 242830
rect 42904 236706 42932 244326
rect 42984 244248 43036 244254
rect 42984 244190 43036 244196
rect 42892 236700 42944 236706
rect 42892 236642 42944 236648
rect 42156 235408 42208 235414
rect 42156 235350 42208 235356
rect 42800 235408 42852 235414
rect 42800 235350 42852 235356
rect 42168 234969 42196 235350
rect 42156 234660 42208 234666
rect 42156 234602 42208 234608
rect 42168 234328 42196 234602
rect 42156 234252 42208 234258
rect 42156 234194 42208 234200
rect 42168 233681 42196 234194
rect 42156 233368 42208 233374
rect 42156 233310 42208 233316
rect 42168 233104 42196 233310
rect 42156 231124 42208 231130
rect 42156 231066 42208 231072
rect 42168 230656 42196 231066
rect 42156 230580 42208 230586
rect 42156 230522 42208 230528
rect 42168 229976 42196 230522
rect 42996 229906 43024 244190
rect 43088 230586 43116 244394
rect 43180 234258 43208 248639
rect 43272 234666 43300 249455
rect 43350 249112 43406 249121
rect 43350 249047 43406 249056
rect 43364 243166 43392 249047
rect 43352 243160 43404 243166
rect 43352 243102 43404 243108
rect 43352 243024 43404 243030
rect 43352 242966 43404 242972
rect 43260 234660 43312 234666
rect 43260 234602 43312 234608
rect 43168 234252 43220 234258
rect 43168 234194 43220 234200
rect 43076 230580 43128 230586
rect 43076 230522 43128 230528
rect 42156 229900 42208 229906
rect 42156 229842 42208 229848
rect 42984 229900 43036 229906
rect 42984 229842 43036 229848
rect 42168 229364 42196 229842
rect 43364 229090 43392 242966
rect 42156 229084 42208 229090
rect 42156 229026 42208 229032
rect 43352 229084 43404 229090
rect 43352 229026 43404 229032
rect 42168 228820 42196 229026
rect 42064 227452 42116 227458
rect 42064 227394 42116 227400
rect 42076 226984 42104 227394
rect 42156 226840 42208 226846
rect 42156 226782 42208 226788
rect 42168 226304 42196 226782
rect 41970 225992 42026 226001
rect 41970 225927 42026 225936
rect 41984 225692 42012 225927
rect 41420 216776 41472 216782
rect 41420 216718 41472 216724
rect 31668 215824 31720 215830
rect 31668 215766 31720 215772
rect 29184 215756 29236 215762
rect 29184 215698 29236 215704
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 29196 204513 29224 215698
rect 29182 204504 29238 204513
rect 29182 204439 29238 204448
rect 31680 203697 31708 215766
rect 41432 214305 41460 216718
rect 41604 216708 41656 216714
rect 41604 216650 41656 216656
rect 41512 216640 41564 216646
rect 41512 216582 41564 216588
rect 41524 215121 41552 216582
rect 41510 215112 41566 215121
rect 41510 215047 41566 215056
rect 41616 214713 41644 216650
rect 41602 214704 41658 214713
rect 41602 214639 41658 214648
rect 41418 214296 41474 214305
rect 43456 214266 43484 255575
rect 43810 251560 43866 251569
rect 43810 251495 43866 251504
rect 43628 249824 43680 249830
rect 43628 249766 43680 249772
rect 43536 244520 43588 244526
rect 43536 244462 43588 244468
rect 43548 227458 43576 244462
rect 43640 243250 43668 249766
rect 43824 243370 43852 251495
rect 43902 251152 43958 251161
rect 43902 251087 43958 251096
rect 43812 243364 43864 243370
rect 43812 243306 43864 243312
rect 43640 243222 43760 243250
rect 43628 243160 43680 243166
rect 43628 243102 43680 243108
rect 43640 231130 43668 243102
rect 43732 233374 43760 243222
rect 43720 233368 43772 233374
rect 43720 233310 43772 233316
rect 43628 231124 43680 231130
rect 43628 231066 43680 231072
rect 43536 227452 43588 227458
rect 43536 227394 43588 227400
rect 43916 226846 43944 251087
rect 45388 230450 45416 289847
rect 45376 230444 45428 230450
rect 45376 230386 45428 230392
rect 43904 226840 43956 226846
rect 43904 226782 43956 226788
rect 41418 214231 41474 214240
rect 41512 214260 41564 214266
rect 41512 214202 41564 214208
rect 43444 214260 43496 214266
rect 43444 214202 43496 214208
rect 41420 213920 41472 213926
rect 41418 213888 41420 213897
rect 41472 213888 41474 213897
rect 41418 213823 41474 213832
rect 41524 213081 41552 214202
rect 41510 213072 41566 213081
rect 41510 213007 41566 213016
rect 45480 211313 45508 988042
rect 45744 988032 45796 988038
rect 45744 987974 45796 987980
rect 45560 987964 45612 987970
rect 45560 987906 45612 987912
rect 45572 213926 45600 987906
rect 45652 985040 45704 985046
rect 45652 984982 45704 984988
rect 45560 213920 45612 213926
rect 45560 213862 45612 213868
rect 45664 212129 45692 984982
rect 45756 254425 45784 987974
rect 48228 987420 48280 987426
rect 48228 987362 48280 987368
rect 45928 984972 45980 984978
rect 45928 984914 45980 984920
rect 45836 984904 45888 984910
rect 45836 984846 45888 984852
rect 45848 256902 45876 984846
rect 45836 256896 45888 256902
rect 45836 256838 45888 256844
rect 45940 255241 45968 984914
rect 46112 984632 46164 984638
rect 46112 984574 46164 984580
rect 46020 984156 46072 984162
rect 46020 984098 46072 984104
rect 46032 941526 46060 984098
rect 46020 941520 46072 941526
rect 46020 941462 46072 941468
rect 46020 932068 46072 932074
rect 46020 932010 46072 932016
rect 45926 255232 45982 255241
rect 45926 255167 45982 255176
rect 45742 254416 45798 254425
rect 45742 254351 45798 254360
rect 45928 247716 45980 247722
rect 45928 247658 45980 247664
rect 45836 247308 45888 247314
rect 45836 247250 45888 247256
rect 45744 246492 45796 246498
rect 45744 246434 45796 246440
rect 45756 230518 45784 246434
rect 45848 230586 45876 247250
rect 45940 230654 45968 247658
rect 45928 230648 45980 230654
rect 45928 230590 45980 230596
rect 45836 230580 45888 230586
rect 45836 230522 45888 230528
rect 45744 230512 45796 230518
rect 45744 230454 45796 230460
rect 46032 219706 46060 932010
rect 46124 298489 46152 984574
rect 46388 984496 46440 984502
rect 46388 984438 46440 984444
rect 46204 984428 46256 984434
rect 46204 984370 46256 984376
rect 46216 339969 46244 984370
rect 46296 762884 46348 762890
rect 46296 762826 46348 762832
rect 46202 339960 46258 339969
rect 46202 339895 46258 339904
rect 46204 332852 46256 332858
rect 46204 332794 46256 332800
rect 46110 298480 46166 298489
rect 46110 298415 46166 298424
rect 46110 290728 46166 290737
rect 46110 290663 46166 290672
rect 46124 230722 46152 290663
rect 46216 230858 46244 332794
rect 46204 230852 46256 230858
rect 46204 230794 46256 230800
rect 46112 230716 46164 230722
rect 46112 230658 46164 230664
rect 46020 219700 46072 219706
rect 46020 219642 46072 219648
rect 46308 219570 46336 762826
rect 46400 339561 46428 984438
rect 46478 684040 46534 684049
rect 46478 683975 46534 683984
rect 46386 339552 46442 339561
rect 46386 339487 46442 339496
rect 46386 291136 46442 291145
rect 46386 291071 46442 291080
rect 46400 230790 46428 291071
rect 46492 278594 46520 683975
rect 46570 598496 46626 598505
rect 46570 598431 46626 598440
rect 46480 278588 46532 278594
rect 46480 278530 46532 278536
rect 46584 278526 46612 598431
rect 46754 597680 46810 597689
rect 46754 597615 46810 597624
rect 46664 419484 46716 419490
rect 46664 419426 46716 419432
rect 46572 278520 46624 278526
rect 46572 278462 46624 278468
rect 46676 230994 46704 419426
rect 46768 278458 46796 597615
rect 46848 376100 46900 376106
rect 46848 376042 46900 376048
rect 46756 278452 46808 278458
rect 46756 278394 46808 278400
rect 46664 230988 46716 230994
rect 46664 230930 46716 230936
rect 46860 230926 46888 376042
rect 48240 297673 48268 987362
rect 62672 986876 62724 986882
rect 62672 986818 62724 986824
rect 62488 986808 62540 986814
rect 62488 986750 62540 986756
rect 62304 986740 62356 986746
rect 62304 986682 62356 986688
rect 48320 984564 48372 984570
rect 48320 984506 48372 984512
rect 48332 300121 48360 984506
rect 48412 984360 48464 984366
rect 48412 984302 48464 984308
rect 48424 345030 48452 984302
rect 62212 984088 62264 984094
rect 62212 984030 62264 984036
rect 62120 984020 62172 984026
rect 62120 983962 62172 983968
rect 62028 983952 62080 983958
rect 62028 983894 62080 983900
rect 58438 976032 58494 976041
rect 58438 975967 58494 975976
rect 58452 972942 58480 975967
rect 58440 972936 58492 972942
rect 58440 972878 58492 972884
rect 57978 962976 58034 962985
rect 57978 962911 58034 962920
rect 57992 960566 58020 962911
rect 48504 960560 48556 960566
rect 48504 960502 48556 960508
rect 57980 960560 58032 960566
rect 57980 960502 58032 960508
rect 48516 942750 48544 960502
rect 58438 949920 58494 949929
rect 58438 949855 58494 949864
rect 58452 949482 58480 949855
rect 58440 949476 58492 949482
rect 58440 949418 58492 949424
rect 49700 943084 49752 943090
rect 49700 943026 49752 943032
rect 48504 942744 48556 942750
rect 48504 942686 48556 942692
rect 49712 938398 49740 943026
rect 49700 938392 49752 938398
rect 49700 938334 49752 938340
rect 58440 938392 58492 938398
rect 58440 938334 58492 938340
rect 58452 937009 58480 938334
rect 58438 937000 58494 937009
rect 58438 936935 58494 936944
rect 58438 923808 58494 923817
rect 58438 923743 58494 923752
rect 58452 921874 58480 923743
rect 48596 921868 48648 921874
rect 48596 921810 48648 921816
rect 58440 921868 58492 921874
rect 58440 921810 58492 921816
rect 48504 805996 48556 806002
rect 48504 805938 48556 805944
rect 48412 345024 48464 345030
rect 48412 344966 48464 344972
rect 48412 336796 48464 336802
rect 48412 336738 48464 336744
rect 48318 300112 48374 300121
rect 48318 300047 48374 300056
rect 48226 297664 48282 297673
rect 48226 297599 48282 297608
rect 48424 258398 48452 336738
rect 48412 258392 48464 258398
rect 48412 258334 48464 258340
rect 46848 230920 46900 230926
rect 46848 230862 46900 230868
rect 46388 230784 46440 230790
rect 46388 230726 46440 230732
rect 48516 219774 48544 805938
rect 48608 800494 48636 921810
rect 59174 910752 59230 910761
rect 59174 910687 59230 910696
rect 59188 908138 59216 910687
rect 53840 908132 53892 908138
rect 53840 908074 53892 908080
rect 59176 908132 59228 908138
rect 59176 908074 59228 908080
rect 51080 883244 51132 883250
rect 51080 883186 51132 883192
rect 50988 869440 51040 869446
rect 50988 869382 51040 869388
rect 48688 858424 48740 858430
rect 48688 858366 48740 858372
rect 48596 800488 48648 800494
rect 48596 800430 48648 800436
rect 48596 778388 48648 778394
rect 48596 778330 48648 778336
rect 48608 730969 48636 778330
rect 48700 773974 48728 858366
rect 48780 844620 48832 844626
rect 48780 844562 48832 844568
rect 48792 774790 48820 844562
rect 48780 774784 48832 774790
rect 48780 774726 48832 774732
rect 48688 773968 48740 773974
rect 48688 773910 48740 773916
rect 48780 767372 48832 767378
rect 48780 767314 48832 767320
rect 48688 739764 48740 739770
rect 48688 739706 48740 739712
rect 48594 730960 48650 730969
rect 48594 730895 48650 730904
rect 48596 719636 48648 719642
rect 48596 719578 48648 719584
rect 48504 219768 48556 219774
rect 48504 219710 48556 219716
rect 48608 219638 48636 719578
rect 48700 688430 48728 739706
rect 48688 688424 48740 688430
rect 48688 688366 48740 688372
rect 48688 676660 48740 676666
rect 48688 676602 48740 676608
rect 48596 219632 48648 219638
rect 48596 219574 48648 219580
rect 46296 219564 46348 219570
rect 46296 219506 46348 219512
rect 48700 219502 48728 676602
rect 48792 670750 48820 767314
rect 51000 760578 51028 869382
rect 51092 817358 51120 883186
rect 51080 817352 51132 817358
rect 51080 817294 51132 817300
rect 53748 817148 53800 817154
rect 53748 817090 53800 817096
rect 51080 805996 51132 806002
rect 51080 805938 51132 805944
rect 50988 760572 51040 760578
rect 50988 760514 51040 760520
rect 51092 730561 51120 805938
rect 51264 792192 51316 792198
rect 51264 792134 51316 792140
rect 51276 731377 51304 792134
rect 51262 731368 51318 731377
rect 51262 731303 51318 731312
rect 51078 730552 51134 730561
rect 51078 730487 51134 730496
rect 51172 725960 51224 725966
rect 51172 725902 51224 725908
rect 50988 714876 51040 714882
rect 50988 714818 51040 714824
rect 48872 673532 48924 673538
rect 48872 673474 48924 673480
rect 48780 670744 48832 670750
rect 48780 670686 48832 670692
rect 48884 644570 48912 673474
rect 48964 662448 49016 662454
rect 48964 662390 49016 662396
rect 48872 644564 48924 644570
rect 48872 644506 48924 644512
rect 48872 634840 48924 634846
rect 48872 634782 48924 634788
rect 48780 633276 48832 633282
rect 48780 633218 48832 633224
rect 48688 219496 48740 219502
rect 48688 219438 48740 219444
rect 48792 219434 48820 633218
rect 48884 601934 48912 634782
rect 48872 601928 48924 601934
rect 48872 601870 48924 601876
rect 48872 590028 48924 590034
rect 48872 589970 48924 589976
rect 48884 231130 48912 589970
rect 48976 585206 49004 662390
rect 51000 629338 51028 714818
rect 51184 687750 51212 725902
rect 53760 716650 53788 817090
rect 53852 816921 53880 908074
rect 58438 897832 58494 897841
rect 58438 897767 58494 897776
rect 58452 897054 58480 897767
rect 53932 897048 53984 897054
rect 53932 896990 53984 896996
rect 58440 897048 58492 897054
rect 58440 896990 58492 896996
rect 53944 817698 53972 896990
rect 58438 884776 58494 884785
rect 58438 884711 58494 884720
rect 58452 883250 58480 884711
rect 58440 883244 58492 883250
rect 58440 883186 58492 883192
rect 58438 871720 58494 871729
rect 58438 871655 58494 871664
rect 58452 869446 58480 871655
rect 58440 869440 58492 869446
rect 58440 869382 58492 869388
rect 58438 858664 58494 858673
rect 58438 858599 58494 858608
rect 58452 858430 58480 858599
rect 58440 858424 58492 858430
rect 58440 858366 58492 858372
rect 58438 845608 58494 845617
rect 58438 845543 58494 845552
rect 58452 844626 58480 845543
rect 58440 844620 58492 844626
rect 58440 844562 58492 844568
rect 57978 832552 58034 832561
rect 57978 832487 58034 832496
rect 57992 830822 58020 832487
rect 54024 830816 54076 830822
rect 54024 830758 54076 830764
rect 57980 830816 58032 830822
rect 57980 830758 58032 830764
rect 53932 817692 53984 817698
rect 53932 817634 53984 817640
rect 53838 816912 53894 816921
rect 53838 816847 53894 816856
rect 54036 774450 54064 830758
rect 59174 819496 59230 819505
rect 59174 819431 59230 819440
rect 59188 817154 59216 819431
rect 59176 817148 59228 817154
rect 59176 817090 59228 817096
rect 58438 806576 58494 806585
rect 58438 806511 58494 806520
rect 58452 806002 58480 806511
rect 58440 805996 58492 806002
rect 58440 805938 58492 805944
rect 58070 793520 58126 793529
rect 58070 793455 58126 793464
rect 58084 792198 58112 793455
rect 58072 792192 58124 792198
rect 58072 792134 58124 792140
rect 58438 780464 58494 780473
rect 58438 780399 58494 780408
rect 58452 778394 58480 780399
rect 58440 778388 58492 778394
rect 58440 778330 58492 778336
rect 54024 774444 54076 774450
rect 54024 774386 54076 774392
rect 58438 767408 58494 767417
rect 58438 767343 58440 767352
rect 58492 767343 58494 767352
rect 58440 767314 58492 767320
rect 58346 754352 58402 754361
rect 58346 754287 58402 754296
rect 58360 753574 58388 754287
rect 53840 753568 53892 753574
rect 53840 753510 53892 753516
rect 58348 753568 58400 753574
rect 58348 753510 58400 753516
rect 53748 716644 53800 716650
rect 53748 716586 53800 716592
rect 53748 701072 53800 701078
rect 53748 701014 53800 701020
rect 51172 687744 51224 687750
rect 51172 687686 51224 687692
rect 51080 687268 51132 687274
rect 51080 687210 51132 687216
rect 51092 645182 51120 687210
rect 51080 645176 51132 645182
rect 51080 645118 51132 645124
rect 53760 644842 53788 701014
rect 53852 688090 53880 753510
rect 58438 741296 58494 741305
rect 58438 741231 58494 741240
rect 58452 739770 58480 741231
rect 58440 739764 58492 739770
rect 58440 739706 58492 739712
rect 58438 728240 58494 728249
rect 58438 728175 58494 728184
rect 58452 725966 58480 728175
rect 58440 725960 58492 725966
rect 58440 725902 58492 725908
rect 58438 715320 58494 715329
rect 58438 715255 58494 715264
rect 58452 714882 58480 715255
rect 58440 714876 58492 714882
rect 58440 714818 58492 714824
rect 58622 702264 58678 702273
rect 58622 702199 58678 702208
rect 58636 701078 58664 702199
rect 58624 701072 58676 701078
rect 58624 701014 58676 701020
rect 58438 689208 58494 689217
rect 58438 689143 58494 689152
rect 53840 688084 53892 688090
rect 53840 688026 53892 688032
rect 58452 687274 58480 689143
rect 58440 687268 58492 687274
rect 58440 687210 58492 687216
rect 58438 676152 58494 676161
rect 58438 676087 58494 676096
rect 58452 673538 58480 676087
rect 58440 673532 58492 673538
rect 58440 673474 58492 673480
rect 58438 663096 58494 663105
rect 58438 663031 58494 663040
rect 58452 662454 58480 663031
rect 58440 662448 58492 662454
rect 58440 662390 58492 662396
rect 59174 650040 59230 650049
rect 59174 649975 59230 649984
rect 59188 648650 59216 649975
rect 53840 648644 53892 648650
rect 53840 648586 53892 648592
rect 59176 648644 59228 648650
rect 59176 648586 59228 648592
rect 53748 644836 53800 644842
rect 53748 644778 53800 644784
rect 50988 629332 51040 629338
rect 50988 629274 51040 629280
rect 51080 623824 51132 623830
rect 51080 623766 51132 623772
rect 50988 610020 51040 610026
rect 50988 609962 51040 609968
rect 48964 585200 49016 585206
rect 48964 585142 49016 585148
rect 48964 582412 49016 582418
rect 48964 582354 49016 582360
rect 48976 558822 49004 582354
rect 48964 558816 49016 558822
rect 48964 558758 49016 558764
rect 49056 557592 49108 557598
rect 49056 557534 49108 557540
rect 48964 546916 49016 546922
rect 48964 546858 49016 546864
rect 48872 231124 48924 231130
rect 48872 231066 48924 231072
rect 48976 231062 49004 546858
rect 49068 410718 49096 557534
rect 51000 541754 51028 609962
rect 51092 601361 51120 623766
rect 51078 601352 51134 601361
rect 51078 601287 51134 601296
rect 53852 600953 53880 648586
rect 58438 637120 58494 637129
rect 58438 637055 58494 637064
rect 58452 634846 58480 637055
rect 58440 634840 58492 634846
rect 58440 634782 58492 634788
rect 58438 624064 58494 624073
rect 58438 623999 58494 624008
rect 58452 623830 58480 623999
rect 58440 623824 58492 623830
rect 58440 623766 58492 623772
rect 58438 611008 58494 611017
rect 58438 610943 58494 610952
rect 58452 610026 58480 610943
rect 58440 610020 58492 610026
rect 58440 609962 58492 609968
rect 53838 600944 53894 600953
rect 53838 600879 53894 600888
rect 59174 597952 59230 597961
rect 59174 597887 59230 597896
rect 59188 596222 59216 597887
rect 53748 596216 53800 596222
rect 53748 596158 53800 596164
rect 59176 596216 59228 596222
rect 59176 596158 59228 596164
rect 53760 558550 53788 596158
rect 58438 584896 58494 584905
rect 58438 584831 58494 584840
rect 58452 582418 58480 584831
rect 58440 582412 58492 582418
rect 58440 582354 58492 582360
rect 58438 571840 58494 571849
rect 58438 571775 58494 571784
rect 58346 558784 58402 558793
rect 58346 558719 58402 558728
rect 53748 558544 53800 558550
rect 53748 558486 53800 558492
rect 58360 557598 58388 558719
rect 58452 558482 58480 571775
rect 58440 558476 58492 558482
rect 58440 558418 58492 558424
rect 58348 557592 58400 557598
rect 58348 557534 58400 557540
rect 58346 545864 58402 545873
rect 58346 545799 58402 545808
rect 58360 543794 58388 545799
rect 53840 543788 53892 543794
rect 53840 543730 53892 543736
rect 58348 543788 58400 543794
rect 58348 543730 58400 543736
rect 50988 541748 51040 541754
rect 50988 541690 51040 541696
rect 51264 518968 51316 518974
rect 51264 518910 51316 518916
rect 50988 505164 51040 505170
rect 50988 505106 51040 505112
rect 49148 491360 49200 491366
rect 49148 491302 49200 491308
rect 49056 410712 49108 410718
rect 49056 410654 49108 410660
rect 49056 400240 49108 400246
rect 49056 400182 49108 400188
rect 49068 281110 49096 400182
rect 49160 387190 49188 491302
rect 49240 414044 49292 414050
rect 49240 413986 49292 413992
rect 49148 387184 49200 387190
rect 49148 387126 49200 387132
rect 49148 375420 49200 375426
rect 49148 375362 49200 375368
rect 49160 301646 49188 375362
rect 49252 344350 49280 413986
rect 51000 366858 51028 505106
rect 51172 480276 51224 480282
rect 51172 480218 51224 480224
rect 51080 438932 51132 438938
rect 51080 438874 51132 438880
rect 50988 366852 51040 366858
rect 50988 366794 51040 366800
rect 50988 347812 51040 347818
rect 50988 347754 51040 347760
rect 49240 344344 49292 344350
rect 49240 344286 49292 344292
rect 49148 301640 49200 301646
rect 49148 301582 49200 301588
rect 49056 281104 49108 281110
rect 49056 281046 49108 281052
rect 51000 257582 51028 347754
rect 51092 343942 51120 438874
rect 51184 388006 51212 480218
rect 51276 430545 51304 518910
rect 53748 452668 53800 452674
rect 53748 452610 53800 452616
rect 51262 430536 51318 430545
rect 51262 430471 51318 430480
rect 51172 388000 51224 388006
rect 51172 387942 51224 387948
rect 51172 361616 51224 361622
rect 51172 361558 51224 361564
rect 51080 343936 51132 343942
rect 51080 343878 51132 343884
rect 51184 300966 51212 361558
rect 53760 320142 53788 452610
rect 53852 430137 53880 543730
rect 59266 532808 59322 532817
rect 59266 532743 59322 532752
rect 58438 519752 58494 519761
rect 58438 519687 58494 519696
rect 58452 518974 58480 519687
rect 58440 518968 58492 518974
rect 58440 518910 58492 518916
rect 58438 506696 58494 506705
rect 58438 506631 58494 506640
rect 58452 505170 58480 506631
rect 58440 505164 58492 505170
rect 58440 505106 58492 505112
rect 57978 493640 58034 493649
rect 57978 493575 58034 493584
rect 57992 491366 58020 493575
rect 57980 491360 58032 491366
rect 57980 491302 58032 491308
rect 58438 480584 58494 480593
rect 58438 480519 58494 480528
rect 58452 480282 58480 480519
rect 58440 480276 58492 480282
rect 58440 480218 58492 480224
rect 58714 467528 58770 467537
rect 58714 467463 58770 467472
rect 58728 466478 58756 467463
rect 54024 466472 54076 466478
rect 54024 466414 54076 466420
rect 58716 466472 58768 466478
rect 58716 466414 58768 466420
rect 53838 430128 53894 430137
rect 53838 430063 53894 430072
rect 53932 427916 53984 427922
rect 53932 427858 53984 427864
rect 53840 389224 53892 389230
rect 53840 389166 53892 389172
rect 53748 320136 53800 320142
rect 53748 320078 53800 320084
rect 51172 300960 51224 300966
rect 51172 300902 51224 300908
rect 53852 300529 53880 389166
rect 53944 344486 53972 427858
rect 54036 387666 54064 466414
rect 59174 454608 59230 454617
rect 59174 454543 59230 454552
rect 59188 452674 59216 454543
rect 59176 452668 59228 452674
rect 59176 452610 59228 452616
rect 58438 441552 58494 441561
rect 58438 441487 58494 441496
rect 58452 438938 58480 441487
rect 58440 438932 58492 438938
rect 58440 438874 58492 438880
rect 59280 430846 59308 532743
rect 59268 430840 59320 430846
rect 59268 430782 59320 430788
rect 58254 428496 58310 428505
rect 58254 428431 58310 428440
rect 58268 427922 58296 428431
rect 58256 427916 58308 427922
rect 58256 427858 58308 427864
rect 58438 415440 58494 415449
rect 58438 415375 58494 415384
rect 58452 414050 58480 415375
rect 58440 414044 58492 414050
rect 58440 413986 58492 413992
rect 58438 402384 58494 402393
rect 58438 402319 58494 402328
rect 58452 400246 58480 402319
rect 58440 400240 58492 400246
rect 58440 400182 58492 400188
rect 57978 389328 58034 389337
rect 57978 389263 58034 389272
rect 57992 389230 58020 389263
rect 57980 389224 58032 389230
rect 57980 389166 58032 389172
rect 54024 387660 54076 387666
rect 54024 387602 54076 387608
rect 62040 383081 62068 983894
rect 62132 386345 62160 983962
rect 62118 386336 62174 386345
rect 62118 386271 62174 386280
rect 62224 383489 62252 984030
rect 62316 939457 62344 986682
rect 62396 985380 62448 985386
rect 62396 985322 62448 985328
rect 62302 939448 62358 939457
rect 62302 939383 62358 939392
rect 62304 817080 62356 817086
rect 62304 817022 62356 817028
rect 62210 383480 62266 383489
rect 62210 383415 62266 383424
rect 62026 383072 62082 383081
rect 62026 383007 62082 383016
rect 58438 376272 58494 376281
rect 58438 376207 58494 376216
rect 58452 375426 58480 376207
rect 58440 375420 58492 375426
rect 58440 375362 58492 375368
rect 58438 363352 58494 363361
rect 58438 363287 58494 363296
rect 58452 361622 58480 363287
rect 58440 361616 58492 361622
rect 58440 361558 58492 361564
rect 58438 350296 58494 350305
rect 58438 350231 58494 350240
rect 58452 347818 58480 350231
rect 58440 347812 58492 347818
rect 58440 347754 58492 347760
rect 53932 344480 53984 344486
rect 53932 344422 53984 344428
rect 58438 337240 58494 337249
rect 58438 337175 58494 337184
rect 58452 336802 58480 337175
rect 58440 336796 58492 336802
rect 58440 336738 58492 336744
rect 58162 324184 58218 324193
rect 58162 324119 58218 324128
rect 58176 323542 58204 324119
rect 53932 323536 53984 323542
rect 53932 323478 53984 323484
rect 58164 323536 58216 323542
rect 58164 323478 58216 323484
rect 53838 300520 53894 300529
rect 53838 300455 53894 300464
rect 53944 258058 53972 323478
rect 59266 311128 59322 311137
rect 59266 311063 59322 311072
rect 53932 258052 53984 258058
rect 53932 257994 53984 258000
rect 50988 257576 51040 257582
rect 50988 257518 51040 257524
rect 52276 256760 52328 256766
rect 52276 256702 52328 256708
rect 52184 245676 52236 245682
rect 52184 245618 52236 245624
rect 52092 237448 52144 237454
rect 52092 237390 52144 237396
rect 48964 231056 49016 231062
rect 48964 230998 49016 231004
rect 48780 219428 48832 219434
rect 48780 219370 48832 219376
rect 46940 218068 46992 218074
rect 46940 218010 46992 218016
rect 46952 212537 46980 218010
rect 48228 215892 48280 215898
rect 48228 215834 48280 215840
rect 46938 212528 46994 212537
rect 46938 212463 46994 212472
rect 45650 212120 45706 212129
rect 45650 212055 45706 212064
rect 45466 211304 45522 211313
rect 45466 211239 45522 211248
rect 32954 209808 33010 209817
rect 32954 209743 33010 209752
rect 31666 203688 31722 203697
rect 31666 203623 31722 203632
rect 32968 200054 32996 209743
rect 33046 208176 33102 208185
rect 33046 208111 33102 208120
rect 33060 200258 33088 208111
rect 42890 206816 42946 206825
rect 42890 206751 42946 206760
rect 42798 205184 42854 205193
rect 42798 205119 42854 205128
rect 33048 200252 33100 200258
rect 33048 200194 33100 200200
rect 41880 200252 41932 200258
rect 41880 200194 41932 200200
rect 32956 200048 33008 200054
rect 32956 199990 33008 199996
rect 41892 197470 41920 200194
rect 42524 200048 42576 200054
rect 42524 199990 42576 199996
rect 41880 197464 41932 197470
rect 41880 197406 41932 197412
rect 41880 197192 41932 197198
rect 41880 197134 41932 197140
rect 41892 196656 41920 197134
rect 42536 195294 42564 199990
rect 42156 195288 42208 195294
rect 42156 195230 42208 195236
rect 42524 195288 42576 195294
rect 42524 195230 42576 195236
rect 42168 194820 42196 195230
rect 42064 193520 42116 193526
rect 42064 193462 42116 193468
rect 42076 192984 42104 193462
rect 42812 192234 42840 205119
rect 42904 193526 42932 206751
rect 43074 206408 43130 206417
rect 43074 206343 43130 206352
rect 42982 205592 43038 205601
rect 42982 205527 43038 205536
rect 42892 193520 42944 193526
rect 42892 193462 42944 193468
rect 42156 192228 42208 192234
rect 42156 192170 42208 192176
rect 42800 192228 42852 192234
rect 42800 192170 42852 192176
rect 42168 191760 42196 192170
rect 42064 191480 42116 191486
rect 42064 191422 42116 191428
rect 42076 191148 42104 191422
rect 42996 191010 43024 205527
rect 43088 191486 43116 206343
rect 48240 204785 48268 215834
rect 48226 204776 48282 204785
rect 48226 204711 48282 204720
rect 43076 191480 43128 191486
rect 43076 191422 43128 191428
rect 42156 191004 42208 191010
rect 42156 190946 42208 190952
rect 42984 191004 43036 191010
rect 42984 190946 43036 190952
rect 42168 190468 42196 190946
rect 42154 190224 42210 190233
rect 42154 190159 42210 190168
rect 42168 189924 42196 190159
rect 41878 187640 41934 187649
rect 41878 187575 41934 187584
rect 41892 187445 41920 187575
rect 42154 187096 42210 187105
rect 42154 187031 42210 187040
rect 42168 186796 42196 187031
rect 41970 186416 42026 186425
rect 41970 186351 42026 186360
rect 41984 186184 42012 186351
rect 42154 185872 42210 185881
rect 42154 185807 42210 185816
rect 42168 185605 42196 185807
rect 42154 184240 42210 184249
rect 42154 184175 42210 184184
rect 42168 183765 42196 184175
rect 41786 183696 41842 183705
rect 41786 183631 41842 183640
rect 41800 183124 41828 183631
rect 41786 182744 41842 182753
rect 41786 182679 41842 182688
rect 41800 182477 41828 182679
rect 52104 51066 52132 237390
rect 52092 51060 52144 51066
rect 52092 51002 52144 51008
rect 52196 42906 52224 245618
rect 52288 47122 52316 256702
rect 57610 227760 57666 227769
rect 52736 227724 52788 227730
rect 57610 227695 57666 227704
rect 52736 227666 52788 227672
rect 52748 217410 52776 227666
rect 56046 227624 56102 227633
rect 56046 227559 56102 227568
rect 55126 225040 55182 225049
rect 55126 224975 55182 224984
rect 53564 222420 53616 222426
rect 53564 222362 53616 222368
rect 53576 217410 53604 222362
rect 54390 222184 54446 222193
rect 54390 222119 54446 222128
rect 54404 217410 54432 222119
rect 55140 217410 55168 224975
rect 56060 217410 56088 227559
rect 56874 224904 56930 224913
rect 56874 224839 56930 224848
rect 56888 217410 56916 224839
rect 57624 217410 57652 227695
rect 59176 222216 59228 222222
rect 59176 222158 59228 222164
rect 58624 219836 58676 219842
rect 58624 219778 58676 219784
rect 58636 217410 58664 219778
rect 59188 217410 59216 222158
rect 52440 217382 52776 217410
rect 53268 217382 53604 217410
rect 54096 217382 54432 217410
rect 54924 217382 55168 217410
rect 55752 217382 56088 217410
rect 56580 217382 56916 217410
rect 57408 217382 57652 217410
rect 58328 217382 58664 217410
rect 59156 217382 59216 217410
rect 59280 216782 59308 311063
rect 59358 298208 59414 298217
rect 59358 298143 59414 298152
rect 59268 216776 59320 216782
rect 59268 216718 59320 216724
rect 59372 216646 59400 298143
rect 59450 285152 59506 285161
rect 59450 285087 59506 285096
rect 59464 216714 59492 285087
rect 62316 278361 62344 817022
rect 62408 772818 62436 985322
rect 62500 938505 62528 986750
rect 62580 983136 62632 983142
rect 62580 983078 62632 983084
rect 62486 938496 62542 938505
rect 62486 938431 62542 938440
rect 62488 817012 62540 817018
rect 62488 816954 62540 816960
rect 62396 772812 62448 772818
rect 62396 772754 62448 772760
rect 62396 728748 62448 728754
rect 62396 728690 62448 728696
rect 62302 278352 62358 278361
rect 62302 278287 62358 278296
rect 62408 278186 62436 728690
rect 62396 278180 62448 278186
rect 62396 278122 62448 278128
rect 62500 278089 62528 816954
rect 62592 596193 62620 983078
rect 62684 950842 62712 986818
rect 62856 985448 62908 985454
rect 62856 985390 62908 985396
rect 62764 983068 62816 983074
rect 62764 983010 62816 983016
rect 62672 950836 62724 950842
rect 62672 950778 62724 950784
rect 62672 814292 62724 814298
rect 62672 814234 62724 814240
rect 62578 596184 62634 596193
rect 62578 596119 62634 596128
rect 62578 430672 62634 430681
rect 62578 430607 62634 430616
rect 62592 278390 62620 430607
rect 62580 278384 62632 278390
rect 62580 278326 62632 278332
rect 62684 278225 62712 814234
rect 62776 598942 62804 983010
rect 62868 814201 62896 985390
rect 73448 983620 73476 989402
rect 89640 983620 89668 990762
rect 92972 989466 93000 1004702
rect 98274 1004663 98276 1004672
rect 98328 1004663 98330 1004672
rect 99102 1004728 99158 1004737
rect 99102 1004663 99104 1004672
rect 98276 1004634 98328 1004640
rect 99156 1004663 99158 1004672
rect 105634 1004728 105636 1004737
rect 105688 1004728 105690 1004737
rect 105634 1004663 105690 1004672
rect 125508 1004692 125560 1004698
rect 99104 1004634 99156 1004640
rect 125508 1004634 125560 1004640
rect 118700 999932 118752 999938
rect 118700 999874 118752 999880
rect 104348 999864 104400 999870
rect 102782 999832 102838 999841
rect 93052 999796 93104 999802
rect 102782 999767 102784 999776
rect 93052 999738 93104 999744
rect 102836 999767 102838 999776
rect 104346 999832 104348 999841
rect 104400 999832 104402 999841
rect 104346 999767 104402 999776
rect 102784 999738 102836 999744
rect 93064 999190 93092 999738
rect 100668 999728 100720 999734
rect 100666 999696 100668 999705
rect 100720 999696 100722 999705
rect 100666 999631 100722 999640
rect 102322 999696 102378 999705
rect 102322 999631 102324 999640
rect 102376 999631 102378 999640
rect 102324 999602 102376 999608
rect 101956 999592 102008 999598
rect 101494 999560 101550 999569
rect 95148 999524 95200 999530
rect 101494 999495 101496 999504
rect 95148 999466 95200 999472
rect 101548 999495 101550 999504
rect 101954 999560 101956 999569
rect 102008 999560 102010 999569
rect 101954 999495 102010 999504
rect 101496 999466 101548 999472
rect 93052 999184 93104 999190
rect 93052 999126 93104 999132
rect 95160 995353 95188 999466
rect 97908 999456 97960 999462
rect 103152 999456 103204 999462
rect 97908 999398 97960 999404
rect 99470 999424 99526 999433
rect 95700 999320 95752 999326
rect 95700 999262 95752 999268
rect 95332 999252 95384 999258
rect 95332 999194 95384 999200
rect 95344 995489 95372 999194
rect 95516 999184 95568 999190
rect 95516 999126 95568 999132
rect 95528 995625 95556 999126
rect 95712 996441 95740 999262
rect 95698 996432 95754 996441
rect 95698 996367 95754 996376
rect 95514 995616 95570 995625
rect 95514 995551 95570 995560
rect 97354 995616 97410 995625
rect 97354 995551 97410 995560
rect 95330 995480 95386 995489
rect 95330 995415 95386 995424
rect 95146 995344 95202 995353
rect 95146 995279 95202 995288
rect 97368 993857 97396 995551
rect 97920 994129 97948 999398
rect 99470 999359 99472 999368
rect 99524 999359 99526 999368
rect 103150 999424 103152 999433
rect 103204 999424 103206 999433
rect 103150 999359 103206 999368
rect 99472 999330 99524 999336
rect 101128 999320 101180 999326
rect 100298 999288 100354 999297
rect 100298 999223 100300 999232
rect 100352 999223 100354 999232
rect 101126 999288 101128 999297
rect 101180 999288 101182 999297
rect 101126 999223 101182 999232
rect 100300 999194 100352 999200
rect 99932 999184 99984 999190
rect 99930 999152 99932 999161
rect 99984 999152 99986 999161
rect 118712 999122 118740 999874
rect 99930 999087 99986 999096
rect 118700 999116 118752 999122
rect 118700 999058 118752 999064
rect 122104 999116 122156 999122
rect 122104 999058 122156 999064
rect 107658 997248 107714 997257
rect 107658 997183 107660 997192
rect 107712 997183 107714 997192
rect 115938 997248 115994 997257
rect 115938 997183 115940 997192
rect 107660 997154 107712 997160
rect 115992 997183 115994 997192
rect 115940 997154 115992 997160
rect 108486 996160 108542 996169
rect 108486 996095 108488 996104
rect 108540 996095 108542 996104
rect 113364 996124 113416 996130
rect 108488 996066 108540 996072
rect 113364 996066 113416 996072
rect 113270 995888 113326 995897
rect 113270 995823 113326 995832
rect 110418 995752 110474 995761
rect 110418 995687 110474 995696
rect 104162 995616 104218 995625
rect 104162 995551 104218 995560
rect 104346 995616 104402 995625
rect 104346 995551 104402 995560
rect 97906 994120 97962 994129
rect 97906 994055 97962 994064
rect 97354 993848 97410 993857
rect 97354 993783 97410 993792
rect 104176 993682 104204 995551
rect 104360 993721 104388 995551
rect 104346 993712 104402 993721
rect 104164 993676 104216 993682
rect 104346 993647 104402 993656
rect 104164 993618 104216 993624
rect 92960 989460 93012 989466
rect 92960 989402 93012 989408
rect 105820 989460 105872 989466
rect 105820 989402 105872 989408
rect 105832 983620 105860 989402
rect 110432 984162 110460 995687
rect 110510 995616 110566 995625
rect 110510 995551 110566 995560
rect 110524 986814 110552 995551
rect 110602 995480 110658 995489
rect 110602 995415 110658 995424
rect 110512 986808 110564 986814
rect 110512 986750 110564 986756
rect 110616 986746 110644 995415
rect 113284 989466 113312 995823
rect 113272 989460 113324 989466
rect 113272 989402 113324 989408
rect 113376 986882 113404 996066
rect 113364 986876 113416 986882
rect 113364 986818 113416 986824
rect 110604 986740 110656 986746
rect 110604 986682 110656 986688
rect 110420 984156 110472 984162
rect 110420 984098 110472 984104
rect 122116 983620 122144 999058
rect 125520 986950 125548 1004634
rect 125612 996193 125640 1005110
rect 143814 1005071 143870 1005080
rect 143722 1005000 143778 1005009
rect 143644 1004958 143722 1004986
rect 125692 1004828 125744 1004834
rect 125692 1004770 125744 1004776
rect 125600 996187 125652 996193
rect 125600 996129 125652 996135
rect 125704 996125 125732 1004770
rect 125784 1004760 125836 1004766
rect 125784 1004702 125836 1004708
rect 125692 996119 125744 996125
rect 125692 996061 125744 996067
rect 125796 996057 125824 1004702
rect 125784 996051 125836 996057
rect 125784 995993 125836 995999
rect 143644 995858 143672 1004958
rect 143722 1004935 143778 1004944
rect 143828 1004714 143856 1005071
rect 143736 1004686 143856 1004714
rect 143736 995920 143764 1004686
rect 143908 1001904 143960 1001910
rect 143908 1001846 143960 1001852
rect 143816 999184 143868 999190
rect 143816 999126 143868 999132
rect 143724 995914 143776 995920
rect 136272 995852 136324 995858
rect 136272 995794 136324 995800
rect 136824 995852 136876 995858
rect 136824 995794 136876 995800
rect 137928 995852 137980 995858
rect 137928 995794 137980 995800
rect 143632 995852 143684 995858
rect 143724 995856 143776 995862
rect 143632 995794 143684 995800
rect 136284 995738 136312 995794
rect 136836 995738 136864 995794
rect 137940 995738 137968 995794
rect 143828 995790 143856 999126
rect 139216 995784 139268 995790
rect 135930 995710 136312 995738
rect 136482 995710 136864 995738
rect 137770 995710 137968 995738
rect 138966 995732 139216 995738
rect 143816 995784 143868 995790
rect 142802 995752 142858 995761
rect 138966 995726 139268 995732
rect 138966 995710 139256 995726
rect 140806 995722 141096 995738
rect 140806 995716 141108 995722
rect 140806 995710 141056 995716
rect 142646 995710 142802 995738
rect 143816 995726 143868 995732
rect 142802 995687 142858 995696
rect 141056 995658 141108 995664
rect 143920 995654 143948 1001846
rect 144000 999116 144052 999122
rect 144000 999058 144052 999064
rect 144012 997257 144040 999058
rect 144092 997756 144144 997762
rect 144092 997698 144144 997704
rect 143998 997248 144054 997257
rect 143998 997183 144054 997192
rect 144000 997144 144052 997150
rect 144000 997086 144052 997092
rect 133144 995648 133196 995654
rect 132158 995586 132448 995602
rect 132802 995596 133144 995602
rect 143908 995648 143960 995654
rect 137374 995616 137430 995625
rect 132802 995590 133196 995596
rect 132158 995580 132460 995586
rect 132158 995574 132408 995580
rect 132802 995574 133184 995590
rect 137126 995574 137374 995602
rect 143908 995590 143960 995596
rect 137374 995551 137430 995560
rect 132408 995522 132460 995528
rect 130016 995512 130068 995518
rect 129766 995460 130016 995466
rect 144012 995489 144040 997086
rect 144104 995518 144132 997698
rect 144092 995512 144144 995518
rect 133694 995480 133750 995489
rect 129766 995454 130068 995460
rect 128464 993682 128492 995452
rect 129108 993750 129136 995452
rect 129766 995438 130056 995454
rect 131606 995450 131896 995466
rect 131606 995444 131908 995450
rect 131606 995438 131856 995444
rect 133446 995438 133694 995466
rect 143998 995480 144054 995489
rect 140162 995438 140544 995466
rect 133694 995415 133750 995424
rect 131856 995386 131908 995392
rect 140516 993750 140544 995438
rect 144092 995454 144144 995460
rect 143998 995415 144054 995424
rect 129096 993744 129148 993750
rect 129096 993686 129148 993692
rect 140504 993744 140556 993750
rect 140504 993686 140556 993692
rect 128452 993676 128504 993682
rect 128452 993618 128504 993624
rect 144840 988786 144868 1005450
rect 145104 1005440 145156 1005446
rect 145104 1005382 145156 1005388
rect 145012 1005372 145064 1005378
rect 145012 1005314 145064 1005320
rect 144920 1005304 144972 1005310
rect 144920 1005246 144972 1005252
rect 144932 995586 144960 1005246
rect 144920 995580 144972 995586
rect 144920 995522 144972 995528
rect 145024 993818 145052 1005314
rect 145116 995450 145144 1005382
rect 145208 995989 145236 1007422
rect 154578 1007383 154634 1007392
rect 501328 1007412 501380 1007418
rect 501328 1007354 501380 1007360
rect 517336 1007412 517388 1007418
rect 517336 1007354 517388 1007360
rect 501340 1007321 501368 1007354
rect 501326 1007312 501382 1007321
rect 501326 1007247 501382 1007256
rect 424690 1006088 424746 1006097
rect 424690 1006023 424692 1006032
rect 424744 1006023 424746 1006032
rect 466460 1006052 466512 1006058
rect 424692 1005994 424744 1006000
rect 466460 1005994 466512 1006000
rect 423862 1005952 423918 1005961
rect 423862 1005887 423864 1005896
rect 423916 1005887 423918 1005896
rect 440148 1005916 440200 1005922
rect 423864 1005858 423916 1005864
rect 440148 1005858 440200 1005864
rect 424324 1005848 424376 1005854
rect 424322 1005816 424324 1005825
rect 424376 1005816 424378 1005825
rect 424322 1005751 424378 1005760
rect 356060 1005712 356112 1005718
rect 356058 1005680 356060 1005689
rect 374276 1005712 374328 1005718
rect 356112 1005680 356114 1005689
rect 356058 1005615 356114 1005624
rect 356518 1005680 356574 1005689
rect 374276 1005654 374328 1005660
rect 356518 1005615 356520 1005624
rect 356572 1005615 356574 1005624
rect 356520 1005586 356572 1005592
rect 200028 1005576 200080 1005582
rect 160282 1005544 160338 1005553
rect 207204 1005576 207256 1005582
rect 200028 1005518 200080 1005524
rect 207202 1005544 207204 1005553
rect 207256 1005544 207258 1005553
rect 160282 1005479 160284 1005488
rect 160336 1005479 160338 1005488
rect 195336 1005508 195388 1005514
rect 160284 1005450 160336 1005456
rect 195336 1005450 195388 1005456
rect 154948 1005440 155000 1005446
rect 153750 1005408 153806 1005417
rect 153750 1005343 153752 1005352
rect 153804 1005343 153806 1005352
rect 154946 1005408 154948 1005417
rect 155000 1005408 155002 1005417
rect 154946 1005343 155002 1005352
rect 153752 1005314 153804 1005320
rect 153292 1005304 153344 1005310
rect 151266 1005272 151322 1005281
rect 148876 1005236 148928 1005242
rect 151266 1005207 151268 1005216
rect 148876 1005178 148928 1005184
rect 151320 1005207 151322 1005216
rect 153290 1005272 153292 1005281
rect 153344 1005272 153346 1005281
rect 153290 1005207 153346 1005216
rect 151268 1005178 151320 1005184
rect 148888 1005145 148916 1005178
rect 148874 1005136 148930 1005145
rect 148874 1005071 148930 1005080
rect 149702 1005136 149758 1005145
rect 149702 1005071 149704 1005080
rect 149756 1005071 149758 1005080
rect 150438 1005136 150494 1005145
rect 150438 1005071 150440 1005080
rect 149704 1005042 149756 1005048
rect 150492 1005071 150494 1005080
rect 175188 1005100 175240 1005106
rect 150440 1005042 150492 1005048
rect 175188 1005042 175240 1005048
rect 148876 1005032 148928 1005038
rect 148874 1005000 148876 1005009
rect 150900 1005032 150952 1005038
rect 148928 1005000 148930 1005009
rect 148140 1004964 148192 1004970
rect 148874 1004935 148930 1004944
rect 150898 1005000 150900 1005009
rect 150952 1005000 150954 1005009
rect 150898 1004935 150954 1004944
rect 154118 1005000 154174 1005009
rect 154118 1004935 154120 1004944
rect 148140 1004906 148192 1004912
rect 154172 1004935 154174 1004944
rect 159454 1005000 159510 1005009
rect 159454 1004935 159456 1004944
rect 154120 1004906 154172 1004912
rect 159508 1004935 159510 1004944
rect 173900 1004964 173952 1004970
rect 159456 1004906 159508 1004912
rect 173900 1004906 173952 1004912
rect 147586 1004864 147642 1004873
rect 147586 1004799 147642 1004808
rect 145196 995983 145248 995989
rect 145196 995925 145248 995931
rect 147600 995625 147628 1004799
rect 147770 1004728 147826 1004737
rect 147770 1004663 147826 1004672
rect 147784 997150 147812 1004663
rect 147772 997144 147824 997150
rect 147772 997086 147824 997092
rect 148152 996441 148180 1004906
rect 148876 1004896 148928 1004902
rect 148874 1004864 148876 1004873
rect 152096 1004896 152148 1004902
rect 148928 1004864 148930 1004873
rect 148784 1004828 148836 1004834
rect 148874 1004799 148930 1004808
rect 152094 1004864 152096 1004873
rect 152148 1004864 152150 1004873
rect 152094 1004799 152150 1004808
rect 152922 1004864 152978 1004873
rect 152922 1004799 152924 1004808
rect 148784 1004770 148836 1004776
rect 152976 1004799 152978 1004808
rect 156970 1004864 157026 1004873
rect 156970 1004799 156972 1004808
rect 152924 1004770 152976 1004776
rect 157024 1004799 157026 1004808
rect 156972 1004770 157024 1004776
rect 148796 1001910 148824 1004770
rect 148876 1004760 148928 1004766
rect 148874 1004728 148876 1004737
rect 151728 1004760 151780 1004766
rect 148928 1004728 148930 1004737
rect 151726 1004728 151728 1004737
rect 157800 1004760 157852 1004766
rect 151780 1004728 151782 1004737
rect 148874 1004663 148930 1004672
rect 148968 1004692 149020 1004698
rect 151726 1004663 151782 1004672
rect 152554 1004728 152610 1004737
rect 157798 1004728 157800 1004737
rect 157852 1004728 157854 1004737
rect 152554 1004663 152556 1004672
rect 148968 1004634 149020 1004640
rect 152608 1004663 152610 1004672
rect 154488 1004692 154540 1004698
rect 152556 1004634 152608 1004640
rect 157798 1004663 157854 1004672
rect 160650 1004728 160706 1004737
rect 160650 1004663 160652 1004672
rect 154488 1004634 154540 1004640
rect 160704 1004663 160706 1004672
rect 160652 1004634 160704 1004640
rect 148784 1001904 148836 1001910
rect 148784 1001846 148836 1001852
rect 148980 999190 149008 1004634
rect 148968 999184 149020 999190
rect 148968 999126 149020 999132
rect 154120 999184 154172 999190
rect 154120 999126 154172 999132
rect 148138 996432 148194 996441
rect 148138 996367 148194 996376
rect 154132 995722 154160 999126
rect 154120 995716 154172 995722
rect 154120 995658 154172 995664
rect 147586 995616 147642 995625
rect 147586 995551 147642 995560
rect 145104 995444 145156 995450
rect 145104 995386 145156 995392
rect 145012 993812 145064 993818
rect 145012 993754 145064 993760
rect 151820 993744 151872 993750
rect 151820 993686 151872 993692
rect 151832 989466 151860 993686
rect 151820 989460 151872 989466
rect 151820 989402 151872 989408
rect 138296 988780 138348 988786
rect 138296 988722 138348 988728
rect 144828 988780 144880 988786
rect 144828 988722 144880 988728
rect 125508 986944 125560 986950
rect 125508 986886 125560 986892
rect 138308 983620 138336 988722
rect 154500 983620 154528 1004634
rect 155776 999592 155828 999598
rect 155774 999560 155776 999569
rect 160284 999592 160336 999598
rect 155828 999560 155830 999569
rect 155774 999495 155830 999504
rect 159086 999560 159142 999569
rect 160284 999534 160336 999540
rect 159086 999495 159088 999504
rect 159140 999495 159142 999504
rect 159088 999466 159140 999472
rect 155776 999184 155828 999190
rect 155774 999152 155776 999161
rect 155828 999152 155830 999161
rect 155774 999087 155830 999096
rect 158258 999152 158314 999161
rect 158258 999087 158260 999096
rect 158312 999087 158314 999096
rect 158260 999058 158312 999064
rect 156142 997792 156198 997801
rect 156142 997727 156144 997736
rect 156196 997727 156198 997736
rect 156144 997698 156196 997704
rect 157800 996187 157852 996193
rect 156970 996155 157026 996164
rect 156970 996090 157026 996099
rect 157798 996155 157800 996164
rect 157852 996155 157854 996164
rect 157798 996090 157854 996099
rect 159454 996155 159510 996164
rect 159454 996090 159456 996099
rect 156984 996057 157012 996090
rect 159508 996090 159510 996099
rect 159456 996061 159508 996067
rect 156972 996051 157024 996057
rect 156972 995993 157024 995999
rect 160296 993682 160324 999534
rect 162860 999524 162912 999530
rect 162860 999466 162912 999472
rect 162872 997264 162900 999466
rect 162872 997236 168900 997264
rect 162872 997235 162900 997236
rect 168872 997121 168900 997236
rect 168858 997112 168914 997121
rect 168858 997047 168914 997056
rect 173912 996193 173940 1004906
rect 174084 1004828 174136 1004834
rect 174084 1004770 174136 1004776
rect 173992 1004760 174044 1004766
rect 173992 1004702 174044 1004708
rect 173900 996187 173952 996193
rect 173900 996129 173952 996135
rect 174004 996125 174032 1004702
rect 173992 996119 174044 996125
rect 173992 996061 174044 996067
rect 174096 996057 174124 1004770
rect 160468 996051 160520 996057
rect 160468 995993 160520 995999
rect 174084 996051 174136 996057
rect 174084 995993 174136 995999
rect 160284 993676 160336 993682
rect 160284 993618 160336 993624
rect 160480 984162 160508 995993
rect 162950 995752 163006 995761
rect 162950 995687 163006 995696
rect 162858 995616 162914 995625
rect 162858 995551 162914 995560
rect 162872 984298 162900 995551
rect 162860 984292 162912 984298
rect 162860 984234 162912 984240
rect 162964 984230 162992 995687
rect 168378 993728 168434 993737
rect 168378 993663 168434 993672
rect 168392 990690 168420 993663
rect 168380 990684 168432 990690
rect 168380 990626 168432 990632
rect 170404 990684 170456 990690
rect 170404 990626 170456 990632
rect 162952 984224 163004 984230
rect 162952 984166 163004 984172
rect 160468 984156 160520 984162
rect 160468 984098 160520 984104
rect 170416 983634 170444 990626
rect 175200 987018 175228 1005042
rect 195152 1004692 195204 1004698
rect 195152 1004634 195204 1004640
rect 195164 997257 195192 1004634
rect 195244 999388 195296 999394
rect 195244 999330 195296 999336
rect 195150 997248 195206 997257
rect 195150 997183 195206 997192
rect 195256 995853 195284 999330
rect 195348 997121 195376 1005450
rect 195704 1004828 195756 1004834
rect 195704 1004770 195756 1004776
rect 195428 999728 195480 999734
rect 195428 999670 195480 999676
rect 195334 997112 195390 997121
rect 195334 997047 195390 997056
rect 188804 995838 188856 995844
rect 183284 995784 183336 995790
rect 182988 995732 183284 995738
rect 188804 995780 188856 995786
rect 189448 995842 189500 995848
rect 195244 995847 195296 995853
rect 189448 995784 189500 995790
rect 194324 995784 194376 995790
rect 195244 995789 195296 995795
rect 195440 995790 195468 999670
rect 195520 999660 195572 999666
rect 195520 999602 195572 999608
rect 187606 995752 187662 995761
rect 182988 995726 183336 995732
rect 182988 995710 183324 995726
rect 187312 995710 187606 995738
rect 188816 995738 188844 995780
rect 189460 995738 189488 995784
rect 187864 995722 188200 995738
rect 187864 995716 188212 995722
rect 187864 995710 188160 995716
rect 187606 995687 187662 995696
rect 188508 995710 188844 995738
rect 189152 995710 189488 995738
rect 194028 995732 194324 995738
rect 194028 995726 194376 995732
rect 195428 995784 195480 995790
rect 195428 995726 195480 995732
rect 194028 995710 194364 995726
rect 188160 995658 188212 995664
rect 184664 995648 184716 995654
rect 192482 995616 192538 995625
rect 184716 995596 184828 995602
rect 184664 995590 184828 995596
rect 184676 995574 184828 995590
rect 190348 995586 190684 995602
rect 190348 995580 190696 995586
rect 190348 995574 190644 995580
rect 192188 995574 192482 995602
rect 195532 995586 195560 999602
rect 195612 999592 195664 999598
rect 195612 999534 195664 999540
rect 195624 995921 195652 999534
rect 195716 995989 195744 1004770
rect 198464 999524 198516 999530
rect 198464 999466 198516 999472
rect 198372 999456 198424 999462
rect 198372 999398 198424 999404
rect 195704 995983 195756 995989
rect 195704 995925 195756 995931
rect 195612 995915 195664 995921
rect 195612 995857 195664 995863
rect 192482 995551 192538 995560
rect 195520 995580 195572 995586
rect 190644 995522 190696 995528
rect 195520 995522 195572 995528
rect 184480 995512 184532 995518
rect 179860 995438 180196 995466
rect 180504 995438 180840 995466
rect 181148 995438 181484 995466
rect 183540 995450 183876 995466
rect 184184 995460 184480 995466
rect 184184 995454 184532 995460
rect 183540 995444 183888 995450
rect 183540 995438 183836 995444
rect 180168 993818 180196 995438
rect 180156 993812 180208 993818
rect 180156 993754 180208 993760
rect 180812 993750 180840 995438
rect 180800 993744 180852 993750
rect 180800 993686 180852 993692
rect 181456 993682 181484 995438
rect 184184 995438 184520 995454
rect 191544 995438 191880 995466
rect 198384 995450 198412 999398
rect 198476 995518 198504 999466
rect 198648 999252 198700 999258
rect 198648 999194 198700 999200
rect 198556 999184 198608 999190
rect 198556 999126 198608 999132
rect 198568 995654 198596 999126
rect 198660 995722 198688 999194
rect 198648 995716 198700 995722
rect 198648 995658 198700 995664
rect 198556 995648 198608 995654
rect 198556 995590 198608 995596
rect 198464 995512 198516 995518
rect 198464 995454 198516 995460
rect 183836 995386 183888 995392
rect 191852 993721 191880 995438
rect 198372 995444 198424 995450
rect 198372 995386 198424 995392
rect 200040 993818 200068 1005518
rect 207202 1005479 207258 1005488
rect 209594 1005544 209650 1005553
rect 209594 1005479 209596 1005488
rect 209648 1005479 209650 1005488
rect 361026 1005544 361082 1005553
rect 361026 1005479 361028 1005488
rect 209596 1005450 209648 1005456
rect 263852 1005464 263908 1005473
rect 361080 1005479 361082 1005488
rect 361028 1005450 361080 1005456
rect 263908 1005422 266868 1005450
rect 263852 1005399 263908 1005408
rect 264933 1005351 265433 1005379
rect 259828 1005304 259880 1005310
rect 259826 1005272 259828 1005281
rect 259880 1005272 259882 1005281
rect 259826 1005207 259882 1005216
rect 260194 1005272 260250 1005281
rect 260194 1005207 260196 1005216
rect 260248 1005207 260250 1005216
rect 260196 1005178 260248 1005184
rect 201868 1005168 201920 1005174
rect 227628 1005168 227680 1005174
rect 201868 1005110 201920 1005116
rect 208398 1005136 208454 1005145
rect 201880 1004766 201908 1005110
rect 261852 1005168 261904 1005174
rect 227628 1005110 227680 1005116
rect 261850 1005136 261852 1005145
rect 261904 1005136 261906 1005145
rect 208398 1005071 208400 1005080
rect 208452 1005071 208454 1005080
rect 208400 1005042 208452 1005048
rect 211620 1005032 211672 1005038
rect 209226 1005000 209282 1005009
rect 204168 1004964 204220 1004970
rect 209226 1004935 209228 1004944
rect 204168 1004906 204220 1004912
rect 209280 1004935 209282 1004944
rect 211618 1005000 211620 1005009
rect 211672 1005000 211674 1005009
rect 211618 1004935 211674 1004944
rect 209228 1004906 209280 1004912
rect 201040 1004760 201092 1004766
rect 201038 1004728 201040 1004737
rect 201868 1004760 201920 1004766
rect 201092 1004728 201094 1004737
rect 201038 1004663 201094 1004672
rect 201866 1004728 201868 1004737
rect 201920 1004728 201922 1004737
rect 201866 1004663 201922 1004672
rect 203890 999696 203946 999705
rect 203890 999631 203892 999640
rect 203944 999631 203946 999640
rect 203892 999602 203944 999608
rect 203524 999592 203576 999598
rect 203522 999560 203524 999569
rect 203576 999560 203578 999569
rect 203522 999495 203578 999504
rect 202234 999424 202290 999433
rect 202234 999359 202236 999368
rect 202288 999359 202290 999368
rect 202236 999330 202288 999336
rect 200120 999320 200172 999326
rect 200120 999262 200172 999268
rect 202694 999288 202750 999297
rect 200028 993812 200080 993818
rect 200028 993754 200080 993760
rect 200132 993750 200160 999262
rect 202694 999223 202696 999232
rect 202748 999223 202750 999232
rect 202696 999194 202748 999200
rect 203064 999184 203116 999190
rect 203062 999152 203064 999161
rect 203116 999152 203118 999161
rect 203062 999087 203118 999096
rect 200120 993744 200172 993750
rect 191838 993712 191894 993721
rect 181444 993676 181496 993682
rect 200120 993686 200172 993692
rect 191838 993647 191894 993656
rect 181444 993618 181496 993624
rect 204180 990690 204208 1004906
rect 210884 1004896 210936 1004902
rect 206374 1004864 206430 1004873
rect 206374 1004799 206376 1004808
rect 206428 1004799 206430 1004808
rect 210882 1004864 210884 1004873
rect 210936 1004864 210938 1004873
rect 210882 1004799 210938 1004808
rect 206376 1004770 206428 1004776
rect 205914 1004728 205970 1004737
rect 205914 1004663 205916 1004672
rect 205968 1004663 205970 1004672
rect 212458 1004728 212514 1004737
rect 212458 1004663 212514 1004672
rect 205916 1004634 205968 1004640
rect 212472 1004607 212500 1004663
rect 212472 1004579 218100 1004607
rect 218072 999734 218100 1004579
rect 205548 999728 205600 999734
rect 205546 999696 205548 999705
rect 218072 999706 219112 999734
rect 205600 999696 205602 999705
rect 205546 999631 205602 999640
rect 204350 999560 204406 999569
rect 204350 999495 204352 999504
rect 204404 999495 204406 999504
rect 204352 999466 204404 999472
rect 204720 999456 204772 999462
rect 204718 999424 204720 999433
rect 208860 999456 208912 999462
rect 204772 999424 204774 999433
rect 204718 999359 204774 999368
rect 208858 999424 208860 999433
rect 212724 999456 212776 999462
rect 208912 999424 208914 999433
rect 208858 999359 208914 999368
rect 210422 999424 210478 999433
rect 212724 999398 212776 999404
rect 210422 999359 210424 999368
rect 210476 999359 210478 999368
rect 210424 999330 210476 999336
rect 205180 999320 205232 999326
rect 205178 999288 205180 999297
rect 209596 999320 209648 999326
rect 205232 999288 205234 999297
rect 205178 999223 205234 999232
rect 209594 999288 209596 999297
rect 212632 999320 212684 999326
rect 209648 999288 209650 999297
rect 209594 999223 209650 999232
rect 211710 999288 211766 999297
rect 212632 999262 212684 999268
rect 211710 999223 211712 999232
rect 211764 999223 211766 999232
rect 211712 999194 211764 999200
rect 211252 999184 211304 999190
rect 207570 999152 207626 999161
rect 207570 999087 207626 999096
rect 211250 999152 211252 999161
rect 211304 999152 211306 999161
rect 211250 999087 211306 999096
rect 207584 993682 207612 999087
rect 212644 996125 212672 999262
rect 212632 996119 212684 996125
rect 212632 996061 212684 996067
rect 207572 993676 207624 993682
rect 207572 993618 207624 993624
rect 203156 990684 203208 990690
rect 203156 990626 203208 990632
rect 204168 990684 204220 990690
rect 204168 990626 204220 990632
rect 186964 989460 187016 989466
rect 186964 989402 187016 989408
rect 175188 987012 175240 987018
rect 175188 986954 175240 986960
rect 170416 983606 170798 983634
rect 186976 983620 187004 989402
rect 203168 983620 203196 990626
rect 212644 987222 212672 996061
rect 212736 996057 212764 999398
rect 218972 999388 219024 999394
rect 218972 999330 219024 999336
rect 216588 999252 216640 999258
rect 216588 999194 216640 999200
rect 215300 999184 215352 999190
rect 215300 999126 215352 999132
rect 215312 996193 215340 999126
rect 215300 996187 215352 996193
rect 215300 996129 215352 996135
rect 212724 996051 212776 996057
rect 212724 995993 212776 995999
rect 212632 987216 212684 987222
rect 212632 987158 212684 987164
rect 212736 987086 212764 995993
rect 215312 987154 215340 996129
rect 216600 989466 216628 999194
rect 218984 997257 219012 999330
rect 218970 997248 219026 997257
rect 218970 997183 219026 997192
rect 216588 989460 216640 989466
rect 216588 989402 216640 989408
rect 215300 987148 215352 987154
rect 215300 987090 215352 987096
rect 212724 987080 212776 987086
rect 212724 987022 212776 987028
rect 219084 983634 219112 999706
rect 227640 987290 227668 1005110
rect 227812 1005100 227864 1005106
rect 261850 1005071 261906 1005080
rect 263046 1005136 263102 1005145
rect 263046 1005071 263048 1005080
rect 227812 1005042 227864 1005048
rect 263100 1005071 263102 1005080
rect 263048 1005042 263100 1005048
rect 227720 1004964 227772 1004970
rect 227720 1004906 227772 1004912
rect 227732 996057 227760 1004906
rect 227824 996125 227852 1005042
rect 260656 1005032 260708 1005038
rect 260654 1005000 260656 1005009
rect 260708 1005000 260710 1005009
rect 260654 1004935 260710 1004944
rect 262678 1005000 262734 1005009
rect 262678 1004935 262680 1004944
rect 262732 1004935 262734 1004944
rect 262680 1004906 262732 1004912
rect 261024 1004896 261076 1004902
rect 261022 1004864 261024 1004873
rect 261076 1004864 261078 1004873
rect 227904 1004828 227956 1004834
rect 261022 1004799 261078 1004808
rect 262218 1004864 262274 1004873
rect 262218 1004799 262220 1004808
rect 227904 1004770 227956 1004776
rect 262272 1004799 262274 1004808
rect 262220 1004770 262272 1004776
rect 227916 996193 227944 1004770
rect 261484 1004760 261536 1004766
rect 252466 1004728 252522 1004737
rect 252466 1004663 252468 1004672
rect 252520 1004663 252522 1004672
rect 253294 1004728 253350 1004737
rect 253294 1004663 253296 1004672
rect 252468 1004634 252520 1004640
rect 253348 1004663 253350 1004672
rect 261482 1004728 261484 1004737
rect 261536 1004728 261538 1004737
rect 261482 1004663 261538 1004672
rect 263506 1004728 263562 1004737
rect 264933 1004714 264961 1005351
rect 265256 1005236 265308 1005242
rect 265256 1005178 265308 1005184
rect 265072 1004896 265124 1004902
rect 265072 1004838 265124 1004844
rect 263562 1004686 264961 1004714
rect 263506 1004663 263562 1004672
rect 253296 1004634 253348 1004640
rect 258630 999968 258686 999977
rect 246764 999932 246816 999938
rect 258630 999903 258632 999912
rect 246764 999874 246816 999880
rect 258684 999903 258686 999912
rect 258632 999874 258684 999880
rect 246672 999864 246724 999870
rect 246672 999806 246724 999812
rect 246580 999796 246632 999802
rect 246580 999738 246632 999744
rect 246592 999682 246620 999738
rect 246500 999654 246620 999682
rect 227904 996187 227956 996193
rect 227904 996129 227956 996135
rect 227812 996119 227864 996125
rect 227812 996061 227864 996067
rect 227720 996051 227772 996057
rect 227720 995993 227772 995999
rect 246500 995858 246528 999654
rect 240876 995852 240928 995858
rect 240876 995794 240928 995800
rect 245568 995852 245620 995858
rect 245568 995794 245620 995800
rect 246488 995852 246540 995858
rect 246488 995794 246540 995800
rect 239036 995784 239088 995790
rect 235262 995752 235318 995761
rect 234968 995710 235262 995738
rect 235906 995752 235962 995761
rect 235612 995710 235906 995738
rect 235262 995687 235318 995696
rect 238740 995732 239036 995738
rect 240888 995738 240916 995794
rect 242070 995752 242126 995761
rect 238740 995726 239088 995732
rect 238740 995710 239076 995726
rect 240580 995710 240916 995738
rect 241776 995710 242070 995738
rect 235906 995687 235962 995696
rect 245580 995738 245608 995794
rect 246684 995790 246712 999806
rect 243616 995722 243952 995738
rect 243616 995716 243964 995722
rect 243616 995710 243912 995716
rect 242070 995687 242126 995696
rect 245456 995710 245608 995738
rect 246672 995784 246724 995790
rect 246672 995726 246724 995732
rect 246776 995722 246804 999874
rect 257344 999864 257396 999870
rect 256974 999832 257030 999841
rect 256974 999767 256976 999776
rect 257028 999767 257030 999776
rect 257342 999832 257344 999841
rect 257396 999832 257398 999841
rect 257342 999767 257398 999776
rect 256976 999738 257028 999744
rect 246856 999728 246908 999734
rect 257804 999728 257856 999734
rect 246856 999670 246908 999676
rect 254858 999696 254914 999705
rect 246764 995716 246816 995722
rect 243912 995658 243964 995664
rect 246764 995658 246816 995664
rect 239588 995648 239640 995654
rect 239292 995596 239588 995602
rect 240046 995616 240102 995625
rect 239292 995590 239640 995596
rect 239292 995574 239628 995590
rect 239936 995574 240046 995602
rect 240046 995551 240102 995560
rect 236550 995480 236606 995489
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 231596 993682 231624 995438
rect 232240 994129 232268 995438
rect 232226 994120 232282 994129
rect 232226 994055 232282 994064
rect 232884 993993 232912 995438
rect 234402 995353 234430 995452
rect 236256 995438 236550 995466
rect 242972 995438 243308 995466
rect 236550 995415 236606 995424
rect 234388 995344 234444 995353
rect 234388 995279 234444 995288
rect 232870 993984 232926 993993
rect 232870 993919 232926 993928
rect 243280 993857 243308 995438
rect 246868 995353 246896 999670
rect 249708 999660 249760 999666
rect 254858 999631 254860 999640
rect 249708 999602 249760 999608
rect 254912 999631 254914 999640
rect 257802 999696 257804 999705
rect 257856 999696 257858 999705
rect 257802 999631 257858 999640
rect 254860 999602 254912 999608
rect 246948 999388 247000 999394
rect 246948 999330 247000 999336
rect 246960 995926 246988 999330
rect 247960 999116 248012 999122
rect 247960 999058 248012 999064
rect 247972 997257 248000 999058
rect 247958 997248 248014 997257
rect 247958 997183 248014 997192
rect 246948 995920 247000 995926
rect 246948 995862 247000 995868
rect 249720 995625 249748 999602
rect 250444 999592 250496 999598
rect 256148 999592 256200 999598
rect 250444 999534 250496 999540
rect 255686 999560 255742 999569
rect 250260 999524 250312 999530
rect 250260 999466 250312 999472
rect 250076 999456 250128 999462
rect 250076 999398 250128 999404
rect 249892 999320 249944 999326
rect 249892 999262 249944 999268
rect 249706 995616 249762 995625
rect 249706 995551 249762 995560
rect 249904 995489 249932 999262
rect 250088 995761 250116 999398
rect 250272 995897 250300 999466
rect 250456 996033 250484 999534
rect 255686 999495 255688 999504
rect 255740 999495 255742 999504
rect 256146 999560 256148 999569
rect 256200 999560 256202 999569
rect 256146 999495 256202 999504
rect 255688 999466 255740 999472
rect 255320 999456 255372 999462
rect 253662 999424 253718 999433
rect 253662 999359 253664 999368
rect 253716 999359 253718 999368
rect 255318 999424 255320 999433
rect 255372 999424 255374 999433
rect 255318 999359 255374 999368
rect 253664 999330 253716 999336
rect 254492 999320 254544 999326
rect 254490 999288 254492 999297
rect 254544 999288 254546 999297
rect 252468 999252 252520 999258
rect 254490 999223 254546 999232
rect 256514 999288 256570 999297
rect 256514 999223 256516 999232
rect 252468 999194 252520 999200
rect 256568 999223 256570 999232
rect 256516 999194 256568 999200
rect 250628 999184 250680 999190
rect 250628 999126 250680 999132
rect 250442 996024 250498 996033
rect 250442 995959 250498 995968
rect 250258 995888 250314 995897
rect 250258 995823 250314 995832
rect 250074 995752 250130 995761
rect 250074 995687 250130 995696
rect 250640 995654 250668 999126
rect 250628 995648 250680 995654
rect 250628 995590 250680 995596
rect 249890 995480 249946 995489
rect 249890 995415 249946 995424
rect 246854 995344 246910 995353
rect 246854 995279 246910 995288
rect 252480 994129 252508 999194
rect 254124 999184 254176 999190
rect 254122 999152 254124 999161
rect 258540 999184 258592 999190
rect 254176 999152 254178 999161
rect 254122 999087 254178 999096
rect 258538 999152 258540 999161
rect 262220 999184 262272 999190
rect 258592 999152 258594 999161
rect 262220 999126 262272 999132
rect 258538 999087 258594 999096
rect 252466 994120 252522 994129
rect 252466 994055 252522 994064
rect 243266 993848 243322 993857
rect 243266 993783 243322 993792
rect 248326 993712 248382 993721
rect 231584 993676 231636 993682
rect 262232 993682 262260 999126
rect 265084 996057 265112 1004838
rect 265164 1004760 265216 1004766
rect 265164 1004686 265216 1004708
rect 265176 999122 265204 1004686
rect 265164 999116 265216 999122
rect 265164 999058 265216 999064
rect 265268 996125 265296 1005178
rect 265405 1004714 265433 1005351
rect 265534 1005136 265590 1005145
rect 265534 1005071 265536 1005080
rect 265588 1005071 265590 1005080
rect 265536 1005042 265588 1005048
rect 265534 1005000 265590 1005009
rect 265534 1004935 265536 1004944
rect 265588 1004935 265590 1004944
rect 266630 1005000 266686 1005009
rect 266630 1004935 266686 1004944
rect 265536 1004906 265588 1004912
rect 265474 1004728 265530 1004737
rect 265405 1004686 265474 1004714
rect 265474 1004663 265530 1004672
rect 266538 1004728 266594 1004737
rect 266538 1004663 266594 1004672
rect 266552 1003045 266580 1004663
rect 266644 1003165 266672 1004935
rect 266840 1003317 266868 1005422
rect 360198 1005408 360254 1005417
rect 360198 1005343 360200 1005352
rect 360252 1005343 360254 1005352
rect 360200 1005314 360252 1005320
rect 280344 1005304 280396 1005310
rect 280344 1005246 280396 1005252
rect 359738 1005272 359794 1005281
rect 267010 1005136 267066 1005145
rect 267010 1005071 267066 1005080
rect 270468 1005100 270520 1005106
rect 267024 1003451 267052 1005071
rect 270468 1005042 270520 1005048
rect 267024 1003423 269252 1003451
rect 267024 1003418 267052 1003423
rect 266840 1003289 269068 1003317
rect 266644 1003137 267871 1003165
rect 266552 1003017 267780 1003045
rect 265256 996119 265308 996125
rect 265256 996061 265308 996067
rect 267648 996119 267700 996125
rect 267648 996061 267700 996067
rect 265072 996051 265124 996057
rect 265072 995993 265124 995999
rect 267556 996051 267608 996057
rect 267556 995993 267608 995999
rect 248326 993647 248382 993656
rect 262220 993676 262272 993682
rect 231584 993618 231636 993624
rect 235632 989460 235684 989466
rect 235632 989402 235684 989408
rect 227628 987284 227680 987290
rect 227628 987226 227680 987232
rect 219084 983606 219466 983634
rect 235644 983620 235672 989402
rect 248340 988174 248368 993647
rect 262220 993618 262272 993624
rect 248328 988168 248380 988174
rect 248328 988110 248380 988116
rect 251824 988168 251876 988174
rect 251824 988110 251876 988116
rect 251836 983620 251864 988110
rect 267568 987358 267596 995993
rect 267660 987494 267688 996061
rect 267648 987488 267700 987494
rect 267648 987430 267700 987436
rect 267556 987352 267608 987358
rect 267556 987294 267608 987300
rect 267752 983634 267780 1003017
rect 267843 1003031 267871 1003137
rect 267843 1002996 267872 1003031
rect 267844 996193 267872 1002996
rect 267832 996187 267884 996193
rect 267832 996129 267884 996135
rect 269040 989466 269068 1003289
rect 269224 989534 269252 1003423
rect 270480 997257 270508 1005042
rect 280160 1004964 280212 1004970
rect 280160 1004906 280212 1004912
rect 280068 1004692 280120 1004698
rect 280068 1004634 280120 1004640
rect 270466 997248 270522 997257
rect 270466 997183 270522 997192
rect 270408 996187 270460 996193
rect 270408 996129 270460 996135
rect 269212 989528 269264 989534
rect 269212 989470 269264 989476
rect 269028 989460 269080 989466
rect 269028 989402 269080 989408
rect 270420 987562 270448 996129
rect 280080 987630 280108 1004634
rect 280172 996120 280200 1004906
rect 280252 1004828 280304 1004834
rect 280252 1004770 280304 1004776
rect 280264 996188 280292 1004770
rect 280252 996182 280304 996188
rect 280252 996124 280304 996130
rect 280160 996114 280212 996120
rect 280160 996056 280212 996062
rect 280356 996052 280384 1005246
rect 359738 1005207 359740 1005216
rect 359792 1005207 359794 1005216
rect 370412 1005236 370464 1005242
rect 359740 1005178 359792 1005184
rect 370412 1005178 370464 1005184
rect 358174 1005136 358230 1005145
rect 358174 1005071 358176 1005080
rect 358228 1005071 358230 1005080
rect 366732 1005100 366784 1005106
rect 358176 1005042 358228 1005048
rect 366732 1005042 366784 1005048
rect 356888 1005032 356940 1005038
rect 356886 1005000 356888 1005009
rect 356940 1005000 356942 1005009
rect 356886 1004935 356942 1004944
rect 358542 1005000 358598 1005009
rect 358542 1004935 358544 1004944
rect 358596 1004935 358598 1004944
rect 358544 1004906 358596 1004912
rect 357348 1004896 357400 1004902
rect 357346 1004864 357348 1004873
rect 362500 1004896 362552 1004902
rect 357400 1004864 357402 1004873
rect 357346 1004799 357402 1004808
rect 357714 1004864 357770 1004873
rect 362500 1004838 362552 1004844
rect 357714 1004799 357716 1004808
rect 357768 1004799 357770 1004808
rect 357716 1004770 357768 1004776
rect 360568 1004760 360620 1004766
rect 315118 1004728 315174 1004737
rect 350446 1004728 350502 1004737
rect 315118 1004663 315120 1004672
rect 315172 1004663 315174 1004672
rect 331220 1004692 331272 1004698
rect 315120 1004634 315172 1004640
rect 350446 1004663 350502 1004672
rect 353666 1004728 353722 1004737
rect 354034 1004728 354090 1004737
rect 353722 1004686 354034 1004714
rect 353666 1004663 353722 1004672
rect 354034 1004663 354090 1004672
rect 354494 1004728 354550 1004737
rect 355230 1004728 355286 1004737
rect 354550 1004686 355230 1004714
rect 354494 1004663 354550 1004672
rect 355230 1004663 355286 1004672
rect 360566 1004728 360568 1004737
rect 360620 1004728 360622 1004737
rect 360566 1004663 360622 1004672
rect 361394 1004728 361450 1004737
rect 361394 1004663 361396 1004672
rect 331220 1004634 331272 1004640
rect 312176 999864 312228 999870
rect 310150 999832 310206 999841
rect 310150 999767 310152 999776
rect 310204 999767 310206 999776
rect 312174 999832 312176 999841
rect 318892 999864 318944 999870
rect 312228 999832 312230 999841
rect 318892 999806 318944 999812
rect 312174 999767 312230 999776
rect 314936 999796 314988 999802
rect 310152 999738 310204 999744
rect 314936 999738 314988 999744
rect 311440 999728 311492 999734
rect 311438 999696 311440 999705
rect 311492 999696 311494 999705
rect 311438 999631 311494 999640
rect 313830 999696 313886 999705
rect 313830 999631 313832 999640
rect 313884 999631 313886 999640
rect 313832 999602 313884 999608
rect 312636 999592 312688 999598
rect 312634 999560 312636 999569
rect 312688 999560 312690 999569
rect 312634 999495 312690 999504
rect 314658 999560 314714 999569
rect 314714 999530 314884 999546
rect 314714 999524 314896 999530
rect 314714 999518 314844 999524
rect 314658 999495 314714 999504
rect 314844 999466 314896 999472
rect 312634 999152 312690 999161
rect 298744 999116 298796 999122
rect 312634 999087 312636 999096
rect 298744 999058 298796 999064
rect 312688 999087 312690 999096
rect 312636 999058 312688 999064
rect 298756 997257 298784 999058
rect 298742 997248 298798 997257
rect 298742 997183 298798 997192
rect 301780 996328 301832 996334
rect 308128 996328 308180 996334
rect 301780 996270 301832 996276
rect 305734 996296 305790 996305
rect 300216 996260 300268 996266
rect 300216 996202 300268 996208
rect 280344 996046 280396 996052
rect 280344 995988 280396 995994
rect 286784 995852 286836 995858
rect 286784 995794 286836 995800
rect 293592 995842 293644 995848
rect 286796 995738 286824 995794
rect 293592 995784 293644 995790
rect 295064 995842 295116 995848
rect 295064 995784 295116 995790
rect 288070 995752 288126 995761
rect 286534 995710 286824 995738
rect 287822 995710 288070 995738
rect 292486 995752 292542 995761
rect 291502 995722 291792 995738
rect 291502 995716 291804 995722
rect 291502 995710 291752 995716
rect 288070 995687 288126 995696
rect 292146 995710 292486 995738
rect 293604 995738 293632 995784
rect 293342 995710 293632 995738
rect 295076 995738 295104 995784
rect 295076 995710 295182 995738
rect 292486 995687 292542 995696
rect 291752 995658 291804 995664
rect 287520 995648 287572 995654
rect 287178 995596 287520 995602
rect 300228 995625 300256 996202
rect 300766 995888 300822 995897
rect 300766 995823 300822 995832
rect 291106 995616 291162 995625
rect 287178 995590 287572 995596
rect 287178 995574 287560 995590
rect 290858 995574 291106 995602
rect 291106 995551 291162 995560
rect 300214 995616 300270 995625
rect 300214 995551 300270 995560
rect 290554 995480 290610 995489
rect 282840 993750 282868 995452
rect 283484 993886 283512 995452
rect 283472 993880 283524 993886
rect 283472 993822 283524 993828
rect 282828 993744 282880 993750
rect 282828 993686 282880 993692
rect 284128 993682 284156 995452
rect 285968 993818 285996 995452
rect 290306 995438 290554 995466
rect 297270 995480 297326 995489
rect 290554 995415 290610 995424
rect 285956 993812 286008 993818
rect 285956 993754 286008 993760
rect 294524 993721 294552 995452
rect 297022 995438 297270 995466
rect 297270 995415 297326 995424
rect 294510 993712 294566 993721
rect 284116 993676 284168 993682
rect 294510 993647 294566 993656
rect 284116 993618 284168 993624
rect 300492 989528 300544 989534
rect 300492 989470 300544 989476
rect 284300 989460 284352 989466
rect 284300 989402 284352 989408
rect 280068 987624 280120 987630
rect 280068 987566 280120 987572
rect 270408 987556 270460 987562
rect 270408 987498 270460 987504
rect 267752 983606 268134 983634
rect 284312 983620 284340 989402
rect 300504 983620 300532 989470
rect 300780 984706 300808 995823
rect 301792 993886 301820 996270
rect 305734 996231 305736 996240
rect 305788 996231 305790 996240
rect 308126 996296 308128 996305
rect 308180 996296 308182 996305
rect 308126 996231 308182 996240
rect 305736 996202 305788 996208
rect 314304 996198 314332 996229
rect 314292 996192 314344 996198
rect 305274 996160 305330 996169
rect 305274 996095 305330 996104
rect 306470 996160 306526 996169
rect 306470 996095 306526 996104
rect 306930 996160 306986 996169
rect 306930 996095 306986 996104
rect 307298 996160 307354 996169
rect 307298 996095 307354 996104
rect 307758 996160 307814 996169
rect 307758 996095 307814 996104
rect 309322 996160 309378 996169
rect 309322 996095 309378 996104
rect 310150 996160 310206 996169
rect 310150 996095 310206 996104
rect 310610 996160 310666 996169
rect 310610 996095 310666 996104
rect 311806 996160 311862 996169
rect 311806 996095 311862 996104
rect 314290 996160 314292 996169
rect 314344 996160 314346 996169
rect 314290 996095 314346 996104
rect 305288 995625 305316 996095
rect 306484 995722 306512 996095
rect 306944 995916 306972 996095
rect 306932 995910 306984 995916
rect 306932 995852 306984 995858
rect 306472 995716 306524 995722
rect 306472 995658 306524 995664
rect 307312 995654 307340 996095
rect 307772 995984 307800 996095
rect 307760 995978 307812 995984
rect 307760 995920 307812 995926
rect 307300 995648 307352 995654
rect 305274 995616 305330 995625
rect 307300 995590 307352 995596
rect 305274 995551 305330 995560
rect 303528 994772 303580 994778
rect 303528 994714 303580 994720
rect 301780 993880 301832 993886
rect 301780 993822 301832 993828
rect 303540 989466 303568 994714
rect 309336 993818 309364 996095
rect 310164 995858 310192 996095
rect 310152 995852 310204 995858
rect 310152 995794 310204 995800
rect 309324 993812 309376 993818
rect 309324 993754 309376 993760
rect 310624 993682 310652 996095
rect 311820 996052 311848 996095
rect 311808 996046 311860 996052
rect 311808 995988 311860 995994
rect 310612 993676 310664 993682
rect 310612 993618 310664 993624
rect 303528 989460 303580 989466
rect 303528 989402 303580 989408
rect 311820 987766 311848 995988
rect 314304 987902 314332 996095
rect 314948 993750 314976 999738
rect 315948 999728 316000 999734
rect 315948 999670 316000 999676
rect 315120 999592 315172 999598
rect 315120 999534 315172 999540
rect 315132 996130 315160 999534
rect 315120 996124 315172 996130
rect 315120 996066 315172 996072
rect 314936 993744 314988 993750
rect 314936 993686 314988 993692
rect 314292 987896 314344 987902
rect 314292 987838 314344 987844
rect 311808 987760 311860 987766
rect 311808 987702 311860 987708
rect 315960 984774 315988 999670
rect 318708 999660 318760 999666
rect 318708 999602 318760 999608
rect 317512 996124 317564 996130
rect 317512 996066 317564 996072
rect 316774 993848 316830 993857
rect 316774 993783 316830 993792
rect 315948 984768 316000 984774
rect 315948 984710 316000 984716
rect 300768 984700 300820 984706
rect 300768 984642 300820 984648
rect 316788 983620 316816 993783
rect 317524 984842 317552 996066
rect 318720 987698 318748 999602
rect 318904 987834 318932 999806
rect 319076 999524 319128 999530
rect 319076 999466 319128 999472
rect 319088 989534 319116 999466
rect 321466 993580 321522 993589
rect 321466 993515 321522 993524
rect 321480 989602 321508 993515
rect 331232 990690 331260 1004634
rect 331220 990684 331272 990690
rect 331220 990626 331272 990632
rect 332692 990684 332744 990690
rect 332692 990626 332744 990632
rect 321468 989596 321520 989602
rect 321468 989538 321520 989544
rect 319076 989528 319128 989534
rect 319076 989470 319128 989476
rect 318892 987828 318944 987834
rect 318892 987770 318944 987776
rect 318708 987692 318760 987698
rect 318708 987634 318760 987640
rect 317512 984836 317564 984842
rect 317512 984778 317564 984784
rect 332704 983634 332732 990626
rect 349160 989596 349212 989602
rect 349160 989538 349212 989544
rect 332704 983606 332994 983634
rect 349172 983620 349200 989538
rect 350460 985114 350488 1004663
rect 361448 1004663 361450 1004672
rect 361396 1004634 361448 1004640
rect 362512 1001910 362540 1004838
rect 364248 1004828 364300 1004834
rect 364248 1004770 364300 1004776
rect 362500 1001904 362552 1001910
rect 362500 1001846 362552 1001852
rect 364260 1001858 364288 1004770
rect 366364 1004760 366416 1004766
rect 366364 1004702 366416 1004708
rect 365444 1004692 365496 1004698
rect 365444 1004634 365496 1004640
rect 364432 1001904 364484 1001910
rect 364260 1001830 364380 1001858
rect 364432 1001846 364484 1001852
rect 358912 1000544 358964 1000550
rect 358910 1000512 358912 1000521
rect 358964 1000512 358966 1000521
rect 358910 1000447 358966 1000456
rect 361856 999728 361908 999734
rect 361854 999696 361856 999705
rect 361908 999696 361910 999705
rect 361854 999631 361910 999640
rect 362590 999696 362646 999705
rect 362590 999631 362592 999640
rect 362644 999631 362646 999640
rect 362592 999602 362644 999608
rect 363420 999592 363472 999598
rect 363418 999560 363420 999569
rect 363472 999560 363474 999569
rect 363418 999495 363474 999504
rect 362224 999456 362276 999462
rect 362222 999424 362224 999433
rect 362276 999424 362278 999433
rect 362222 999359 362278 999368
rect 364246 999288 364302 999297
rect 364246 999223 364248 999232
rect 364300 999223 364302 999232
rect 364248 999194 364300 999200
rect 355968 999184 356020 999190
rect 358912 999184 358964 999190
rect 355968 999126 356020 999132
rect 358910 999152 358912 999161
rect 363052 999184 363104 999190
rect 358964 999152 358966 999161
rect 355980 993682 356008 999126
rect 358910 999087 358966 999096
rect 363050 999152 363052 999161
rect 363104 999152 363106 999161
rect 363050 999087 363106 999096
rect 364352 998238 364380 1001830
rect 364340 998232 364392 998238
rect 364340 998174 364392 998180
rect 364444 997966 364472 1001846
rect 365456 1000686 365484 1004634
rect 366376 1000822 366404 1004702
rect 366744 1004698 366772 1005042
rect 366732 1004692 366784 1004698
rect 366732 1004634 366784 1004640
rect 366364 1000816 366416 1000822
rect 366364 1000758 366416 1000764
rect 365444 1000680 365496 1000686
rect 365444 1000622 365496 1000628
rect 370424 1000618 370452 1005178
rect 371330 1004728 371386 1004737
rect 371330 1004663 371386 1004672
rect 370412 1000612 370464 1000618
rect 370412 1000554 370464 1000560
rect 368756 999728 368808 999734
rect 368756 999670 368808 999676
rect 368572 999660 368624 999666
rect 368572 999602 368624 999608
rect 365074 999560 365130 999569
rect 365074 999495 365076 999504
rect 365128 999495 365130 999504
rect 365076 999466 365128 999472
rect 367192 999456 367244 999462
rect 364706 999424 364762 999433
rect 367192 999398 367244 999404
rect 364706 999359 364708 999368
rect 364760 999359 364762 999368
rect 364708 999330 364760 999336
rect 365444 999320 365496 999326
rect 365442 999288 365444 999297
rect 365496 999288 365498 999297
rect 365442 999223 365498 999232
rect 367100 999184 367152 999190
rect 367100 999126 367152 999132
rect 364432 997960 364484 997966
rect 364432 997902 364484 997908
rect 366178 993712 366234 993721
rect 355968 993676 356020 993682
rect 366178 993647 366234 993656
rect 355968 993618 356020 993624
rect 366192 989738 366220 993647
rect 366180 989732 366232 989738
rect 366180 989674 366232 989680
rect 365444 989528 365496 989534
rect 365444 989470 365496 989476
rect 350448 985108 350500 985114
rect 350448 985050 350500 985056
rect 365456 983620 365484 989470
rect 367112 985046 367140 999126
rect 367204 988106 367232 999398
rect 368388 999252 368440 999258
rect 368388 999194 368440 999200
rect 368400 993410 368428 999194
rect 368584 993546 368612 999602
rect 368572 993540 368624 993546
rect 368572 993482 368624 993488
rect 368388 993404 368440 993410
rect 368388 993346 368440 993352
rect 367192 988100 367244 988106
rect 367192 988042 367244 988048
rect 367100 985040 367152 985046
rect 367100 984982 367152 984988
rect 368400 984910 368428 993346
rect 368584 984978 368612 993482
rect 368768 993478 368796 999670
rect 368940 999592 368992 999598
rect 368940 999534 368992 999540
rect 368952 997257 368980 999534
rect 369860 999388 369912 999394
rect 369860 999330 369912 999336
rect 368938 997248 368994 997257
rect 368938 997183 368994 997192
rect 368756 993472 368808 993478
rect 368756 993414 368808 993420
rect 368768 988038 368796 993414
rect 368756 988032 368808 988038
rect 368756 987974 368808 987980
rect 369872 987970 369900 999330
rect 371148 999320 371200 999326
rect 371148 999262 371200 999268
rect 371160 989670 371188 999262
rect 371148 989664 371200 989670
rect 371148 989606 371200 989612
rect 371344 989602 371372 1004663
rect 374288 1000482 374316 1005654
rect 377312 1005644 377364 1005650
rect 377312 1005586 377364 1005592
rect 377324 1001774 377352 1005586
rect 377956 1005508 378008 1005514
rect 377956 1005450 378008 1005456
rect 377312 1001768 377364 1001774
rect 377312 1001710 377364 1001716
rect 374276 1000476 374328 1000482
rect 374276 1000418 374328 1000424
rect 371516 999524 371568 999530
rect 371516 999466 371568 999472
rect 371332 989596 371384 989602
rect 371332 989538 371384 989544
rect 371528 989534 371556 999466
rect 377968 999002 377996 1005450
rect 423494 1005408 423550 1005417
rect 380808 1005372 380860 1005378
rect 423494 1005343 423496 1005352
rect 380808 1005314 380860 1005320
rect 423548 1005343 423550 1005352
rect 423496 1005314 423548 1005320
rect 378048 1005032 378100 1005038
rect 378048 1004974 378100 1004980
rect 378060 999190 378088 1004974
rect 380820 1001994 380848 1005314
rect 428372 1005304 428424 1005310
rect 428370 1005272 428372 1005281
rect 428424 1005272 428426 1005281
rect 428370 1005207 428426 1005216
rect 428830 1005136 428886 1005145
rect 428830 1005071 428832 1005080
rect 428884 1005071 428886 1005080
rect 428832 1005042 428884 1005048
rect 425520 1005032 425572 1005038
rect 425518 1005000 425520 1005009
rect 425572 1005000 425574 1005009
rect 383098 1004964 383150 1004970
rect 425518 1004935 425574 1004944
rect 426806 1005000 426862 1005009
rect 426806 1004935 426808 1004944
rect 383098 1004906 383150 1004912
rect 426860 1004935 426862 1004944
rect 426808 1004906 426860 1004912
rect 380820 1001966 380940 1001994
rect 378324 1001768 378376 1001774
rect 378324 1001710 378376 1001716
rect 378048 999184 378100 999190
rect 378048 999126 378100 999132
rect 377968 998974 378180 999002
rect 375196 998232 375248 998238
rect 375196 998174 375248 998180
rect 374460 997960 374512 997966
rect 374460 997902 374512 997908
rect 374472 993750 374500 997902
rect 374460 993744 374512 993750
rect 375208 993721 375236 998174
rect 378152 993857 378180 998974
rect 378336 993886 378364 1001710
rect 380912 1000414 380940 1001966
rect 380992 1000476 381044 1000482
rect 380992 1000418 381044 1000424
rect 380900 1000408 380952 1000414
rect 380900 1000350 380952 1000356
rect 381004 995518 381032 1000418
rect 383110 996441 383138 1004906
rect 427176 1004896 427228 1004902
rect 427174 1004864 427176 1004873
rect 427228 1004864 427230 1004873
rect 427174 1004799 427230 1004808
rect 427542 1004864 427598 1004873
rect 427542 1004799 427544 1004808
rect 427596 1004799 427598 1004808
rect 427544 1004770 427596 1004776
rect 419080 1004760 419132 1004766
rect 421840 1004760 421892 1004766
rect 419080 1004702 419132 1004708
rect 421838 1004728 421840 1004737
rect 422668 1004760 422720 1004766
rect 421892 1004728 421894 1004737
rect 383282 1004692 383334 1004698
rect 383282 1004634 383334 1004640
rect 383190 999184 383242 999190
rect 383190 999126 383242 999132
rect 383096 996432 383152 996441
rect 383096 996367 383152 996376
rect 383202 995586 383230 999126
rect 383294 995722 383322 1004634
rect 383558 1000816 383610 1000822
rect 383610 1000764 383782 1000770
rect 383558 1000758 383782 1000764
rect 383570 1000742 383782 1000758
rect 383374 1000680 383426 1000686
rect 383374 1000622 383426 1000628
rect 383386 995926 383414 1000622
rect 383466 1000612 383518 1000618
rect 383466 1000554 383518 1000560
rect 383478 995994 383506 1000554
rect 383558 1000544 383610 1000550
rect 383610 1000492 383690 1000498
rect 383558 1000486 383690 1000492
rect 383570 1000470 383690 1000486
rect 383558 1000408 383610 1000414
rect 383558 1000350 383610 1000356
rect 383466 995988 383518 995994
rect 383466 995930 383518 995936
rect 383374 995920 383426 995926
rect 383374 995862 383426 995868
rect 383282 995716 383334 995722
rect 383282 995658 383334 995664
rect 383570 995654 383598 1000350
rect 383662 995790 383690 1000470
rect 383754 995858 383782 1000742
rect 400036 999184 400088 999190
rect 400036 999126 400088 999132
rect 399944 999116 399996 999122
rect 399944 999058 399996 999064
rect 399956 997257 399984 999058
rect 399942 997248 399998 997257
rect 399942 997183 399998 997192
rect 400048 995858 400076 999126
rect 383742 995852 383794 995858
rect 383742 995794 383794 995800
rect 384396 995852 384448 995858
rect 384396 995794 384448 995800
rect 385684 995852 385736 995858
rect 385684 995794 385736 995800
rect 391940 995852 391992 995858
rect 391940 995794 391992 995800
rect 396632 995852 396684 995858
rect 396632 995794 396684 995800
rect 400036 995852 400088 995858
rect 400036 995794 400088 995800
rect 383650 995784 383702 995790
rect 383650 995726 383702 995732
rect 384408 995738 384436 995794
rect 384948 995784 385000 995790
rect 384408 995710 384698 995738
rect 385696 995738 385724 995794
rect 388166 995752 388222 995761
rect 385000 995732 385342 995738
rect 384948 995726 385342 995732
rect 384960 995710 385342 995726
rect 385696 995710 385986 995738
rect 391952 995738 391980 995794
rect 396644 995738 396672 995794
rect 388222 995710 388378 995738
rect 388640 995722 389022 995738
rect 388628 995716 389022 995722
rect 388166 995687 388222 995696
rect 388680 995710 389022 995716
rect 391952 995710 392150 995738
rect 396382 995710 396672 995738
rect 388628 995658 388680 995664
rect 383558 995648 383610 995654
rect 383558 995590 383610 995596
rect 387524 995648 387576 995654
rect 387576 995596 387826 995602
rect 387524 995590 387826 995596
rect 383190 995580 383242 995586
rect 387536 995574 387826 995590
rect 389376 995586 389666 995602
rect 389364 995580 389666 995586
rect 383190 995522 383242 995528
rect 389416 995574 389666 995580
rect 389364 995522 389416 995528
rect 380992 995512 381044 995518
rect 380992 995454 381044 995460
rect 393596 995512 393648 995518
rect 393648 995460 393990 995466
rect 393596 995454 393990 995460
rect 392688 993886 392716 995452
rect 378324 993880 378376 993886
rect 378138 993848 378194 993857
rect 378324 993822 378376 993828
rect 392676 993880 392728 993886
rect 392676 993822 392728 993828
rect 378138 993783 378194 993792
rect 393332 993750 393360 995452
rect 393608 995438 393990 995454
rect 393320 993744 393372 993750
rect 374460 993686 374512 993692
rect 375194 993712 375250 993721
rect 395172 993721 395200 995452
rect 397012 993857 397040 995452
rect 396998 993848 397054 993857
rect 396998 993783 397054 993792
rect 393320 993686 393372 993692
rect 395158 993712 395214 993721
rect 375194 993647 375250 993656
rect 398852 993682 398880 995452
rect 395158 993647 395214 993656
rect 398840 993676 398892 993682
rect 398840 993618 398892 993624
rect 381636 989732 381688 989738
rect 381636 989674 381688 989680
rect 371516 989528 371568 989534
rect 371516 989470 371568 989476
rect 369860 987964 369912 987970
rect 369860 987906 369912 987912
rect 368572 984972 368624 984978
rect 368572 984914 368624 984920
rect 368388 984904 368440 984910
rect 368388 984846 368440 984852
rect 381648 983620 381676 989674
rect 397828 989664 397880 989670
rect 397828 989606 397880 989612
rect 397840 983620 397868 989606
rect 414112 989596 414164 989602
rect 414112 989538 414164 989544
rect 414124 983620 414152 989538
rect 419092 984910 419120 1004702
rect 421838 1004663 421894 1004672
rect 422666 1004728 422668 1004737
rect 425152 1004760 425204 1004766
rect 422720 1004728 422722 1004737
rect 422666 1004663 422722 1004672
rect 425150 1004728 425152 1004737
rect 425204 1004728 425206 1004737
rect 425150 1004663 425206 1004672
rect 440160 1002046 440188 1005858
rect 440424 1005848 440476 1005854
rect 440424 1005790 440476 1005796
rect 440148 1002040 440200 1002046
rect 440148 1001982 440200 1001988
rect 440436 1001978 440464 1005790
rect 453948 1005304 454000 1005310
rect 453948 1005246 454000 1005252
rect 440424 1001972 440476 1001978
rect 440424 1001914 440476 1001920
rect 447140 1001904 447192 1001910
rect 447140 1001846 447192 1001852
rect 447324 1001904 447376 1001910
rect 447324 1001846 447376 1001852
rect 428004 1000680 428056 1000686
rect 426346 1000648 426402 1000657
rect 426346 1000583 426348 1000592
rect 426400 1000583 426402 1000592
rect 428002 1000648 428004 1000657
rect 428056 1000648 428058 1000657
rect 428002 1000583 428058 1000592
rect 426348 1000554 426400 1000560
rect 425980 1000544 426032 1000550
rect 425978 1000512 425980 1000521
rect 426032 1000512 426034 1000521
rect 425978 1000447 426034 1000456
rect 430856 999864 430908 999870
rect 430854 999832 430856 999841
rect 439824 999864 439876 999870
rect 430908 999832 430910 999841
rect 430854 999767 430910 999776
rect 431682 999832 431738 999841
rect 439824 999806 439876 999812
rect 431682 999767 431684 999776
rect 431736 999767 431738 999776
rect 437940 999796 437992 999802
rect 431684 999738 431736 999744
rect 437940 999738 437992 999744
rect 429200 999728 429252 999734
rect 429198 999696 429200 999705
rect 434628 999728 434680 999734
rect 429252 999696 429254 999705
rect 429198 999631 429254 999640
rect 430026 999696 430082 999705
rect 434628 999670 434680 999676
rect 430026 999631 430028 999640
rect 430080 999631 430082 999640
rect 430028 999602 430080 999608
rect 431224 999592 431276 999598
rect 431222 999560 431224 999569
rect 431276 999560 431278 999569
rect 431222 999495 431278 999504
rect 432418 999560 432474 999569
rect 432418 999495 432420 999504
rect 432472 999495 432474 999504
rect 432420 999466 432472 999472
rect 432880 999456 432932 999462
rect 429658 999424 429714 999433
rect 429658 999359 429660 999368
rect 429712 999359 429714 999368
rect 432878 999424 432880 999433
rect 432932 999424 432934 999433
rect 432878 999359 432934 999368
rect 433340 999388 433392 999394
rect 429660 999330 429712 999336
rect 433340 999330 433392 999336
rect 430396 999320 430448 999326
rect 430394 999288 430396 999297
rect 430448 999288 430450 999297
rect 430394 999223 430450 999232
rect 432050 999288 432106 999297
rect 432050 999223 432052 999232
rect 432104 999223 432106 999232
rect 432052 999194 432104 999200
rect 433352 993478 433380 999330
rect 433432 999320 433484 999326
rect 433432 999262 433484 999268
rect 433444 993546 433472 999262
rect 434640 993614 434668 999670
rect 434812 999660 434864 999666
rect 434812 999602 434864 999608
rect 433524 993608 433576 993614
rect 433524 993550 433576 993556
rect 434628 993608 434680 993614
rect 434628 993550 434680 993556
rect 433432 993540 433484 993546
rect 433432 993482 433484 993488
rect 433340 993472 433392 993478
rect 433340 993414 433392 993420
rect 430304 989528 430356 989534
rect 430304 989470 430356 989476
rect 419080 984904 419132 984910
rect 419080 984846 419132 984852
rect 430316 983620 430344 989470
rect 433536 987426 433564 993550
rect 434824 993546 434852 999602
rect 436192 999592 436244 999598
rect 436192 999534 436244 999540
rect 436100 999252 436152 999258
rect 436100 999194 436152 999200
rect 433616 993540 433668 993546
rect 433616 993482 433668 993488
rect 434812 993540 434864 993546
rect 434812 993482 434864 993488
rect 433524 987420 433576 987426
rect 433524 987362 433576 987368
rect 433628 984638 433656 993482
rect 436112 993410 436140 999194
rect 436204 999122 436232 999534
rect 437572 999524 437624 999530
rect 437572 999466 437624 999472
rect 437386 999152 437442 999161
rect 436192 999116 436244 999122
rect 437386 999087 437442 999096
rect 436192 999058 436244 999064
rect 436192 993472 436244 993478
rect 436192 993414 436244 993420
rect 436100 993404 436152 993410
rect 436100 993346 436152 993352
rect 433616 984632 433668 984638
rect 433616 984574 433668 984580
rect 436204 984570 436232 993414
rect 437400 989602 437428 999087
rect 437388 989596 437440 989602
rect 437388 989538 437440 989544
rect 437584 989534 437612 999466
rect 437756 999456 437808 999462
rect 437756 999398 437808 999404
rect 437768 989670 437796 999398
rect 437952 993478 437980 999738
rect 439836 997257 439864 999806
rect 444380 999184 444432 999190
rect 444380 999126 444432 999132
rect 439822 997248 439878 997257
rect 439822 997183 439878 997192
rect 437940 993472 437992 993478
rect 437940 993414 437992 993420
rect 444392 990690 444420 999126
rect 447152 993721 447180 1001846
rect 447336 995761 447364 1001846
rect 453960 999122 453988 1005246
rect 464252 1005100 464304 1005106
rect 464252 1005042 464304 1005048
rect 455604 1005032 455656 1005038
rect 455604 1004974 455656 1004980
rect 455512 1004964 455564 1004970
rect 455512 1004906 455564 1004912
rect 455420 1004896 455472 1004902
rect 455420 1004838 455472 1004844
rect 455432 1003338 455460 1004838
rect 455420 1003332 455472 1003338
rect 455420 1003274 455472 1003280
rect 455524 1003270 455552 1004906
rect 455512 1003264 455564 1003270
rect 455512 1003206 455564 1003212
rect 455616 1000754 455644 1004974
rect 455604 1000748 455656 1000754
rect 455604 1000690 455656 1000696
rect 464264 999190 464292 1005042
rect 466472 1004698 466500 1005994
rect 503352 1005848 503404 1005854
rect 502982 1005816 503038 1005825
rect 502982 1005751 502984 1005760
rect 503036 1005751 503038 1005760
rect 503350 1005816 503352 1005825
rect 503404 1005816 503406 1005825
rect 503350 1005751 503406 1005760
rect 502984 1005722 503036 1005728
rect 502524 1005712 502576 1005718
rect 502522 1005680 502524 1005689
rect 502576 1005680 502578 1005689
rect 502522 1005615 502578 1005624
rect 504546 1005680 504602 1005689
rect 504546 1005615 504548 1005624
rect 504600 1005615 504602 1005624
rect 517244 1005644 517296 1005650
rect 504548 1005586 504600 1005592
rect 517244 1005586 517296 1005592
rect 505836 1005576 505888 1005582
rect 505374 1005544 505430 1005553
rect 505374 1005479 505376 1005488
rect 505428 1005479 505430 1005488
rect 505834 1005544 505836 1005553
rect 505888 1005544 505890 1005553
rect 505834 1005479 505890 1005488
rect 505376 1005450 505428 1005456
rect 467840 1005372 467892 1005378
rect 467840 1005314 467892 1005320
rect 466552 1004828 466604 1004834
rect 466552 1004770 466604 1004776
rect 466460 1004692 466512 1004698
rect 466460 1004634 466512 1004640
rect 466564 1001978 466592 1004770
rect 467748 1004760 467800 1004766
rect 467748 1004702 467800 1004708
rect 466552 1001972 466604 1001978
rect 466552 1001914 466604 1001920
rect 464252 999184 464304 999190
rect 464252 999126 464304 999132
rect 453948 999116 454000 999122
rect 453948 999058 454000 999064
rect 462780 999116 462832 999122
rect 462780 999058 462832 999064
rect 447322 995752 447378 995761
rect 447322 995687 447378 995696
rect 447138 993712 447194 993721
rect 462792 993682 462820 999058
rect 467760 998374 467788 1004702
rect 467748 998368 467800 998374
rect 467748 998310 467800 998316
rect 467852 998170 467880 1005314
rect 504180 1005168 504232 1005174
rect 504178 1005136 504180 1005145
rect 504232 1005136 504234 1005145
rect 504178 1005071 504234 1005080
rect 505006 1005000 505062 1005009
rect 505006 1004935 505008 1004944
rect 505060 1004935 505062 1004944
rect 505008 1004906 505060 1004912
rect 500498 1004864 500554 1004873
rect 500498 1004799 500500 1004808
rect 500552 1004799 500554 1004808
rect 509332 1004828 509384 1004834
rect 500500 1004770 500552 1004776
rect 509332 1004770 509384 1004776
rect 496636 1004760 496688 1004766
rect 498844 1004760 498896 1004766
rect 496636 1004702 496688 1004708
rect 498842 1004728 498844 1004737
rect 499672 1004760 499724 1004766
rect 498896 1004728 498898 1004737
rect 472256 1004692 472308 1004698
rect 472256 1004634 472308 1004640
rect 469036 1003332 469088 1003338
rect 469036 1003274 469088 1003280
rect 469048 999134 469076 1003274
rect 469128 1003264 469180 1003270
rect 469128 1003206 469180 1003212
rect 469140 1001858 469168 1003206
rect 469140 1001830 469352 1001858
rect 469048 999106 469260 999134
rect 467840 998164 467892 998170
rect 467840 998106 467892 998112
rect 469232 995382 469260 999106
rect 469220 995376 469272 995382
rect 469220 995318 469272 995324
rect 469324 993818 469352 1001830
rect 472164 1000748 472216 1000754
rect 472164 1000690 472216 1000696
rect 470876 998368 470928 998374
rect 470876 998310 470928 998316
rect 469404 998164 469456 998170
rect 469404 998106 469456 998112
rect 469416 995450 469444 998106
rect 469404 995444 469456 995450
rect 469404 995386 469456 995392
rect 469312 993812 469364 993818
rect 469312 993754 469364 993760
rect 470888 993750 470916 998310
rect 472176 995994 472204 1000690
rect 472164 995988 472216 995994
rect 472164 995930 472216 995936
rect 472268 995654 472296 1004634
rect 472624 1001972 472676 1001978
rect 472624 1001914 472676 1001920
rect 472636 1001858 472664 1001914
rect 472636 1001830 472756 1001858
rect 472624 1000680 472676 1000686
rect 472624 1000622 472676 1000628
rect 472532 1000612 472584 1000618
rect 472532 1000554 472584 1000560
rect 472348 1000544 472400 1000550
rect 472348 1000486 472400 1000492
rect 472256 995648 472308 995654
rect 472256 995590 472308 995596
rect 472360 995586 472388 1000486
rect 472440 999184 472492 999190
rect 472440 999126 472492 999132
rect 472452 995722 472480 999126
rect 472544 995858 472572 1000554
rect 472532 995852 472584 995858
rect 472532 995794 472584 995800
rect 472636 995790 472664 1000622
rect 472728 995926 472756 1001830
rect 488908 999116 488960 999122
rect 488908 999058 488960 999064
rect 488920 997257 488948 999058
rect 488906 997248 488962 997257
rect 488906 997183 488962 997192
rect 472716 995920 472768 995926
rect 472716 995862 472768 995868
rect 474004 995852 474056 995858
rect 474004 995794 474056 995800
rect 476396 995852 476448 995858
rect 476396 995794 476448 995800
rect 477684 995852 477736 995858
rect 477684 995794 477736 995800
rect 472624 995784 472676 995790
rect 472624 995726 472676 995732
rect 473268 995784 473320 995790
rect 474016 995738 474044 995794
rect 476408 995738 476436 995794
rect 477696 995738 477724 995794
rect 481454 995752 481510 995761
rect 473320 995732 473662 995738
rect 473268 995726 473662 995732
rect 472440 995716 472492 995722
rect 473280 995710 473662 995726
rect 474016 995710 474306 995738
rect 474752 995722 474950 995738
rect 474740 995716 474950 995722
rect 472440 995658 472492 995664
rect 474792 995710 474950 995716
rect 476408 995710 476790 995738
rect 477696 995710 477986 995738
rect 481510 995710 481666 995738
rect 481454 995687 481510 995696
rect 474740 995658 474792 995664
rect 481916 995648 481968 995654
rect 476960 995586 477342 995602
rect 481968 995596 482310 995602
rect 481916 995590 482310 995596
rect 472348 995580 472400 995586
rect 472348 995522 472400 995528
rect 476948 995580 477342 995586
rect 477000 995574 477342 995580
rect 481928 995574 482310 995590
rect 482664 995586 482954 995602
rect 482652 995580 482954 995586
rect 476948 995522 477000 995528
rect 482704 995574 482954 995580
rect 482652 995522 482704 995528
rect 470876 993744 470928 993750
rect 478616 993721 478644 995452
rect 480824 995438 481114 995466
rect 480824 995382 480852 995438
rect 480812 995376 480864 995382
rect 480812 995318 480864 995324
rect 484136 993750 484164 995452
rect 484124 993744 484176 993750
rect 470876 993686 470928 993692
rect 478602 993712 478658 993721
rect 447138 993647 447194 993656
rect 462780 993676 462832 993682
rect 484124 993686 484176 993692
rect 478602 993647 478658 993656
rect 462780 993618 462832 993624
rect 444380 990684 444432 990690
rect 444380 990626 444432 990632
rect 446220 990684 446272 990690
rect 446220 990626 446272 990632
rect 437756 989664 437808 989670
rect 437756 989606 437808 989612
rect 437572 989528 437624 989534
rect 437572 989470 437624 989476
rect 436192 984564 436244 984570
rect 436192 984506 436244 984512
rect 446232 983634 446260 990626
rect 462780 989664 462832 989670
rect 462780 989606 462832 989612
rect 446232 983606 446522 983634
rect 462792 983620 462820 989606
rect 478972 989596 479024 989602
rect 478972 989538 479024 989544
rect 478984 983620 479012 989538
rect 485332 989505 485360 995452
rect 485976 993682 486004 995452
rect 487816 993818 487844 995452
rect 487804 993812 487856 993818
rect 487804 993754 487856 993760
rect 485964 993676 486016 993682
rect 485964 993618 486016 993624
rect 495164 989528 495216 989534
rect 485318 989496 485374 989505
rect 495164 989470 495216 989476
rect 485318 989431 485374 989440
rect 495176 983620 495204 989470
rect 496648 984570 496676 1004702
rect 498842 1004663 498898 1004672
rect 499670 1004728 499672 1004737
rect 501696 1004760 501748 1004766
rect 499724 1004728 499726 1004737
rect 499670 1004663 499726 1004672
rect 501694 1004728 501696 1004737
rect 509240 1004760 509292 1004766
rect 501748 1004728 501750 1004737
rect 501694 1004663 501750 1004672
rect 502154 1004728 502210 1004737
rect 509240 1004702 509292 1004708
rect 502154 1004663 502156 1004672
rect 502208 1004663 502210 1004672
rect 509148 1004692 509200 1004698
rect 502156 1004634 502208 1004640
rect 509148 1004634 509200 1004640
rect 508686 999832 508742 999841
rect 508686 999767 508688 999776
rect 508740 999767 508742 999776
rect 508688 999738 508740 999744
rect 506204 999728 506256 999734
rect 506202 999696 506204 999705
rect 506256 999696 506258 999705
rect 506202 999631 506258 999640
rect 508226 999696 508282 999705
rect 508226 999631 508228 999640
rect 508280 999631 508282 999640
rect 508228 999602 508280 999608
rect 507032 999592 507084 999598
rect 507030 999560 507032 999569
rect 507084 999560 507086 999569
rect 507030 999495 507086 999504
rect 507858 999560 507914 999569
rect 507858 999495 507860 999504
rect 507912 999495 507914 999504
rect 507860 999466 507912 999472
rect 506664 999456 506716 999462
rect 506662 999424 506664 999433
rect 506716 999424 506718 999433
rect 506662 999359 506718 999368
rect 509054 999424 509110 999433
rect 509054 999359 509056 999368
rect 509108 999359 509110 999368
rect 509056 999330 509108 999336
rect 507400 999320 507452 999326
rect 500866 999288 500922 999297
rect 500866 999223 500868 999232
rect 500920 999223 500922 999232
rect 507398 999288 507400 999297
rect 507452 999288 507454 999297
rect 507398 999223 507454 999232
rect 507860 999252 507912 999258
rect 500868 999194 500920 999200
rect 507860 999194 507912 999200
rect 499488 999184 499540 999190
rect 503352 999184 503404 999190
rect 499488 999126 499540 999132
rect 503350 999152 503352 999161
rect 503404 999152 503406 999161
rect 499500 993682 499528 999126
rect 503350 999087 503406 999096
rect 507872 998850 507900 999194
rect 509160 998918 509188 1004634
rect 509252 998986 509280 1004702
rect 509344 999054 509372 1004770
rect 515220 999796 515272 999802
rect 515220 999738 515272 999744
rect 512092 999728 512144 999734
rect 512092 999670 512144 999676
rect 511908 999592 511960 999598
rect 511908 999534 511960 999540
rect 510712 999456 510764 999462
rect 510712 999398 510764 999404
rect 510620 999320 510672 999326
rect 509514 999288 509570 999297
rect 510620 999262 510672 999268
rect 509514 999223 509516 999232
rect 509568 999223 509570 999232
rect 509516 999194 509568 999200
rect 509884 999184 509936 999190
rect 509882 999152 509884 999161
rect 509936 999152 509938 999161
rect 509882 999087 509938 999096
rect 509332 999048 509384 999054
rect 509332 998990 509384 998996
rect 509240 998980 509292 998986
rect 509240 998922 509292 998928
rect 509148 998912 509200 998918
rect 509148 998854 509200 998860
rect 507860 998844 507912 998850
rect 507860 998786 507912 998792
rect 499488 993676 499540 993682
rect 499488 993618 499540 993624
rect 510632 993546 510660 999262
rect 510724 993614 510752 999398
rect 511920 993614 511948 999534
rect 510712 993608 510764 993614
rect 510712 993550 510764 993556
rect 510896 993608 510948 993614
rect 510896 993550 510948 993556
rect 511908 993608 511960 993614
rect 511908 993550 511960 993556
rect 510620 993540 510672 993546
rect 510620 993482 510672 993488
rect 510804 993540 510856 993546
rect 510804 993482 510856 993488
rect 496636 984564 496688 984570
rect 496636 984506 496688 984512
rect 510816 984502 510844 993482
rect 510804 984496 510856 984502
rect 510804 984438 510856 984444
rect 510908 984434 510936 993550
rect 512104 993546 512132 999670
rect 513472 999660 513524 999666
rect 513472 999602 513524 999608
rect 512276 999524 512328 999530
rect 512276 999466 512328 999472
rect 512288 996188 512316 999466
rect 513380 999388 513432 999394
rect 513380 999330 513432 999336
rect 512276 996182 512328 996188
rect 512276 996124 512328 996130
rect 512092 993540 512144 993546
rect 512092 993482 512144 993488
rect 513392 993478 513420 999330
rect 513484 999122 513512 999602
rect 513643 999329 515076 999357
rect 513643 999161 513671 999329
rect 514668 999252 514720 999258
rect 514668 999194 514720 999200
rect 513629 999152 513685 999161
rect 513472 999116 513524 999122
rect 513629 999087 513685 999096
rect 513472 999058 513524 999064
rect 513380 993472 513432 993478
rect 513380 993414 513432 993420
rect 513472 993472 513524 993478
rect 513472 993414 513524 993420
rect 511446 989496 511502 989505
rect 511446 989431 511502 989440
rect 510896 984428 510948 984434
rect 510896 984370 510948 984376
rect 511460 983620 511488 989431
rect 513484 984366 513512 993414
rect 514680 989534 514708 999194
rect 514852 999184 514904 999190
rect 514852 999126 514904 999132
rect 514864 989670 514892 999126
rect 514852 989664 514904 989670
rect 514852 989606 514904 989612
rect 515048 989602 515076 999329
rect 515232 993478 515260 999738
rect 517256 999161 517284 1005586
rect 517348 1004698 517376 1007354
rect 520188 1005848 520240 1005854
rect 520188 1005790 520240 1005796
rect 520004 1005780 520056 1005786
rect 520004 1005722 520056 1005728
rect 519176 1005712 519228 1005718
rect 519176 1005654 519228 1005660
rect 517612 1005576 517664 1005582
rect 517612 1005518 517664 1005524
rect 517428 1005508 517480 1005514
rect 517428 1005450 517480 1005456
rect 517336 1004692 517388 1004698
rect 517336 1004634 517388 1004640
rect 517242 999152 517298 999161
rect 517242 999087 517298 999096
rect 517440 993721 517468 1005450
rect 517624 995625 517652 1005518
rect 519188 1001978 519216 1005654
rect 519176 1001972 519228 1001978
rect 519176 1001914 519228 1001920
rect 520016 999297 520044 1005722
rect 520002 999288 520058 999297
rect 520002 999223 520058 999232
rect 520200 995761 520228 1005790
rect 520372 1005168 520424 1005174
rect 520372 1005110 520424 1005116
rect 551926 1005136 551982 1005145
rect 520186 995752 520242 995761
rect 520186 995687 520242 995696
rect 517610 995616 517666 995625
rect 517610 995551 517666 995560
rect 520384 995489 520412 1005110
rect 551926 1005071 551928 1005080
rect 551980 1005071 551982 1005080
rect 568580 1005100 568632 1005106
rect 551928 1005042 551980 1005048
rect 568580 1005042 568632 1005048
rect 554778 1005000 554834 1005009
rect 522948 1004964 523000 1004970
rect 522948 1004906 523000 1004912
rect 551652 1004964 551704 1004970
rect 554778 1004935 554780 1004944
rect 551652 1004906 551704 1004912
rect 554832 1004935 554834 1004944
rect 554780 1004906 554832 1004912
rect 521292 999048 521344 999054
rect 521292 998990 521344 998996
rect 521304 995586 521332 998990
rect 521476 998980 521528 998986
rect 521476 998922 521528 998928
rect 521384 998912 521436 998918
rect 521384 998854 521436 998860
rect 521292 995580 521344 995586
rect 521292 995522 521344 995528
rect 520370 995480 520426 995489
rect 520370 995415 520426 995424
rect 521396 993818 521424 998854
rect 521488 995654 521516 998922
rect 521568 998844 521620 998850
rect 521568 998786 521620 998792
rect 521580 995722 521608 998786
rect 522960 995858 522988 1004906
rect 549444 1004760 549496 1004766
rect 546406 1004728 546462 1004737
rect 523592 1004692 523644 1004698
rect 546406 1004663 546462 1004672
rect 549442 1004728 549444 1004737
rect 550272 1004760 550324 1004766
rect 549496 1004728 549498 1004737
rect 549442 1004663 549498 1004672
rect 550270 1004728 550272 1004737
rect 551100 1004760 551152 1004766
rect 550324 1004728 550326 1004737
rect 550270 1004663 550326 1004672
rect 551098 1004728 551100 1004737
rect 551152 1004728 551154 1004737
rect 551098 1004663 551154 1004672
rect 523592 1004634 523644 1004640
rect 523604 995926 523632 1004634
rect 523776 1001972 523828 1001978
rect 523776 1001914 523828 1001920
rect 523592 995920 523644 995926
rect 523592 995862 523644 995868
rect 522948 995852 523000 995858
rect 522948 995794 523000 995800
rect 523788 995790 523816 1001914
rect 540336 999320 540388 999326
rect 523866 999288 523922 999297
rect 540336 999262 540388 999268
rect 523866 999223 523922 999232
rect 523880 996577 523908 999223
rect 524050 999152 524106 999161
rect 524050 999087 524106 999096
rect 523866 996568 523922 996577
rect 523866 996503 523922 996512
rect 524064 996441 524092 999087
rect 524050 996432 524106 996441
rect 524050 996367 524106 996376
rect 540348 995858 540376 999262
rect 524788 995852 524840 995858
rect 524788 995794 524840 995800
rect 530124 995852 530176 995858
rect 530124 995794 530176 995800
rect 537024 995852 537076 995858
rect 537024 995794 537076 995800
rect 540336 995852 540388 995858
rect 540336 995794 540388 995800
rect 523776 995784 523828 995790
rect 523776 995726 523828 995732
rect 524800 995738 524828 995794
rect 529020 995784 529072 995790
rect 525430 995752 525486 995761
rect 521568 995716 521620 995722
rect 524800 995710 525090 995738
rect 528006 995752 528062 995761
rect 525486 995710 525734 995738
rect 525430 995687 525486 995696
rect 528558 995752 528614 995761
rect 528062 995710 528218 995738
rect 528006 995687 528062 995696
rect 528614 995710 528770 995738
rect 530136 995738 530164 995794
rect 537036 995738 537064 995794
rect 529072 995732 529414 995738
rect 529020 995726 529414 995732
rect 529032 995710 529414 995726
rect 530058 995710 530164 995738
rect 532712 995722 533094 995738
rect 532700 995716 533094 995722
rect 528558 995687 528614 995696
rect 521568 995658 521620 995664
rect 532752 995710 533094 995716
rect 536774 995710 537064 995738
rect 532700 995658 532752 995664
rect 521476 995648 521528 995654
rect 533436 995648 533488 995654
rect 521476 995590 521528 995596
rect 526074 995616 526130 995625
rect 526130 995574 526378 995602
rect 533488 995596 533738 995602
rect 533436 995590 533738 995596
rect 533448 995574 533738 995590
rect 534000 995586 534382 995602
rect 533988 995580 534382 995586
rect 526074 995551 526130 995560
rect 534040 995574 534382 995580
rect 533988 995522 534040 995528
rect 532146 995480 532202 995489
rect 532202 995438 532542 995466
rect 532146 995415 532202 995424
rect 535564 993818 535592 995452
rect 521384 993812 521436 993818
rect 521384 993754 521436 993760
rect 535552 993812 535604 993818
rect 535552 993754 535604 993760
rect 537404 993721 537432 995452
rect 517426 993712 517482 993721
rect 517426 993647 517482 993656
rect 537390 993712 537446 993721
rect 539244 993682 539272 995452
rect 537390 993647 537446 993656
rect 539232 993676 539284 993682
rect 539232 993618 539284 993624
rect 515220 993472 515272 993478
rect 515220 993414 515272 993420
rect 527640 989664 527692 989670
rect 527640 989606 527692 989612
rect 515036 989596 515088 989602
rect 515036 989538 515088 989544
rect 514668 989528 514720 989534
rect 514668 989470 514720 989476
rect 513472 984360 513524 984366
rect 513472 984302 513524 984308
rect 527652 983620 527680 989606
rect 543832 989596 543884 989602
rect 543832 989538 543884 989544
rect 543844 983620 543872 989538
rect 546420 984366 546448 1004663
rect 548892 999252 548944 999258
rect 548892 999194 548944 999200
rect 548904 997626 548932 999194
rect 549076 999184 549128 999190
rect 549076 999126 549128 999132
rect 549088 997830 549116 999126
rect 549076 997824 549128 997830
rect 549076 997766 549128 997772
rect 548892 997620 548944 997626
rect 548892 997562 548944 997568
rect 551664 993682 551692 1004906
rect 553124 1004896 553176 1004902
rect 553122 1004864 553124 1004873
rect 555516 1004896 555568 1004902
rect 553176 1004864 553178 1004873
rect 553122 1004799 553178 1004808
rect 553950 1004864 554006 1004873
rect 555516 1004838 555568 1004844
rect 567474 1004864 567530 1004873
rect 553950 1004799 553952 1004808
rect 554004 1004799 554006 1004808
rect 553952 1004770 554004 1004776
rect 552756 1004760 552808 1004766
rect 552754 1004728 552756 1004737
rect 552808 1004728 552810 1004737
rect 555146 1004728 555202 1004737
rect 552754 1004663 552810 1004672
rect 554700 1004686 555146 1004714
rect 553492 1003536 553544 1003542
rect 553490 1003504 553492 1003513
rect 553544 1003504 553546 1003513
rect 553490 1003439 553546 1003448
rect 554700 1003338 554728 1004686
rect 555146 1004663 555202 1004672
rect 555528 1003950 555556 1004838
rect 555700 1004828 555752 1004834
rect 567474 1004799 567530 1004808
rect 555700 1004770 555752 1004776
rect 555712 1004222 555740 1004770
rect 555700 1004216 555752 1004222
rect 555700 1004158 555752 1004164
rect 555516 1003944 555568 1003950
rect 555516 1003886 555568 1003892
rect 556160 1003536 556212 1003542
rect 556160 1003478 556212 1003484
rect 554688 1003332 554740 1003338
rect 554688 1003274 554740 1003280
rect 554320 1003264 554372 1003270
rect 554318 1003232 554320 1003241
rect 554372 1003232 554374 1003241
rect 554318 1003167 554374 1003176
rect 556172 1001298 556200 1003478
rect 556160 1001292 556212 1001298
rect 556160 1001234 556212 1001240
rect 555974 1000104 556030 1000113
rect 555974 1000039 555976 1000048
rect 556028 1000039 556030 1000048
rect 567016 1000068 567068 1000074
rect 555976 1000010 556028 1000016
rect 567016 1000010 567068 1000016
rect 564256 1000000 564308 1000006
rect 558458 999968 558514 999977
rect 564256 999942 564308 999948
rect 558458 999903 558460 999912
rect 558512 999903 558514 999912
rect 558460 999874 558512 999880
rect 560852 999864 560904 999870
rect 556342 999832 556398 999841
rect 556342 999767 556344 999776
rect 556396 999767 556398 999776
rect 560850 999832 560852 999841
rect 560904 999832 560906 999841
rect 560850 999767 560906 999776
rect 562140 999796 562192 999802
rect 556344 999738 556396 999744
rect 562140 999738 562192 999744
rect 560484 999728 560536 999734
rect 559194 999696 559250 999705
rect 559194 999631 559196 999640
rect 559248 999631 559250 999640
rect 560482 999696 560484 999705
rect 560536 999696 560538 999705
rect 560482 999631 560538 999640
rect 559196 999602 559248 999608
rect 560024 999592 560076 999598
rect 557998 999560 558054 999569
rect 557998 999495 558000 999504
rect 558052 999495 558054 999504
rect 560022 999560 560024 999569
rect 560076 999560 560078 999569
rect 560022 999495 560078 999504
rect 558000 999466 558052 999472
rect 556804 999456 556856 999462
rect 556802 999424 556804 999433
rect 561772 999456 561824 999462
rect 556856 999424 556858 999433
rect 556802 999359 556858 999368
rect 557170 999424 557226 999433
rect 561772 999398 561824 999404
rect 557170 999359 557172 999368
rect 557224 999359 557226 999368
rect 557172 999330 557224 999336
rect 558828 999320 558880 999326
rect 554318 999288 554374 999297
rect 554318 999223 554320 999232
rect 554372 999223 554374 999232
rect 558826 999288 558828 999297
rect 558880 999288 558882 999297
rect 558826 999223 558882 999232
rect 559654 999288 559710 999297
rect 559654 999223 559656 999232
rect 554320 999194 554372 999200
rect 559708 999223 559710 999232
rect 561310 999288 561366 999297
rect 561366 999246 561720 999274
rect 561310 999223 561366 999232
rect 559656 999194 559708 999200
rect 561692 999190 561720 999246
rect 551928 999184 551980 999190
rect 551926 999152 551928 999161
rect 557632 999184 557684 999190
rect 551980 999152 551982 999161
rect 551926 999087 551982 999096
rect 557630 999152 557632 999161
rect 561588 999184 561640 999190
rect 557684 999152 557686 999161
rect 561588 999126 561640 999132
rect 561680 999184 561732 999190
rect 561680 999126 561732 999132
rect 557630 999087 557686 999096
rect 551652 993676 551704 993682
rect 551652 993618 551704 993624
rect 560116 989528 560168 989534
rect 560116 989470 560168 989476
rect 546408 984360 546460 984366
rect 546408 984302 546460 984308
rect 560128 983620 560156 989470
rect 561600 985833 561628 999126
rect 561784 993721 561812 999398
rect 561956 999388 562008 999394
rect 561956 999330 562008 999336
rect 561968 997694 561996 999330
rect 561956 997688 562008 997694
rect 561956 997630 562008 997636
rect 562152 997354 562180 999738
rect 563060 999524 563112 999530
rect 563060 999466 563112 999472
rect 562140 997348 562192 997354
rect 562140 997290 562192 997296
rect 561770 993712 561826 993721
rect 561770 993647 561826 993656
rect 563072 993546 563100 999466
rect 563152 999320 563204 999326
rect 563152 999262 563204 999268
rect 563164 993614 563192 999262
rect 563244 999252 563296 999258
rect 563244 999194 563296 999200
rect 563256 996188 563284 999194
rect 563244 996182 563296 996188
rect 563244 996124 563296 996130
rect 563152 993608 563204 993614
rect 563152 993550 563204 993556
rect 563060 993540 563112 993546
rect 563060 993482 563112 993488
rect 564268 990826 564296 999942
rect 564532 999932 564584 999938
rect 564532 999874 564584 999880
rect 564348 999660 564400 999666
rect 564348 999602 564400 999608
rect 564256 990820 564308 990826
rect 564256 990762 564308 990768
rect 561034 985824 561090 985833
rect 561034 985759 561090 985768
rect 561586 985824 561642 985833
rect 561586 985759 561642 985768
rect 561048 984094 561076 985759
rect 564360 984094 564388 999602
rect 564544 999134 564572 999874
rect 565820 999728 565872 999734
rect 565820 999670 565872 999676
rect 564716 999592 564768 999598
rect 564716 999534 564768 999540
rect 564452 999106 564572 999134
rect 564452 985969 564480 999106
rect 564438 985960 564494 985969
rect 564438 985895 564494 985904
rect 561036 984088 561088 984094
rect 561036 984030 561088 984036
rect 564348 984088 564400 984094
rect 564348 984030 564400 984036
rect 564452 983958 564480 985895
rect 564728 985522 564756 999534
rect 565832 993478 565860 999670
rect 567028 993753 567056 1000010
rect 567292 999864 567344 999870
rect 567292 999806 567344 999812
rect 567108 999184 567160 999190
rect 567108 999126 567160 999132
rect 567014 993744 567070 993753
rect 567014 993679 567070 993688
rect 565820 993472 565872 993478
rect 565820 993414 565872 993420
rect 567120 989670 567148 999126
rect 567108 989664 567160 989670
rect 567108 989606 567160 989612
rect 567304 989534 567332 999806
rect 567488 989602 567516 1004799
rect 568592 1002114 568620 1005042
rect 571248 1004896 571300 1004902
rect 571248 1004838 571300 1004844
rect 569868 1004216 569920 1004222
rect 569868 1004158 569920 1004164
rect 568580 1002108 568632 1002114
rect 568580 1002050 568632 1002056
rect 569880 997490 569908 1004158
rect 569960 1003944 570012 1003950
rect 569960 1003886 570012 1003892
rect 569868 997484 569920 997490
rect 569868 997426 569920 997432
rect 569972 993857 570000 1003886
rect 571260 1001858 571288 1004838
rect 571616 1003332 571668 1003338
rect 571616 1003274 571668 1003280
rect 571432 1003264 571484 1003270
rect 571432 1003206 571484 1003212
rect 571260 1001830 571380 1001858
rect 571248 1001292 571300 1001298
rect 571248 1001234 571300 1001240
rect 571260 996554 571288 1001234
rect 571352 997558 571380 1001830
rect 571340 997552 571392 997558
rect 571340 997494 571392 997500
rect 571444 997422 571472 1003206
rect 571524 1002108 571576 1002114
rect 571524 1002050 571576 1002056
rect 571536 997762 571564 1002050
rect 571524 997756 571576 997762
rect 571524 997698 571576 997704
rect 571432 997416 571484 997422
rect 571432 997358 571484 997364
rect 571260 996526 571380 996554
rect 571352 994129 571380 996526
rect 571338 994120 571394 994129
rect 571338 994055 571394 994064
rect 569958 993848 570014 993857
rect 569958 993783 570014 993792
rect 571628 993750 571656 1003274
rect 590660 1001972 590712 1001978
rect 590660 1001914 590712 1001920
rect 625804 1001972 625856 1001978
rect 625804 1001914 625856 1001920
rect 575572 997824 575624 997830
rect 575572 997766 575624 997772
rect 575584 994265 575612 997766
rect 590672 997694 590700 1001914
rect 625816 1001858 625844 1001914
rect 625816 1001830 625936 1001858
rect 590752 999456 590804 999462
rect 590752 999398 590804 999404
rect 625436 999456 625488 999462
rect 625436 999398 625488 999404
rect 590660 997688 590712 997694
rect 590660 997630 590712 997636
rect 590764 997558 590792 999398
rect 607128 999320 607180 999326
rect 607128 999262 607180 999268
rect 602252 999252 602304 999258
rect 602252 999194 602304 999200
rect 590752 997552 590804 997558
rect 590752 997494 590804 997500
rect 602264 997422 602292 999194
rect 607140 997490 607168 999262
rect 612740 999184 612792 999190
rect 612740 999126 612792 999132
rect 612752 997626 612780 999126
rect 623780 997756 623832 997762
rect 623780 997698 623832 997704
rect 612740 997620 612792 997626
rect 612740 997562 612792 997568
rect 607128 997484 607180 997490
rect 607128 997426 607180 997432
rect 602252 997416 602304 997422
rect 602252 997358 602304 997364
rect 623688 997348 623740 997354
rect 623688 997290 623740 997296
rect 623700 995858 623728 997290
rect 623688 995852 623740 995858
rect 623688 995794 623740 995800
rect 623792 995586 623820 997698
rect 625448 995654 625476 999398
rect 625620 999320 625672 999326
rect 625620 999262 625672 999268
rect 625632 995994 625660 999262
rect 625712 999252 625764 999258
rect 625712 999194 625764 999200
rect 625620 995988 625672 995994
rect 625620 995930 625672 995936
rect 625724 995722 625752 999194
rect 625804 999184 625856 999190
rect 625804 999126 625856 999132
rect 625816 995790 625844 999126
rect 625908 995926 625936 1001830
rect 625896 995920 625948 995926
rect 625896 995862 625948 995868
rect 626540 995852 626592 995858
rect 626540 995794 626592 995800
rect 627828 995852 627880 995858
rect 627828 995794 627880 995800
rect 630864 995852 630916 995858
rect 630864 995794 630916 995800
rect 625804 995784 625856 995790
rect 625804 995726 625856 995732
rect 626552 995738 626580 995794
rect 627184 995784 627236 995790
rect 625712 995716 625764 995722
rect 626552 995710 626888 995738
rect 627840 995738 627868 995794
rect 630876 995738 630904 995794
rect 627236 995732 627532 995738
rect 627184 995726 627532 995732
rect 627196 995710 627532 995726
rect 627840 995710 628176 995738
rect 630232 995722 630568 995738
rect 630220 995716 630568 995722
rect 625712 995658 625764 995664
rect 630272 995710 630568 995716
rect 630876 995710 631212 995738
rect 630220 995658 630272 995664
rect 625436 995648 625488 995654
rect 625436 995590 625488 995596
rect 631508 995648 631560 995654
rect 631560 995596 631856 995602
rect 631508 995590 631856 995596
rect 623780 995580 623832 995586
rect 631520 995574 631856 995590
rect 635844 995586 636180 995602
rect 635832 995580 636180 995586
rect 623780 995522 623832 995528
rect 635884 995574 636180 995580
rect 635832 995522 635884 995528
rect 629680 995438 630016 995466
rect 634004 995438 634340 995466
rect 634832 995438 634892 995466
rect 635200 995438 635536 995466
rect 637040 995438 637376 995466
rect 575570 994256 575626 994265
rect 575570 994191 575626 994200
rect 629680 993993 629708 995438
rect 629666 993984 629722 993993
rect 629666 993919 629722 993928
rect 634004 993750 634032 995438
rect 634832 994265 634860 995438
rect 634818 994256 634874 994265
rect 634818 994191 634874 994200
rect 635200 993857 635228 995438
rect 637040 994129 637068 995438
rect 638558 995217 638586 995452
rect 638880 995438 639216 995466
rect 640720 995438 641056 995466
rect 638544 995208 638600 995217
rect 638544 995143 638600 995152
rect 637026 994120 637082 994129
rect 637026 994055 637082 994064
rect 635186 993848 635242 993857
rect 635186 993783 635242 993792
rect 571616 993744 571668 993750
rect 571616 993686 571668 993692
rect 633992 993744 634044 993750
rect 638880 993721 638908 995438
rect 633992 993686 634044 993692
rect 638866 993712 638922 993721
rect 640720 993682 640748 995438
rect 638866 993647 638922 993656
rect 640708 993676 640760 993682
rect 640708 993618 640760 993624
rect 576308 990820 576360 990826
rect 576308 990762 576360 990768
rect 567476 989596 567528 989602
rect 567476 989538 567528 989544
rect 567292 989528 567344 989534
rect 567292 989470 567344 989476
rect 564532 985516 564584 985522
rect 564532 985458 564584 985464
rect 564716 985516 564768 985522
rect 564716 985458 564768 985464
rect 564544 984026 564572 985458
rect 564532 984020 564584 984026
rect 564532 983962 564584 983968
rect 564440 983952 564492 983958
rect 564440 983894 564492 983900
rect 576320 983620 576348 990762
rect 641166 990584 641222 990593
rect 641166 990519 641222 990528
rect 592500 989664 592552 989670
rect 592500 989606 592552 989612
rect 592512 983620 592540 989606
rect 608784 989596 608836 989602
rect 608784 989538 608836 989544
rect 608796 983620 608824 989538
rect 624976 989528 625028 989534
rect 624976 989470 625028 989476
rect 624988 983620 625016 989470
rect 641180 983620 641208 990519
rect 666560 989460 666612 989466
rect 666560 989402 666612 989408
rect 651380 987624 651432 987630
rect 651380 987566 651432 987572
rect 649908 984088 649960 984094
rect 649908 984030 649960 984036
rect 63132 983000 63184 983006
rect 63132 982942 63184 982948
rect 62948 982932 63000 982938
rect 62948 982874 63000 982880
rect 62854 814192 62910 814201
rect 62854 814127 62910 814136
rect 62856 772880 62908 772886
rect 62856 772822 62908 772828
rect 62764 598936 62816 598942
rect 62764 598878 62816 598884
rect 62764 427848 62816 427854
rect 62764 427790 62816 427796
rect 62776 278322 62804 427790
rect 62764 278316 62816 278322
rect 62764 278258 62816 278264
rect 62670 278216 62726 278225
rect 62670 278151 62726 278160
rect 62486 278080 62542 278089
rect 62486 278015 62542 278024
rect 62868 277953 62896 772822
rect 62960 681698 62988 982874
rect 63038 730280 63094 730289
rect 63038 730215 63094 730224
rect 62948 681692 63000 681698
rect 62948 681634 63000 681640
rect 62946 427952 63002 427961
rect 62946 427887 63002 427896
rect 62960 278254 62988 427887
rect 62948 278248 63000 278254
rect 62948 278190 63000 278196
rect 62854 277944 62910 277953
rect 62854 277879 62910 277888
rect 63052 277817 63080 730215
rect 63144 684321 63172 982942
rect 649920 935678 649948 984030
rect 649908 935672 649960 935678
rect 649908 935614 649960 935620
rect 63130 684312 63186 684321
rect 63130 684247 63186 684256
rect 63222 386744 63278 386753
rect 63222 386679 63278 386688
rect 63132 386436 63184 386442
rect 63132 386378 63184 386384
rect 63144 278118 63172 386378
rect 63132 278112 63184 278118
rect 63132 278054 63184 278060
rect 63236 278050 63264 386679
rect 63314 383752 63370 383761
rect 63314 383687 63370 383696
rect 63224 278044 63276 278050
rect 63224 277986 63276 277992
rect 63328 277982 63356 383687
rect 63316 277976 63368 277982
rect 63316 277918 63368 277924
rect 63038 277808 63094 277817
rect 63038 277743 63094 277752
rect 65904 271862 65932 277780
rect 67008 271930 67036 277780
rect 66996 271924 67048 271930
rect 66996 271866 67048 271872
rect 65892 271856 65944 271862
rect 65892 271798 65944 271804
rect 68204 266354 68232 277780
rect 69400 269113 69428 277780
rect 70596 271833 70624 277780
rect 70582 271824 70638 271833
rect 70582 271759 70638 271768
rect 71792 269210 71820 277780
rect 71780 269204 71832 269210
rect 71780 269146 71832 269152
rect 69386 269104 69442 269113
rect 69386 269039 69442 269048
rect 72988 266490 73016 277780
rect 74092 269414 74120 277780
rect 75288 271998 75316 277780
rect 75276 271992 75328 271998
rect 76484 271969 76512 277780
rect 75276 271934 75328 271940
rect 76470 271960 76526 271969
rect 76470 271895 76526 271904
rect 74080 269408 74132 269414
rect 74080 269350 74132 269356
rect 77680 269249 77708 277780
rect 78876 269385 78904 277780
rect 78862 269376 78918 269385
rect 80072 269346 80100 277780
rect 78862 269311 78918 269320
rect 80060 269340 80112 269346
rect 80060 269282 80112 269288
rect 81268 269278 81296 277780
rect 81256 269272 81308 269278
rect 77666 269240 77722 269249
rect 81256 269214 81308 269220
rect 77666 269175 77722 269184
rect 82372 268054 82400 277780
rect 83568 272105 83596 277780
rect 83554 272096 83610 272105
rect 83554 272031 83610 272040
rect 84764 269521 84792 277780
rect 85960 272241 85988 277780
rect 85946 272232 86002 272241
rect 85946 272167 86002 272176
rect 87156 269657 87184 277780
rect 87142 269648 87198 269657
rect 87142 269583 87198 269592
rect 84750 269512 84806 269521
rect 84750 269447 84806 269456
rect 82360 268048 82412 268054
rect 82360 267990 82412 267996
rect 88352 267918 88380 277780
rect 89548 272066 89576 277780
rect 89536 272060 89588 272066
rect 89536 272002 89588 272008
rect 90652 269793 90680 277780
rect 91848 272377 91876 277780
rect 91834 272368 91890 272377
rect 91834 272303 91890 272312
rect 93044 272202 93072 277780
rect 93032 272196 93084 272202
rect 93032 272138 93084 272144
rect 90638 269784 90694 269793
rect 90638 269719 90694 269728
rect 94240 269550 94268 277780
rect 94228 269544 94280 269550
rect 94228 269486 94280 269492
rect 88340 267912 88392 267918
rect 88340 267854 88392 267860
rect 95436 267850 95464 277780
rect 96632 269929 96660 277780
rect 97736 272785 97764 277780
rect 97722 272776 97778 272785
rect 97722 272711 97778 272720
rect 98932 272513 98960 277780
rect 100128 272649 100156 277780
rect 100114 272640 100170 272649
rect 100114 272575 100170 272584
rect 98918 272504 98974 272513
rect 98918 272439 98974 272448
rect 101324 270065 101352 277780
rect 101310 270056 101366 270065
rect 101310 269991 101366 270000
rect 96618 269920 96674 269929
rect 96618 269855 96674 269864
rect 102520 269686 102548 277780
rect 103716 270201 103744 277780
rect 104912 272134 104940 277780
rect 106016 272921 106044 277780
rect 107212 273057 107240 277780
rect 107198 273048 107254 273057
rect 107198 272983 107254 272992
rect 106002 272912 106058 272921
rect 106002 272847 106058 272856
rect 104900 272128 104952 272134
rect 104900 272070 104952 272076
rect 108408 270337 108436 277780
rect 108394 270328 108450 270337
rect 108394 270263 108450 270272
rect 103702 270192 103758 270201
rect 103702 270127 103758 270136
rect 109604 269754 109632 277780
rect 110800 269890 110828 277780
rect 111996 273193 112024 277780
rect 111982 273184 112038 273193
rect 111982 273119 112038 273128
rect 110788 269884 110840 269890
rect 110788 269826 110840 269832
rect 109592 269748 109644 269754
rect 109592 269690 109644 269696
rect 102508 269680 102560 269686
rect 102508 269622 102560 269628
rect 95424 267844 95476 267850
rect 95424 267786 95476 267792
rect 72976 266484 73028 266490
rect 72976 266426 73028 266432
rect 113192 266422 113220 277780
rect 114296 269822 114324 277780
rect 115492 271697 115520 277780
rect 115478 271688 115534 271697
rect 115478 271623 115534 271632
rect 114284 269816 114336 269822
rect 114284 269758 114336 269764
rect 116688 266558 116716 277780
rect 117884 272270 117912 277780
rect 117872 272264 117924 272270
rect 117872 272206 117924 272212
rect 119080 269958 119108 277780
rect 120276 271794 120304 277780
rect 120264 271788 120316 271794
rect 120264 271730 120316 271736
rect 121380 270473 121408 277780
rect 122576 271561 122604 277780
rect 122562 271552 122618 271561
rect 122562 271487 122618 271496
rect 121366 270464 121422 270473
rect 121366 270399 121422 270408
rect 119068 269952 119120 269958
rect 119068 269894 119120 269900
rect 123772 266626 123800 277780
rect 124968 272338 124996 277780
rect 124956 272332 125008 272338
rect 124956 272274 125008 272280
rect 126164 270026 126192 277780
rect 126152 270020 126204 270026
rect 126152 269962 126204 269968
rect 127360 268841 127388 277780
rect 128556 268977 128584 277780
rect 129660 272406 129688 277780
rect 129648 272400 129700 272406
rect 129648 272342 129700 272348
rect 130856 271726 130884 277780
rect 132052 272474 132080 277780
rect 132040 272468 132092 272474
rect 132040 272410 132092 272416
rect 130844 271720 130896 271726
rect 130844 271662 130896 271668
rect 133248 270162 133276 277780
rect 133236 270156 133288 270162
rect 133236 270098 133288 270104
rect 134444 270094 134472 277780
rect 135640 270230 135668 277780
rect 136836 272610 136864 277780
rect 136824 272604 136876 272610
rect 136824 272546 136876 272552
rect 137940 272542 137968 277780
rect 139136 272678 139164 277780
rect 139124 272672 139176 272678
rect 139124 272614 139176 272620
rect 137928 272536 137980 272542
rect 137928 272478 137980 272484
rect 140332 270366 140360 277780
rect 140320 270360 140372 270366
rect 140320 270302 140372 270308
rect 141528 270298 141556 277780
rect 141516 270292 141568 270298
rect 141516 270234 141568 270240
rect 135628 270224 135680 270230
rect 135628 270166 135680 270172
rect 134432 270088 134484 270094
rect 134432 270030 134484 270036
rect 128542 268968 128598 268977
rect 128542 268903 128598 268912
rect 127346 268832 127402 268841
rect 127346 268767 127402 268776
rect 142724 268705 142752 277780
rect 143920 272950 143948 277780
rect 143908 272944 143960 272950
rect 143908 272886 143960 272892
rect 145024 272746 145052 277780
rect 146220 272814 146248 277780
rect 146208 272808 146260 272814
rect 146208 272750 146260 272756
rect 145012 272740 145064 272746
rect 145012 272682 145064 272688
rect 147416 270434 147444 277780
rect 148612 272882 148640 277780
rect 149808 273086 149836 277780
rect 149796 273080 149848 273086
rect 149796 273022 149848 273028
rect 151004 273018 151032 277780
rect 150992 273012 151044 273018
rect 150992 272954 151044 272960
rect 148600 272876 148652 272882
rect 148600 272818 148652 272824
rect 147404 270428 147456 270434
rect 147404 270370 147456 270376
rect 152200 269074 152228 277780
rect 152188 269068 152240 269074
rect 152188 269010 152240 269016
rect 142710 268696 142766 268705
rect 142710 268631 142766 268640
rect 153304 268569 153332 277780
rect 154500 270502 154528 277780
rect 155696 273154 155724 277780
rect 155684 273148 155736 273154
rect 155684 273090 155736 273096
rect 156892 271794 156920 277780
rect 156788 271788 156840 271794
rect 156788 271730 156840 271736
rect 156880 271788 156932 271794
rect 156880 271730 156932 271736
rect 154488 270496 154540 270502
rect 154488 270438 154540 270444
rect 153290 268560 153346 268569
rect 156800 268530 156828 271730
rect 158088 271522 158116 277780
rect 158076 271516 158128 271522
rect 158076 271458 158128 271464
rect 159284 269006 159312 277780
rect 159272 269000 159324 269006
rect 159272 268942 159324 268948
rect 160480 268938 160508 277780
rect 160468 268932 160520 268938
rect 160468 268874 160520 268880
rect 161584 268870 161612 277780
rect 162780 271318 162808 277780
rect 163976 271658 164004 277780
rect 163964 271652 164016 271658
rect 163964 271594 164016 271600
rect 165172 271590 165200 277780
rect 165160 271584 165212 271590
rect 165160 271526 165212 271532
rect 162768 271312 162820 271318
rect 162768 271254 162820 271260
rect 161572 268864 161624 268870
rect 161572 268806 161624 268812
rect 166368 268802 166396 277780
rect 166356 268796 166408 268802
rect 166356 268738 166408 268744
rect 167564 268734 167592 277780
rect 167552 268728 167604 268734
rect 167552 268670 167604 268676
rect 168668 268598 168696 277780
rect 169864 271114 169892 277780
rect 171060 271454 171088 277780
rect 171048 271448 171100 271454
rect 171048 271390 171100 271396
rect 172256 271386 172284 277780
rect 172244 271380 172296 271386
rect 172244 271322 172296 271328
rect 169852 271108 169904 271114
rect 169852 271050 169904 271056
rect 173452 268666 173480 277780
rect 173440 268660 173492 268666
rect 173440 268602 173492 268608
rect 168656 268592 168708 268598
rect 168656 268534 168708 268540
rect 153290 268495 153346 268504
rect 156788 268524 156840 268530
rect 156788 268466 156840 268472
rect 174648 268462 174676 277780
rect 175844 270978 175872 277780
rect 176948 271046 176976 277780
rect 177856 273148 177908 273154
rect 177856 273090 177908 273096
rect 177868 271794 177896 273090
rect 178144 272066 178172 277780
rect 178040 272060 178092 272066
rect 178040 272002 178092 272008
rect 178132 272060 178184 272066
rect 178132 272002 178184 272008
rect 177856 271788 177908 271794
rect 177856 271730 177908 271736
rect 177948 271788 178000 271794
rect 177948 271730 178000 271736
rect 177960 271522 177988 271730
rect 177948 271516 178000 271522
rect 177948 271458 178000 271464
rect 178052 271250 178080 272002
rect 178132 271516 178184 271522
rect 178132 271458 178184 271464
rect 178144 271318 178172 271458
rect 178132 271312 178184 271318
rect 178132 271254 178184 271260
rect 178040 271244 178092 271250
rect 178040 271186 178092 271192
rect 179340 271182 179368 277780
rect 180064 271380 180116 271386
rect 180064 271322 180116 271328
rect 179328 271176 179380 271182
rect 179328 271118 179380 271124
rect 180076 271114 180104 271322
rect 180064 271108 180116 271114
rect 180064 271050 180116 271056
rect 176936 271040 176988 271046
rect 176936 270982 176988 270988
rect 175832 270972 175884 270978
rect 175832 270914 175884 270920
rect 179328 270972 179380 270978
rect 179328 270914 179380 270920
rect 174636 268456 174688 268462
rect 174636 268398 174688 268404
rect 179340 268394 179368 270914
rect 179328 268388 179380 268394
rect 179328 268330 179380 268336
rect 180536 268326 180564 277780
rect 180524 268320 180576 268326
rect 180524 268262 180576 268268
rect 181732 268258 181760 277780
rect 182928 271114 182956 277780
rect 182916 271108 182968 271114
rect 182916 271050 182968 271056
rect 181720 268252 181772 268258
rect 181720 268194 181772 268200
rect 184124 268122 184152 277780
rect 184940 272196 184992 272202
rect 184940 272138 184992 272144
rect 184952 268433 184980 272138
rect 185228 270978 185256 277780
rect 185216 270972 185268 270978
rect 185216 270914 185268 270920
rect 186424 270910 186452 277780
rect 186412 270904 186464 270910
rect 186412 270846 186464 270852
rect 187620 270774 187648 277780
rect 188816 272202 188844 277780
rect 188804 272196 188856 272202
rect 188804 272138 188856 272144
rect 188620 271244 188672 271250
rect 188620 271186 188672 271192
rect 187608 270768 187660 270774
rect 187608 270710 187660 270716
rect 188632 269618 188660 271186
rect 190012 270842 190040 277780
rect 190000 270836 190052 270842
rect 190000 270778 190052 270784
rect 191208 270706 191236 277780
rect 192116 271856 192168 271862
rect 192116 271798 192168 271804
rect 191196 270700 191248 270706
rect 191196 270642 191248 270648
rect 188620 269612 188672 269618
rect 188620 269554 188672 269560
rect 184938 268424 184994 268433
rect 184938 268359 184994 268368
rect 184112 268116 184164 268122
rect 184112 268058 184164 268064
rect 123760 266620 123812 266626
rect 123760 266562 123812 266568
rect 116676 266552 116728 266558
rect 116676 266494 116728 266500
rect 113180 266416 113232 266422
rect 113180 266358 113232 266364
rect 68192 266348 68244 266354
rect 68192 266290 68244 266296
rect 192128 264330 192156 271798
rect 192312 270570 192340 277780
rect 192484 271924 192536 271930
rect 192484 271866 192536 271872
rect 192300 270564 192352 270570
rect 192300 270506 192352 270512
rect 192496 264330 192524 271866
rect 193508 269142 193536 277780
rect 194138 271824 194194 271833
rect 194138 271759 194194 271768
rect 194506 271824 194562 271833
rect 194506 271759 194508 271768
rect 193496 269136 193548 269142
rect 193496 269078 193548 269084
rect 193678 269104 193734 269113
rect 193678 269039 193734 269048
rect 193220 266348 193272 266354
rect 193220 266290 193272 266296
rect 192128 264302 192418 264330
rect 192496 264302 192786 264330
rect 193232 264316 193260 266290
rect 193692 264316 193720 269039
rect 194152 264316 194180 271759
rect 194560 271759 194562 271768
rect 194508 271730 194560 271736
rect 194704 271726 194732 277780
rect 195428 271992 195480 271998
rect 195428 271934 195480 271940
rect 194692 271720 194744 271726
rect 194692 271662 194744 271668
rect 194600 269204 194652 269210
rect 194600 269146 194652 269152
rect 194612 264316 194640 269146
rect 195060 266484 195112 266490
rect 195060 266426 195112 266432
rect 195072 264316 195100 266426
rect 195440 264316 195468 271934
rect 195900 269498 195928 277780
rect 197110 277766 197400 277794
rect 197268 272060 197320 272066
rect 197268 272002 197320 272008
rect 196346 271960 196402 271969
rect 196346 271895 196402 271904
rect 195808 269470 195928 269498
rect 195808 269210 195836 269470
rect 195888 269408 195940 269414
rect 195888 269350 195940 269356
rect 195796 269204 195848 269210
rect 195796 269146 195848 269152
rect 195900 264316 195928 269350
rect 196360 264316 196388 271895
rect 197176 271856 197228 271862
rect 197176 271798 197228 271804
rect 196806 269240 196862 269249
rect 196806 269175 196862 269184
rect 196820 264316 196848 269175
rect 197188 267986 197216 271798
rect 197280 271250 197308 272002
rect 197268 271244 197320 271250
rect 197268 271186 197320 271192
rect 197372 269346 197400 277766
rect 198292 271862 198320 277780
rect 199106 272096 199162 272105
rect 199488 272066 199516 277780
rect 199934 272232 199990 272241
rect 199934 272167 199990 272176
rect 199106 272031 199162 272040
rect 199476 272060 199528 272066
rect 198280 271856 198332 271862
rect 198280 271798 198332 271804
rect 198648 270564 198700 270570
rect 198648 270506 198700 270512
rect 198660 269482 198688 270506
rect 199014 269512 199070 269521
rect 198648 269476 198700 269482
rect 199014 269447 199070 269456
rect 198648 269418 198700 269424
rect 197726 269376 197782 269385
rect 197268 269340 197320 269346
rect 197268 269282 197320 269288
rect 197360 269340 197412 269346
rect 197726 269311 197782 269320
rect 197360 269282 197412 269288
rect 197176 267980 197228 267986
rect 197176 267922 197228 267928
rect 197280 264316 197308 269282
rect 197740 264316 197768 269311
rect 198096 269272 198148 269278
rect 198096 269214 198148 269220
rect 198108 264316 198136 269214
rect 198556 268048 198608 268054
rect 198556 267990 198608 267996
rect 198568 264316 198596 267990
rect 199028 264316 199056 269447
rect 199120 264330 199148 272031
rect 199476 272002 199528 272008
rect 199120 264302 199502 264330
rect 199948 264316 199976 272167
rect 200394 269648 200450 269657
rect 200394 269583 200450 269592
rect 200408 264316 200436 269583
rect 200592 269278 200620 277780
rect 201314 272776 201370 272785
rect 201314 272711 201370 272720
rect 200764 269612 200816 269618
rect 200764 269554 200816 269560
rect 200580 269272 200632 269278
rect 200580 269214 200632 269220
rect 200776 264316 200804 269554
rect 201328 268054 201356 272711
rect 201788 271998 201816 277780
rect 202142 272368 202198 272377
rect 202142 272303 202198 272312
rect 201776 271992 201828 271998
rect 201776 271934 201828 271940
rect 201682 269784 201738 269793
rect 201682 269719 201738 269728
rect 201316 268048 201368 268054
rect 201316 267990 201368 267996
rect 201224 267912 201276 267918
rect 201224 267854 201276 267860
rect 201236 264316 201264 267854
rect 201696 264316 201724 269719
rect 202156 264316 202184 272303
rect 202696 272128 202748 272134
rect 202696 272070 202748 272076
rect 202604 269544 202656 269550
rect 202604 269486 202656 269492
rect 202616 264316 202644 269486
rect 202708 267782 202736 272070
rect 202788 270768 202840 270774
rect 202788 270710 202840 270716
rect 202800 270570 202828 270710
rect 202788 270564 202840 270570
rect 202788 270506 202840 270512
rect 202984 269550 203012 277780
rect 203522 273048 203578 273057
rect 203522 272983 203578 272992
rect 202972 269544 203024 269550
rect 202972 269486 203024 269492
rect 203062 268424 203118 268433
rect 203062 268359 203118 268368
rect 202696 267776 202748 267782
rect 202696 267718 202748 267724
rect 203076 264316 203104 268359
rect 203536 268161 203564 272983
rect 204180 269414 204208 277780
rect 204810 272504 204866 272513
rect 204810 272439 204866 272448
rect 204350 269920 204406 269929
rect 204350 269855 204406 269864
rect 204168 269408 204220 269414
rect 204168 269350 204220 269356
rect 203522 268152 203578 268161
rect 203522 268087 203578 268096
rect 203892 268048 203944 268054
rect 203892 267990 203944 267996
rect 203524 267844 203576 267850
rect 203524 267786 203576 267792
rect 203536 264316 203564 267786
rect 203904 264316 203932 267990
rect 204364 264316 204392 269855
rect 204824 264316 204852 272439
rect 205376 272134 205404 277780
rect 205730 272640 205786 272649
rect 205730 272575 205786 272584
rect 205548 272264 205600 272270
rect 205548 272206 205600 272212
rect 205364 272128 205416 272134
rect 205364 272070 205416 272076
rect 205270 270056 205326 270065
rect 205270 269991 205326 270000
rect 205284 264316 205312 269991
rect 205560 267850 205588 272206
rect 205548 267844 205600 267850
rect 205548 267786 205600 267792
rect 205744 264316 205772 272575
rect 206468 270496 206520 270502
rect 206468 270438 206520 270444
rect 206192 269680 206244 269686
rect 206192 269622 206244 269628
rect 206204 264316 206232 269622
rect 206480 268054 206508 270438
rect 206572 268190 206600 277780
rect 207478 272912 207534 272921
rect 207478 272847 207534 272856
rect 206744 270768 206796 270774
rect 206744 270710 206796 270716
rect 206756 270638 206784 270710
rect 206744 270632 206796 270638
rect 206744 270574 206796 270580
rect 207018 270192 207074 270201
rect 207018 270127 207074 270136
rect 206560 268184 206612 268190
rect 206560 268126 206612 268132
rect 206468 268048 206520 268054
rect 206468 267990 206520 267996
rect 206560 267776 206612 267782
rect 206560 267718 206612 267724
rect 206572 264316 206600 267718
rect 207032 264316 207060 270127
rect 207492 264316 207520 272847
rect 207768 269618 207796 277780
rect 208886 277766 209176 277794
rect 208490 271824 208546 271833
rect 208490 271759 208546 271768
rect 208504 271726 208532 271759
rect 208492 271720 208544 271726
rect 208492 271662 208544 271668
rect 208032 270360 208084 270366
rect 207938 270328 207994 270337
rect 208308 270360 208360 270366
rect 208084 270308 208308 270314
rect 208032 270302 208360 270308
rect 208044 270286 208348 270302
rect 207938 270263 207994 270272
rect 207756 269612 207808 269618
rect 207756 269554 207808 269560
rect 207952 264316 207980 270263
rect 208400 270224 208452 270230
rect 208228 270184 208400 270212
rect 208228 270094 208256 270184
rect 208400 270166 208452 270172
rect 208216 270088 208268 270094
rect 208216 270030 208268 270036
rect 208860 269748 208912 269754
rect 208860 269690 208912 269696
rect 208398 268152 208454 268161
rect 208398 268087 208454 268096
rect 208412 264316 208440 268087
rect 208872 264316 208900 269690
rect 209148 269686 209176 277766
rect 209226 273184 209282 273193
rect 209226 273119 209282 273128
rect 209136 269680 209188 269686
rect 209136 269622 209188 269628
rect 209240 264316 209268 273119
rect 210068 269890 210096 277780
rect 210606 271688 210662 271697
rect 210606 271623 210662 271632
rect 209688 269884 209740 269890
rect 209688 269826 209740 269832
rect 210056 269884 210108 269890
rect 210056 269826 210108 269832
rect 209700 264316 209728 269826
rect 210148 266416 210200 266422
rect 210148 266358 210200 266364
rect 210160 264316 210188 266358
rect 210620 264316 210648 271623
rect 211068 269816 211120 269822
rect 211068 269758 211120 269764
rect 211080 264316 211108 269758
rect 211264 267918 211292 277780
rect 211896 269952 211948 269958
rect 211896 269894 211948 269900
rect 211252 267912 211304 267918
rect 211252 267854 211304 267860
rect 211528 266552 211580 266558
rect 211528 266494 211580 266500
rect 211540 264316 211568 266494
rect 211908 264316 211936 269894
rect 212460 269754 212488 277780
rect 213274 271552 213330 271561
rect 213274 271487 213330 271496
rect 212448 269748 212500 269754
rect 212448 269690 212500 269696
rect 212816 268524 212868 268530
rect 212816 268466 212868 268472
rect 212356 267844 212408 267850
rect 212356 267786 212408 267792
rect 212368 264316 212396 267786
rect 212828 264316 212856 268466
rect 213288 264316 213316 271487
rect 213656 270026 213684 277780
rect 213734 270464 213790 270473
rect 213734 270399 213790 270408
rect 213644 270020 213696 270026
rect 213644 269962 213696 269968
rect 213748 264316 213776 270399
rect 214656 269952 214708 269958
rect 214656 269894 214708 269900
rect 214196 266620 214248 266626
rect 214196 266562 214248 266568
rect 214208 264316 214236 266562
rect 214668 264316 214696 269894
rect 214852 269822 214880 277780
rect 215668 272400 215720 272406
rect 215668 272342 215720 272348
rect 215024 272332 215076 272338
rect 215024 272274 215076 272280
rect 214840 269816 214892 269822
rect 214840 269758 214892 269764
rect 215036 264316 215064 272274
rect 215482 268832 215538 268841
rect 215482 268767 215538 268776
rect 215496 264316 215524 268767
rect 215680 264330 215708 272342
rect 215956 270162 215984 277780
rect 215944 270156 215996 270162
rect 215944 270098 215996 270104
rect 217152 269958 217180 277780
rect 217692 272468 217744 272474
rect 217692 272410 217744 272416
rect 217324 270088 217376 270094
rect 217324 270030 217376 270036
rect 217140 269952 217192 269958
rect 217140 269894 217192 269900
rect 216402 268968 216458 268977
rect 216402 268903 216458 268912
rect 215680 264302 215970 264330
rect 216416 264316 216444 268903
rect 216864 267980 216916 267986
rect 216864 267922 216916 267928
rect 216876 264316 216904 267922
rect 217336 264316 217364 270030
rect 217704 264316 217732 272410
rect 218348 270230 218376 277780
rect 218612 272604 218664 272610
rect 218612 272546 218664 272552
rect 218152 270224 218204 270230
rect 218152 270166 218204 270172
rect 218336 270224 218388 270230
rect 218336 270166 218388 270172
rect 218164 264316 218192 270166
rect 218624 264316 218652 272546
rect 219440 272536 219492 272542
rect 219440 272478 219492 272484
rect 219072 270292 219124 270298
rect 219072 270234 219124 270240
rect 219084 264316 219112 270234
rect 219452 264330 219480 272478
rect 219544 268530 219572 277780
rect 220360 272672 220412 272678
rect 220360 272614 220412 272620
rect 219992 270360 220044 270366
rect 219992 270302 220044 270308
rect 219532 268524 219584 268530
rect 219532 268466 219584 268472
rect 219452 264302 219558 264330
rect 220004 264316 220032 270302
rect 220372 264316 220400 272614
rect 220740 270366 220768 277780
rect 221280 272944 221332 272950
rect 221280 272886 221332 272892
rect 220820 270428 220872 270434
rect 220820 270370 220872 270376
rect 220728 270360 220780 270366
rect 220728 270302 220780 270308
rect 220832 264316 220860 270370
rect 221292 264316 221320 272886
rect 221936 270298 221964 277780
rect 223028 272808 223080 272814
rect 223028 272750 223080 272756
rect 222200 272740 222252 272746
rect 222200 272682 222252 272688
rect 221924 270292 221976 270298
rect 221924 270234 221976 270240
rect 221738 268696 221794 268705
rect 221738 268631 221794 268640
rect 221752 264316 221780 268631
rect 222212 264316 222240 272682
rect 222660 270496 222712 270502
rect 222660 270438 222712 270444
rect 222672 264316 222700 270438
rect 223040 264316 223068 272750
rect 223132 270094 223160 277780
rect 223948 273012 224000 273018
rect 223948 272954 224000 272960
rect 223212 272876 223264 272882
rect 223212 272818 223264 272824
rect 223120 270088 223172 270094
rect 223120 270030 223172 270036
rect 223224 264330 223252 272818
rect 223224 264302 223514 264330
rect 223960 264316 223988 272954
rect 224236 270434 224264 277780
rect 224408 273080 224460 273086
rect 224408 273022 224460 273028
rect 224224 270428 224276 270434
rect 224224 270370 224276 270376
rect 224420 264316 224448 273022
rect 225432 270502 225460 277780
rect 225880 273216 225932 273222
rect 225880 273158 225932 273164
rect 225420 270496 225472 270502
rect 225420 270438 225472 270444
rect 224868 269068 224920 269074
rect 224868 269010 224920 269016
rect 224880 264316 224908 269010
rect 225786 268560 225842 268569
rect 225786 268495 225842 268504
rect 225328 268048 225380 268054
rect 225328 267990 225380 267996
rect 225340 264316 225368 267990
rect 225800 264316 225828 268495
rect 225892 264330 225920 273158
rect 226524 271788 226576 271794
rect 226524 271730 226576 271736
rect 226432 271040 226484 271046
rect 226432 270982 226484 270988
rect 226444 269550 226472 270982
rect 226340 269544 226392 269550
rect 226340 269486 226392 269492
rect 226432 269544 226484 269550
rect 226432 269486 226484 269492
rect 226352 269074 226380 269486
rect 226340 269068 226392 269074
rect 226340 269010 226392 269016
rect 226536 264330 226564 271730
rect 226628 271046 226656 277780
rect 227076 272264 227128 272270
rect 227076 272206 227128 272212
rect 226616 271040 226668 271046
rect 226616 270982 226668 270988
rect 225892 264302 226182 264330
rect 226536 264302 226642 264330
rect 227088 264316 227116 272206
rect 227824 270570 227852 277780
rect 228824 271516 228876 271522
rect 228824 271458 228876 271464
rect 227812 270564 227864 270570
rect 227812 270506 227864 270512
rect 227536 269000 227588 269006
rect 227536 268942 227588 268948
rect 227548 264316 227576 268942
rect 228456 268932 228508 268938
rect 228456 268874 228508 268880
rect 227996 268864 228048 268870
rect 227996 268806 228048 268812
rect 228008 264316 228036 268806
rect 228468 264316 228496 268874
rect 228836 264316 228864 271458
rect 229020 270638 229048 277780
rect 230216 272474 230244 277780
rect 230204 272468 230256 272474
rect 230204 272410 230256 272416
rect 229744 271652 229796 271658
rect 229744 271594 229796 271600
rect 229468 271584 229520 271590
rect 229468 271526 229520 271532
rect 229376 270768 229428 270774
rect 229376 270710 229428 270716
rect 229008 270632 229060 270638
rect 229008 270574 229060 270580
rect 229388 268870 229416 270710
rect 229376 268864 229428 268870
rect 229376 268806 229428 268812
rect 229480 264330 229508 271526
rect 229310 264302 229508 264330
rect 229756 264316 229784 271594
rect 231412 271522 231440 277780
rect 232516 272610 232544 277780
rect 232504 272604 232556 272610
rect 232504 272546 232556 272552
rect 233712 271658 233740 277780
rect 234908 272814 234936 277780
rect 236104 272882 236132 277780
rect 236092 272876 236144 272882
rect 236092 272818 236144 272824
rect 234896 272808 234948 272814
rect 234896 272750 234948 272756
rect 237300 272746 237328 277780
rect 237288 272740 237340 272746
rect 237288 272682 237340 272688
rect 238496 272202 238524 277780
rect 239600 272950 239628 277780
rect 239588 272944 239640 272950
rect 239588 272886 239640 272892
rect 234804 272196 234856 272202
rect 234804 272138 234856 272144
rect 238484 272196 238536 272202
rect 238484 272138 238536 272144
rect 233700 271652 233752 271658
rect 233700 271594 233752 271600
rect 231400 271516 231452 271522
rect 231400 271458 231452 271464
rect 232412 271448 232464 271454
rect 232412 271390 232464 271396
rect 231492 271380 231544 271386
rect 231492 271322 231544 271328
rect 230204 270700 230256 270706
rect 230204 270642 230256 270648
rect 230216 268938 230244 270642
rect 230204 268932 230256 268938
rect 230204 268874 230256 268880
rect 230204 268796 230256 268802
rect 230204 268738 230256 268744
rect 230216 264316 230244 268738
rect 231124 268728 231176 268734
rect 231124 268670 231176 268676
rect 230664 268592 230716 268598
rect 230664 268534 230716 268540
rect 230676 264316 230704 268534
rect 231136 264316 231164 268670
rect 231504 264316 231532 271322
rect 231768 271312 231820 271318
rect 231768 271254 231820 271260
rect 231780 270484 231808 271254
rect 231952 271244 232004 271250
rect 231952 271186 232004 271192
rect 231780 270456 231900 270484
rect 231872 264330 231900 270456
rect 231964 268054 231992 271186
rect 232044 271108 232096 271114
rect 232044 271050 232096 271056
rect 231952 268048 232004 268054
rect 231952 267990 232004 267996
rect 232056 267986 232084 271050
rect 232136 270904 232188 270910
rect 232136 270846 232188 270852
rect 232148 269006 232176 270846
rect 232136 269000 232188 269006
rect 232136 268942 232188 268948
rect 232044 267980 232096 267986
rect 232044 267922 232096 267928
rect 231872 264302 231978 264330
rect 232424 264316 232452 271390
rect 234528 271176 234580 271182
rect 234528 271118 234580 271124
rect 232504 270836 232556 270842
rect 232504 270778 232556 270784
rect 232516 267782 232544 270778
rect 234540 270484 234568 271118
rect 234712 270972 234764 270978
rect 234712 270914 234764 270920
rect 234540 270456 234660 270484
rect 234160 269544 234212 269550
rect 234160 269486 234212 269492
rect 232872 268660 232924 268666
rect 232872 268602 232924 268608
rect 232504 267776 232556 267782
rect 232504 267718 232556 267724
rect 232884 264316 232912 268602
rect 233792 268456 233844 268462
rect 233792 268398 233844 268404
rect 233332 268388 233384 268394
rect 233332 268330 233384 268336
rect 233344 264316 233372 268330
rect 233804 264316 233832 268398
rect 234172 264316 234200 269486
rect 234632 264316 234660 270456
rect 234724 267850 234752 270914
rect 234816 268462 234844 272138
rect 240140 272128 240192 272134
rect 240140 272070 240192 272076
rect 239956 269476 240008 269482
rect 239956 269418 240008 269424
rect 237288 269000 237340 269006
rect 237288 268942 237340 268948
rect 234804 268456 234856 268462
rect 234804 268398 234856 268404
rect 235540 268320 235592 268326
rect 235540 268262 235592 268268
rect 235080 268048 235132 268054
rect 235080 267990 235132 267996
rect 234712 267844 234764 267850
rect 234712 267786 234764 267792
rect 235092 264316 235120 267990
rect 235552 264316 235580 268262
rect 236460 268252 236512 268258
rect 236460 268194 236512 268200
rect 235724 267980 235776 267986
rect 235724 267922 235776 267928
rect 235736 264330 235764 267922
rect 235736 264302 236026 264330
rect 236472 264316 236500 268194
rect 236920 268116 236972 268122
rect 236920 268058 236972 268064
rect 236932 264316 236960 268058
rect 237300 264316 237328 268942
rect 238208 268932 238260 268938
rect 238208 268874 238260 268880
rect 237748 267844 237800 267850
rect 237748 267786 237800 267792
rect 237760 264316 237788 267786
rect 238220 264316 238248 268874
rect 239588 268864 239640 268870
rect 239588 268806 239640 268812
rect 239128 268456 239180 268462
rect 239128 268398 239180 268404
rect 238668 267776 238720 267782
rect 238668 267718 238720 267724
rect 238680 264316 238708 267718
rect 239140 264316 239168 268398
rect 239600 264316 239628 268806
rect 239968 264316 239996 269418
rect 240152 268598 240180 272070
rect 240796 271726 240824 277780
rect 240876 271856 240928 271862
rect 240876 271798 240928 271804
rect 240784 271720 240836 271726
rect 240784 271662 240836 271668
rect 240416 269136 240468 269142
rect 240416 269078 240468 269084
rect 240140 268592 240192 268598
rect 240140 268534 240192 268540
rect 240428 264316 240456 269078
rect 240888 264316 240916 271798
rect 241992 271794 242020 277780
rect 243188 273086 243216 277780
rect 243176 273080 243228 273086
rect 243176 273022 243228 273028
rect 242624 272060 242676 272066
rect 242624 272002 242676 272008
rect 242256 271924 242308 271930
rect 242256 271866 242308 271872
rect 241980 271788 242032 271794
rect 241980 271730 242032 271736
rect 241796 269340 241848 269346
rect 241796 269282 241848 269288
rect 241336 269204 241388 269210
rect 241336 269146 241388 269152
rect 241348 264316 241376 269146
rect 241808 264316 241836 269282
rect 242268 264316 242296 271866
rect 242636 264316 242664 272002
rect 243544 271992 243596 271998
rect 243544 271934 243596 271940
rect 243084 269272 243136 269278
rect 243084 269214 243136 269220
rect 243096 264316 243124 269214
rect 243556 264316 243584 271934
rect 244384 271862 244412 277780
rect 244372 271856 244424 271862
rect 244372 271798 244424 271804
rect 245580 271590 245608 277780
rect 246776 271726 246804 277780
rect 246764 271720 246816 271726
rect 246764 271662 246816 271668
rect 247880 271658 247908 277780
rect 247868 271652 247920 271658
rect 247868 271594 247920 271600
rect 245568 271584 245620 271590
rect 245568 271526 245620 271532
rect 249076 271182 249104 277780
rect 250272 271590 250300 277780
rect 250168 271584 250220 271590
rect 250168 271526 250220 271532
rect 250260 271584 250312 271590
rect 250260 271526 250312 271532
rect 249064 271176 249116 271182
rect 249064 271118 249116 271124
rect 250180 270978 250208 271526
rect 251468 271250 251496 277780
rect 251456 271244 251508 271250
rect 251456 271186 251508 271192
rect 250168 270972 250220 270978
rect 250168 270914 250220 270920
rect 252664 270706 252692 277780
rect 253860 271114 253888 277780
rect 254216 272468 254268 272474
rect 254216 272410 254268 272416
rect 253848 271108 253900 271114
rect 253848 271050 253900 271056
rect 252928 271040 252980 271046
rect 252928 270982 252980 270988
rect 252652 270700 252704 270706
rect 252652 270642 252704 270648
rect 252468 270496 252520 270502
rect 252468 270438 252520 270444
rect 252008 270428 252060 270434
rect 252008 270370 252060 270376
rect 250720 270360 250772 270366
rect 250720 270302 250772 270308
rect 249800 270224 249852 270230
rect 249800 270166 249852 270172
rect 248880 270156 248932 270162
rect 248880 270098 248932 270104
rect 248052 270020 248104 270026
rect 248052 269962 248104 269968
rect 246672 269884 246724 269890
rect 246672 269826 246724 269832
rect 246212 269680 246264 269686
rect 246212 269622 246264 269628
rect 245752 269612 245804 269618
rect 245752 269554 245804 269560
rect 244464 269408 244516 269414
rect 244464 269350 244516 269356
rect 244004 269068 244056 269074
rect 244004 269010 244056 269016
rect 244016 264316 244044 269010
rect 244476 264316 244504 269350
rect 244924 268592 244976 268598
rect 244924 268534 244976 268540
rect 244936 264316 244964 268534
rect 245292 268184 245344 268190
rect 245292 268126 245344 268132
rect 245304 264316 245332 268126
rect 245764 264316 245792 269554
rect 246224 264316 246252 269622
rect 246684 264316 246712 269826
rect 247592 269748 247644 269754
rect 247592 269690 247644 269696
rect 247132 267912 247184 267918
rect 247132 267854 247184 267860
rect 247144 264316 247172 267854
rect 247604 264316 247632 269690
rect 248064 264316 248092 269962
rect 248420 269816 248472 269822
rect 248420 269758 248472 269764
rect 248432 264316 248460 269758
rect 248892 264316 248920 270098
rect 249340 269952 249392 269958
rect 249340 269894 249392 269900
rect 249352 264316 249380 269894
rect 249812 264316 249840 270166
rect 250260 268660 250312 268666
rect 250260 268602 250312 268608
rect 250272 264316 250300 268602
rect 250732 264316 250760 270302
rect 251088 270292 251140 270298
rect 251088 270234 251140 270240
rect 251100 264316 251128 270234
rect 251548 270088 251600 270094
rect 251548 270030 251600 270036
rect 251560 264316 251588 270030
rect 252020 264316 252048 270370
rect 252480 264316 252508 270438
rect 252940 264316 252968 270982
rect 253756 270632 253808 270638
rect 253756 270574 253808 270580
rect 253388 270564 253440 270570
rect 253388 270506 253440 270512
rect 253400 264316 253428 270506
rect 253768 264316 253796 270574
rect 254228 264316 254256 272410
rect 255056 271522 255084 277780
rect 256056 272808 256108 272814
rect 256056 272750 256108 272756
rect 255136 272604 255188 272610
rect 255136 272546 255188 272552
rect 254676 271516 254728 271522
rect 254676 271458 254728 271464
rect 255044 271516 255096 271522
rect 255044 271458 255096 271464
rect 254688 264316 254716 271458
rect 255148 264316 255176 272546
rect 255596 271788 255648 271794
rect 255596 271730 255648 271736
rect 255608 264316 255636 271730
rect 256068 264316 256096 272750
rect 256160 271318 256188 277780
rect 256424 272876 256476 272882
rect 256424 272818 256476 272824
rect 256148 271312 256200 271318
rect 256148 271254 256200 271260
rect 256436 264316 256464 272818
rect 257160 272740 257212 272746
rect 257160 272682 257212 272688
rect 257172 264330 257200 272682
rect 257252 272196 257304 272202
rect 257252 272138 257304 272144
rect 257264 271266 257292 272138
rect 257356 271386 257384 277780
rect 257804 272944 257856 272950
rect 257804 272886 257856 272892
rect 257344 271380 257396 271386
rect 257344 271322 257396 271328
rect 257264 271238 257384 271266
rect 256910 264302 257200 264330
rect 257356 264316 257384 271238
rect 257816 264316 257844 272886
rect 258264 271856 258316 271862
rect 258264 271798 258316 271804
rect 258276 264316 258304 271798
rect 258552 271454 258580 277780
rect 259184 273080 259236 273086
rect 259184 273022 259236 273028
rect 258724 271924 258776 271930
rect 258724 271866 258776 271872
rect 258540 271448 258592 271454
rect 258540 271390 258592 271396
rect 258736 264316 258764 271866
rect 259196 264316 259224 273022
rect 259552 271992 259604 271998
rect 259552 271934 259604 271940
rect 259564 264316 259592 271934
rect 259748 270842 259776 277780
rect 260944 273086 260972 277780
rect 260932 273080 260984 273086
rect 260932 273022 260984 273028
rect 262140 271794 262168 277780
rect 263244 273222 263272 277780
rect 263232 273216 263284 273222
rect 263232 273158 263284 273164
rect 264440 273154 264468 277780
rect 264428 273148 264480 273154
rect 264428 273090 264480 273096
rect 262128 271788 262180 271794
rect 262128 271730 262180 271736
rect 260472 271720 260524 271726
rect 260472 271662 260524 271668
rect 260012 270972 260064 270978
rect 260012 270914 260064 270920
rect 259736 270836 259788 270842
rect 259736 270778 259788 270784
rect 260024 264316 260052 270914
rect 260484 264316 260512 271662
rect 260932 271652 260984 271658
rect 260932 271594 260984 271600
rect 260944 264316 260972 271594
rect 261852 271584 261904 271590
rect 261852 271526 261904 271532
rect 261392 271176 261444 271182
rect 261392 271118 261444 271124
rect 261404 264316 261432 271118
rect 261864 264316 261892 271526
rect 263600 271516 263652 271522
rect 263600 271458 263652 271464
rect 262220 271244 262272 271250
rect 262220 271186 262272 271192
rect 262232 264316 262260 271186
rect 263140 271108 263192 271114
rect 263140 271050 263192 271056
rect 262864 270700 262916 270706
rect 262864 270642 262916 270648
rect 262876 264330 262904 270642
rect 262706 264302 262904 264330
rect 263152 264316 263180 271050
rect 263612 264316 263640 271458
rect 264888 271448 264940 271454
rect 264888 271390 264940 271396
rect 264520 271380 264572 271386
rect 264520 271322 264572 271328
rect 264060 271312 264112 271318
rect 264060 271254 264112 271260
rect 264072 264316 264100 271254
rect 264532 264316 264560 271322
rect 264900 264316 264928 271390
rect 265348 270836 265400 270842
rect 265348 270778 265400 270784
rect 265360 264316 265388 270778
rect 265636 270502 265664 277780
rect 266728 273216 266780 273222
rect 266728 273158 266780 273164
rect 265808 273080 265860 273086
rect 265808 273022 265860 273028
rect 265624 270496 265676 270502
rect 265624 270438 265676 270444
rect 265820 264316 265848 273022
rect 266268 271788 266320 271794
rect 266268 271730 266320 271736
rect 266280 264316 266308 271730
rect 266740 264316 266768 273158
rect 266832 271114 266860 277780
rect 268042 277766 268516 277794
rect 267188 273148 267240 273154
rect 267188 273090 267240 273096
rect 266820 271108 266872 271114
rect 266820 271050 266872 271056
rect 267200 264316 267228 273090
rect 268016 271108 268068 271114
rect 268016 271050 268068 271056
rect 267556 270496 267608 270502
rect 267556 270438 267608 270444
rect 267568 264316 267596 270438
rect 268028 264316 268056 271050
rect 268488 264316 268516 277766
rect 268948 277766 269238 277794
rect 268948 264316 268976 277766
rect 269856 270496 269908 270502
rect 269856 270438 269908 270444
rect 269396 269000 269448 269006
rect 269396 268942 269448 268948
rect 269408 264316 269436 268942
rect 269868 264316 269896 270438
rect 270316 270428 270368 270434
rect 270316 270370 270368 270376
rect 270328 264316 270356 270370
rect 270420 269006 270448 277780
rect 271524 270502 271552 277780
rect 271512 270496 271564 270502
rect 271512 270438 271564 270444
rect 272064 270496 272116 270502
rect 272064 270438 272116 270444
rect 270684 270360 270736 270366
rect 270684 270302 270736 270308
rect 270408 269000 270460 269006
rect 270408 268942 270460 268948
rect 270696 264316 270724 270302
rect 271144 270292 271196 270298
rect 271144 270234 271196 270240
rect 271156 264316 271184 270234
rect 271604 270088 271656 270094
rect 271604 270030 271656 270036
rect 271616 264316 271644 270030
rect 272076 264316 272104 270438
rect 272720 270434 272748 277780
rect 272708 270428 272760 270434
rect 272708 270370 272760 270376
rect 272984 270428 273036 270434
rect 272984 270370 273036 270376
rect 272524 270224 272576 270230
rect 272524 270166 272576 270172
rect 272536 264316 272564 270166
rect 272996 264316 273024 270370
rect 273916 270366 273944 277780
rect 273904 270360 273956 270366
rect 273904 270302 273956 270308
rect 274272 270360 274324 270366
rect 274272 270302 274324 270308
rect 273720 270156 273772 270162
rect 273720 270098 273772 270104
rect 273732 264330 273760 270098
rect 273812 268728 273864 268734
rect 273812 268670 273864 268676
rect 273378 264302 273760 264330
rect 273824 264316 273852 268670
rect 274284 264316 274312 270302
rect 275112 270298 275140 277780
rect 275100 270292 275152 270298
rect 275100 270234 275152 270240
rect 276308 270094 276336 277780
rect 277504 270502 277532 277780
rect 277492 270496 277544 270502
rect 277492 270438 277544 270444
rect 277400 270292 277452 270298
rect 277400 270234 277452 270240
rect 276296 270088 276348 270094
rect 276296 270030 276348 270036
rect 276940 269952 276992 269958
rect 276940 269894 276992 269900
rect 276480 268456 276532 268462
rect 276480 268398 276532 268404
rect 275192 268388 275244 268394
rect 275192 268330 275244 268336
rect 274732 268320 274784 268326
rect 274732 268262 274784 268268
rect 274744 264316 274772 268262
rect 275204 264316 275232 268330
rect 275652 268252 275704 268258
rect 275652 268194 275704 268200
rect 275664 264316 275692 268194
rect 276296 267912 276348 267918
rect 276296 267854 276348 267860
rect 276308 264330 276336 267854
rect 276046 264302 276336 264330
rect 276492 264316 276520 268398
rect 276952 264316 276980 269894
rect 277412 264316 277440 270234
rect 278700 270230 278728 277780
rect 279804 270434 279832 277780
rect 279792 270428 279844 270434
rect 279792 270370 279844 270376
rect 278688 270224 278740 270230
rect 278688 270166 278740 270172
rect 278780 270224 278832 270230
rect 278780 270166 278832 270172
rect 278688 270088 278740 270094
rect 278688 270030 278740 270036
rect 278320 270020 278372 270026
rect 278320 269962 278372 269968
rect 277860 269680 277912 269686
rect 277860 269622 277912 269628
rect 277872 264316 277900 269622
rect 278332 264316 278360 269962
rect 278700 264316 278728 270030
rect 278792 269958 278820 270166
rect 281000 270162 281028 277780
rect 280988 270156 281040 270162
rect 280988 270098 281040 270104
rect 281540 270020 281592 270026
rect 281540 269962 281592 269968
rect 278780 269952 278832 269958
rect 278780 269894 278832 269900
rect 279608 269952 279660 269958
rect 279608 269894 279660 269900
rect 279148 269884 279200 269890
rect 279148 269826 279200 269832
rect 279160 264316 279188 269826
rect 279620 264316 279648 269894
rect 280528 269816 280580 269822
rect 280528 269758 280580 269764
rect 280068 269748 280120 269754
rect 280068 269690 280120 269696
rect 280080 264316 280108 269690
rect 280540 264316 280568 269758
rect 281552 269686 281580 269962
rect 281540 269680 281592 269686
rect 281540 269622 281592 269628
rect 281816 269680 281868 269686
rect 281816 269622 281868 269628
rect 281448 269612 281500 269618
rect 281448 269554 281500 269560
rect 280988 269544 281040 269550
rect 280988 269486 281040 269492
rect 281000 264316 281028 269486
rect 281460 264316 281488 269554
rect 281828 264316 281856 269622
rect 282196 268734 282224 277780
rect 283392 270366 283420 277780
rect 284208 272060 284260 272066
rect 284208 272002 284260 272008
rect 283380 270360 283432 270366
rect 283380 270302 283432 270308
rect 282736 269476 282788 269482
rect 282736 269418 282788 269424
rect 282276 269408 282328 269414
rect 282276 269350 282328 269356
rect 282184 268728 282236 268734
rect 282184 268670 282236 268676
rect 282288 264316 282316 269350
rect 282748 264316 282776 269418
rect 283656 269340 283708 269346
rect 283656 269282 283708 269288
rect 283196 269272 283248 269278
rect 283196 269214 283248 269220
rect 283208 264316 283236 269214
rect 283668 264316 283696 269282
rect 284220 264330 284248 272002
rect 284484 269136 284536 269142
rect 284484 269078 284536 269084
rect 284142 264302 284248 264330
rect 284496 264316 284524 269078
rect 284588 268326 284616 277780
rect 285404 271992 285456 271998
rect 285404 271934 285456 271940
rect 284944 269204 284996 269210
rect 284944 269146 284996 269152
rect 284576 268320 284628 268326
rect 284576 268262 284628 268268
rect 284956 264316 284984 269146
rect 285416 264316 285444 271934
rect 285784 268394 285812 277780
rect 286784 271312 286836 271318
rect 286784 271254 286836 271260
rect 286692 271108 286744 271114
rect 286692 271050 286744 271056
rect 285864 270972 285916 270978
rect 285864 270914 285916 270920
rect 285772 268388 285824 268394
rect 285772 268330 285824 268336
rect 285876 264316 285904 270914
rect 286704 264330 286732 271050
rect 286350 264302 286732 264330
rect 286796 264316 286824 271254
rect 286888 268258 286916 277780
rect 287612 271380 287664 271386
rect 287612 271322 287664 271328
rect 287152 271176 287204 271182
rect 287152 271118 287204 271124
rect 286876 268252 286928 268258
rect 286876 268194 286928 268200
rect 287164 264316 287192 271118
rect 287624 264316 287652 271322
rect 288084 267918 288112 277780
rect 288532 271448 288584 271454
rect 288532 271390 288584 271396
rect 288164 271244 288216 271250
rect 288164 271186 288216 271192
rect 288072 267912 288124 267918
rect 288072 267854 288124 267860
rect 288176 264330 288204 271186
rect 288098 264302 288204 264330
rect 288544 264316 288572 271390
rect 289280 268462 289308 277780
rect 290280 271924 290332 271930
rect 290280 271866 290332 271872
rect 289544 271856 289596 271862
rect 289544 271798 289596 271804
rect 289360 271516 289412 271522
rect 289360 271458 289412 271464
rect 289268 268456 289320 268462
rect 289268 268398 289320 268404
rect 289372 264330 289400 271458
rect 289556 264330 289584 271798
rect 289820 271652 289872 271658
rect 289820 271594 289872 271600
rect 289018 264302 289400 264330
rect 289478 264302 289584 264330
rect 289832 264316 289860 271594
rect 290292 264316 290320 271866
rect 290476 270230 290504 277780
rect 290740 271720 290792 271726
rect 290740 271662 290792 271668
rect 290464 270224 290516 270230
rect 290464 270166 290516 270172
rect 290752 264316 290780 271662
rect 291200 271584 291252 271590
rect 291200 271526 291252 271532
rect 291212 264316 291240 271526
rect 291672 270298 291700 277780
rect 292120 273216 292172 273222
rect 292120 273158 292172 273164
rect 291752 271788 291804 271794
rect 291752 271730 291804 271736
rect 291660 270292 291712 270298
rect 291660 270234 291712 270240
rect 291764 264330 291792 271730
rect 291686 264302 291792 264330
rect 292132 264316 292160 273158
rect 292580 273148 292632 273154
rect 292580 273090 292632 273096
rect 292592 264316 292620 273090
rect 292868 270026 292896 277780
rect 293408 273080 293460 273086
rect 293408 273022 293460 273028
rect 292856 270020 292908 270026
rect 292856 269962 292908 269968
rect 292948 269068 293000 269074
rect 292948 269010 293000 269016
rect 292960 264316 292988 269010
rect 293420 264316 293448 273022
rect 293868 273012 293920 273018
rect 293868 272954 293920 272960
rect 293880 264316 293908 272954
rect 294064 270094 294092 277780
rect 295064 272332 295116 272338
rect 295064 272274 295116 272280
rect 294328 270428 294380 270434
rect 294328 270370 294380 270376
rect 294052 270088 294104 270094
rect 294052 270030 294104 270036
rect 294340 264316 294368 270370
rect 295076 264330 295104 272274
rect 295168 270162 295196 277780
rect 296076 272740 296128 272746
rect 296076 272682 296128 272688
rect 295248 272536 295300 272542
rect 295248 272478 295300 272484
rect 295156 270156 295208 270162
rect 295156 270098 295208 270104
rect 294814 264302 295104 264330
rect 295260 264316 295288 272478
rect 295616 269000 295668 269006
rect 295616 268942 295668 268948
rect 295628 264316 295656 268942
rect 296088 264316 296116 272682
rect 296364 269890 296392 277780
rect 296996 270360 297048 270366
rect 296996 270302 297048 270308
rect 296536 270224 296588 270230
rect 296536 270166 296588 270172
rect 296352 269884 296404 269890
rect 296352 269826 296404 269832
rect 296548 264316 296576 270166
rect 297008 264316 297036 270302
rect 297456 270292 297508 270298
rect 297456 270234 297508 270240
rect 297468 264316 297496 270234
rect 297560 269958 297588 277780
rect 298284 270156 298336 270162
rect 298284 270098 298336 270104
rect 297548 269952 297600 269958
rect 297548 269894 297600 269900
rect 297916 267912 297968 267918
rect 297916 267854 297968 267860
rect 297928 264316 297956 267854
rect 298296 264316 298324 270098
rect 298756 269754 298784 277780
rect 299204 270088 299256 270094
rect 299204 270030 299256 270036
rect 298744 269748 298796 269754
rect 298744 269690 298796 269696
rect 298744 267980 298796 267986
rect 298744 267922 298796 267928
rect 298756 264316 298784 267922
rect 299216 264316 299244 270030
rect 299952 269822 299980 277780
rect 300768 272808 300820 272814
rect 300768 272750 300820 272756
rect 300676 272672 300728 272678
rect 300676 272614 300728 272620
rect 299940 269816 299992 269822
rect 299940 269758 299992 269764
rect 299664 267164 299716 267170
rect 299664 267106 299716 267112
rect 299676 264316 299704 267106
rect 300688 264974 300716 272614
rect 300504 264946 300716 264974
rect 300504 264330 300532 264946
rect 300780 264330 300808 272750
rect 301148 269550 301176 277780
rect 301412 272604 301464 272610
rect 301412 272546 301464 272552
rect 301136 269544 301188 269550
rect 301136 269486 301188 269492
rect 300952 267096 301004 267102
rect 300952 267038 301004 267044
rect 300150 264302 300532 264330
rect 300610 264302 300808 264330
rect 300964 264316 300992 267038
rect 301424 264316 301452 272546
rect 301872 272468 301924 272474
rect 301872 272410 301924 272416
rect 301884 264316 301912 272410
rect 302344 269618 302372 277780
rect 303344 272264 303396 272270
rect 303344 272206 303396 272212
rect 302332 269612 302384 269618
rect 302332 269554 302384 269560
rect 302332 267028 302384 267034
rect 302332 266970 302384 266976
rect 302344 264316 302372 266970
rect 303356 264974 303384 272206
rect 303448 269686 303476 277780
rect 303528 272400 303580 272406
rect 303528 272342 303580 272348
rect 303436 269680 303488 269686
rect 303436 269622 303488 269628
rect 303172 264946 303384 264974
rect 303172 264330 303200 264946
rect 303540 264330 303568 272342
rect 304080 270496 304132 270502
rect 304080 270438 304132 270444
rect 303712 266960 303764 266966
rect 303712 266902 303764 266908
rect 302818 264302 303200 264330
rect 303278 264302 303568 264330
rect 303724 264316 303752 266902
rect 304092 264316 304120 270438
rect 304644 269414 304672 277780
rect 304908 272944 304960 272950
rect 304908 272886 304960 272892
rect 304632 269408 304684 269414
rect 304632 269350 304684 269356
rect 304920 267918 304948 272886
rect 305460 269952 305512 269958
rect 305460 269894 305512 269900
rect 304908 267912 304960 267918
rect 304908 267854 304960 267860
rect 304540 267844 304592 267850
rect 304540 267786 304592 267792
rect 304552 264316 304580 267786
rect 305000 266892 305052 266898
rect 305000 266834 305052 266840
rect 305012 264316 305040 266834
rect 305472 264316 305500 269894
rect 305840 269482 305868 277780
rect 306288 272196 306340 272202
rect 306288 272138 306340 272144
rect 305828 269476 305880 269482
rect 305828 269418 305880 269424
rect 306300 264330 306328 272138
rect 306748 269884 306800 269890
rect 306748 269826 306800 269832
rect 306380 266824 306432 266830
rect 306380 266766 306432 266772
rect 305946 264302 306328 264330
rect 306392 264316 306420 266766
rect 306760 264316 306788 269826
rect 307036 269278 307064 277780
rect 307852 272876 307904 272882
rect 307852 272818 307904 272824
rect 307208 269816 307260 269822
rect 307208 269758 307260 269764
rect 307024 269272 307076 269278
rect 307024 269214 307076 269220
rect 307220 264316 307248 269758
rect 307864 267986 307892 272818
rect 308128 269748 308180 269754
rect 308128 269690 308180 269696
rect 307852 267980 307904 267986
rect 307852 267922 307904 267928
rect 307668 266756 307720 266762
rect 307668 266698 307720 266704
rect 307680 264316 307708 266698
rect 308140 264316 308168 269690
rect 308232 269346 308260 277780
rect 308956 272128 309008 272134
rect 308956 272070 309008 272076
rect 308220 269340 308272 269346
rect 308220 269282 308272 269288
rect 308968 264330 308996 272070
rect 309428 272066 309456 277780
rect 309416 272060 309468 272066
rect 309416 272002 309468 272008
rect 310532 269142 310560 277780
rect 311624 272060 311676 272066
rect 311624 272002 311676 272008
rect 310796 269612 310848 269618
rect 310796 269554 310848 269560
rect 310520 269136 310572 269142
rect 310520 269078 310572 269084
rect 309876 268932 309928 268938
rect 309876 268874 309928 268880
rect 309416 268388 309468 268394
rect 309416 268330 309468 268336
rect 309048 266688 309100 266694
rect 309048 266630 309100 266636
rect 308614 264302 308996 264330
rect 309060 264316 309088 266630
rect 309428 264316 309456 268330
rect 309888 264316 309916 268874
rect 310336 266620 310388 266626
rect 310336 266562 310388 266568
rect 310348 264316 310376 266562
rect 310808 264316 310836 269554
rect 311636 264330 311664 272002
rect 311728 269210 311756 277780
rect 312924 271998 312952 277780
rect 312912 271992 312964 271998
rect 312912 271934 312964 271940
rect 314120 270978 314148 277780
rect 314292 271992 314344 271998
rect 314292 271934 314344 271940
rect 314108 270972 314160 270978
rect 314108 270914 314160 270920
rect 312084 269544 312136 269550
rect 312084 269486 312136 269492
rect 311716 269204 311768 269210
rect 311716 269146 311768 269152
rect 311716 266552 311768 266558
rect 311716 266494 311768 266500
rect 311282 264302 311664 264330
rect 311728 264316 311756 266494
rect 312096 264316 312124 269486
rect 313464 269476 313516 269482
rect 313464 269418 313516 269424
rect 312544 268320 312596 268326
rect 312544 268262 312596 268268
rect 312556 264316 312584 268262
rect 313004 266484 313056 266490
rect 313004 266426 313056 266432
rect 313016 264316 313044 266426
rect 313476 264316 313504 269418
rect 314304 264330 314332 271934
rect 315316 271114 315344 277780
rect 316512 271318 316540 277780
rect 316500 271312 316552 271318
rect 316500 271254 316552 271260
rect 317708 271182 317736 277780
rect 318812 271386 318840 277780
rect 318892 274848 318944 274854
rect 318892 274790 318944 274796
rect 318800 271380 318852 271386
rect 318800 271322 318852 271328
rect 317696 271176 317748 271182
rect 317696 271118 317748 271124
rect 315304 271108 315356 271114
rect 315304 271050 315356 271056
rect 314844 269408 314896 269414
rect 314844 269350 314896 269356
rect 314384 265260 314436 265266
rect 314384 265202 314436 265208
rect 313950 264302 314332 264330
rect 314396 264316 314424 265202
rect 314856 264316 314884 269350
rect 315212 269340 315264 269346
rect 315212 269282 315264 269288
rect 315224 264316 315252 269282
rect 317880 269272 317932 269278
rect 317880 269214 317932 269220
rect 316132 268252 316184 268258
rect 316132 268194 316184 268200
rect 315672 266416 315724 266422
rect 315672 266358 315724 266364
rect 315684 264316 315712 266358
rect 316144 264316 316172 268194
rect 316592 268184 316644 268190
rect 316592 268126 316644 268132
rect 316604 264316 316632 268126
rect 317052 266348 317104 266354
rect 317052 266290 317104 266296
rect 317064 264316 317092 266290
rect 317512 265804 317564 265810
rect 317512 265746 317564 265752
rect 317524 264316 317552 265746
rect 317892 264316 317920 269214
rect 318340 265328 318392 265334
rect 318340 265270 318392 265276
rect 318352 264316 318380 265270
rect 318904 264330 318932 274790
rect 320008 271250 320036 277780
rect 320180 274780 320232 274786
rect 320180 274722 320232 274728
rect 319996 271244 320048 271250
rect 319996 271186 320048 271192
rect 319260 268048 319312 268054
rect 319260 267990 319312 267996
rect 318826 264302 318932 264330
rect 319272 264316 319300 267990
rect 319720 265192 319772 265198
rect 319720 265134 319772 265140
rect 319732 264316 319760 265134
rect 320192 264316 320220 274722
rect 321008 274712 321060 274718
rect 321008 274654 321060 274660
rect 320548 269204 320600 269210
rect 320548 269146 320600 269152
rect 320560 264316 320588 269146
rect 321020 264316 321048 274654
rect 321204 271454 321232 277780
rect 322400 271522 322428 277780
rect 322848 274644 322900 274650
rect 322848 274586 322900 274592
rect 322388 271516 322440 271522
rect 322388 271458 322440 271464
rect 321192 271448 321244 271454
rect 321192 271390 321244 271396
rect 321928 267980 321980 267986
rect 321928 267922 321980 267928
rect 321468 265396 321520 265402
rect 321468 265338 321520 265344
rect 321480 264316 321508 265338
rect 321940 264316 321968 267922
rect 322860 264974 322888 274586
rect 323596 271862 323624 277780
rect 323676 273624 323728 273630
rect 323676 273566 323728 273572
rect 323584 271856 323636 271862
rect 323584 271798 323636 271804
rect 323216 269136 323268 269142
rect 323216 269078 323268 269084
rect 322940 265464 322992 265470
rect 322940 265406 322992 265412
rect 322768 264946 322888 264974
rect 322768 264330 322796 264946
rect 322952 264330 322980 265406
rect 322414 264302 322796 264330
rect 322874 264302 322980 264330
rect 323228 264316 323256 269078
rect 323688 264316 323716 273566
rect 324792 271658 324820 277780
rect 325424 273760 325476 273766
rect 325424 273702 325476 273708
rect 324780 271652 324832 271658
rect 324780 271594 324832 271600
rect 324596 270632 324648 270638
rect 324596 270574 324648 270580
rect 324136 265532 324188 265538
rect 324136 265474 324188 265480
rect 324148 264316 324176 265474
rect 324608 264316 324636 270574
rect 325436 264330 325464 273702
rect 325988 271930 326016 277780
rect 326804 273828 326856 273834
rect 326804 273770 326856 273776
rect 326344 273692 326396 273698
rect 326344 273634 326396 273640
rect 325976 271924 326028 271930
rect 325976 271866 326028 271872
rect 325608 271856 325660 271862
rect 325608 271798 325660 271804
rect 325620 267986 325648 271798
rect 325976 268456 326028 268462
rect 325976 268398 326028 268404
rect 325608 267980 325660 267986
rect 325608 267922 325660 267928
rect 325516 265600 325568 265606
rect 325516 265542 325568 265548
rect 325082 264302 325464 264330
rect 325528 264316 325556 265542
rect 325988 264316 326016 268398
rect 326356 264316 326384 273634
rect 326712 271924 326764 271930
rect 326712 271866 326764 271872
rect 326436 270768 326488 270774
rect 326436 270710 326488 270716
rect 326448 268190 326476 270710
rect 326436 268184 326488 268190
rect 326436 268126 326488 268132
rect 326724 268054 326752 271866
rect 326712 268048 326764 268054
rect 326712 267990 326764 267996
rect 326816 264316 326844 273770
rect 327092 271726 327120 277780
rect 327724 273964 327776 273970
rect 327724 273906 327776 273912
rect 327080 271720 327132 271726
rect 327080 271662 327132 271668
rect 327264 270904 327316 270910
rect 327264 270846 327316 270852
rect 327276 264316 327304 270846
rect 327736 264316 327764 273906
rect 328288 271590 328316 277780
rect 329104 273896 329156 273902
rect 329104 273838 329156 273844
rect 328276 271584 328328 271590
rect 328276 271526 328328 271532
rect 329012 270836 329064 270842
rect 329012 270778 329064 270784
rect 329024 269006 329052 270778
rect 329012 269000 329064 269006
rect 329012 268942 329064 268948
rect 328644 268864 328696 268870
rect 328644 268806 328696 268812
rect 328000 267912 328052 267918
rect 328000 267854 328052 267860
rect 328012 264330 328040 267854
rect 328012 264302 328210 264330
rect 328656 264316 328684 268806
rect 329116 264330 329144 273838
rect 329484 271794 329512 277780
rect 330392 273556 330444 273562
rect 330392 273498 330444 273504
rect 329472 271788 329524 271794
rect 329472 271730 329524 271736
rect 329932 270972 329984 270978
rect 329932 270914 329984 270920
rect 329472 265736 329524 265742
rect 329472 265678 329524 265684
rect 329038 264302 329144 264330
rect 329484 264316 329512 265678
rect 329944 264316 329972 270914
rect 330404 264316 330432 273498
rect 330680 273222 330708 277780
rect 331680 274032 331732 274038
rect 331680 273974 331732 273980
rect 330668 273216 330720 273222
rect 330668 273158 330720 273164
rect 331312 271040 331364 271046
rect 331312 270982 331364 270988
rect 331128 270700 331180 270706
rect 331128 270642 331180 270648
rect 330852 269000 330904 269006
rect 330852 268942 330904 268948
rect 330864 264316 330892 268942
rect 331140 268938 331168 270642
rect 331128 268932 331180 268938
rect 331128 268874 331180 268880
rect 331324 264316 331352 270982
rect 331692 264316 331720 273974
rect 331876 273154 331904 277780
rect 332140 274168 332192 274174
rect 332140 274110 332192 274116
rect 331864 273148 331916 273154
rect 331864 273090 331916 273096
rect 331956 273148 332008 273154
rect 331956 273090 332008 273096
rect 331968 272338 331996 273090
rect 331956 272332 332008 272338
rect 331956 272274 332008 272280
rect 332152 264316 332180 274110
rect 332508 272944 332560 272950
rect 332508 272886 332560 272892
rect 332520 272338 332548 272886
rect 332508 272332 332560 272338
rect 332508 272274 332560 272280
rect 333072 269074 333100 277780
rect 333428 274236 333480 274242
rect 333428 274178 333480 274184
rect 333060 269068 333112 269074
rect 333060 269010 333112 269016
rect 332784 268456 332836 268462
rect 332784 268398 332836 268404
rect 332508 268388 332560 268394
rect 332508 268330 332560 268336
rect 332600 268388 332652 268394
rect 332600 268330 332652 268336
rect 332520 267782 332548 268330
rect 332508 267776 332560 267782
rect 332508 267718 332560 267724
rect 332612 264316 332640 268330
rect 332692 268252 332744 268258
rect 332692 268194 332744 268200
rect 332704 267918 332732 268194
rect 332796 268122 332824 268398
rect 332784 268116 332836 268122
rect 332784 268058 332836 268064
rect 332692 267912 332744 267918
rect 332692 267854 332744 267860
rect 333440 264330 333468 274178
rect 334176 273086 334204 277780
rect 334348 274304 334400 274310
rect 334348 274246 334400 274252
rect 334164 273080 334216 273086
rect 334164 273022 334216 273028
rect 333980 271176 334032 271182
rect 333980 271118 334032 271124
rect 333520 268456 333572 268462
rect 333520 268398 333572 268404
rect 333086 264302 333468 264330
rect 333532 264316 333560 268398
rect 333992 264316 334020 271118
rect 334360 264316 334388 274246
rect 335372 273018 335400 277780
rect 335728 274372 335780 274378
rect 335728 274314 335780 274320
rect 335360 273012 335412 273018
rect 335360 272954 335412 272960
rect 334808 271108 334860 271114
rect 334808 271050 334860 271056
rect 334820 264316 334848 271050
rect 335268 268524 335320 268530
rect 335268 268466 335320 268472
rect 335280 264316 335308 268466
rect 335740 264316 335768 274314
rect 336464 271312 336516 271318
rect 336464 271254 336516 271260
rect 336188 268592 336240 268598
rect 336188 268534 336240 268540
rect 336200 264316 336228 268534
rect 336476 264330 336504 271254
rect 336568 270434 336596 277780
rect 337108 274440 337160 274446
rect 337108 274382 337160 274388
rect 336740 271720 336792 271726
rect 336740 271662 336792 271668
rect 336556 270428 336608 270434
rect 336556 270370 336608 270376
rect 336752 270366 336780 271662
rect 336740 270360 336792 270366
rect 336740 270302 336792 270308
rect 336476 264302 336674 264330
rect 337120 264316 337148 274382
rect 337764 273154 337792 277780
rect 337752 273148 337804 273154
rect 337752 273090 337804 273096
rect 338960 272542 338988 277780
rect 339500 273216 339552 273222
rect 339500 273158 339552 273164
rect 338948 272536 339000 272542
rect 338948 272478 339000 272484
rect 339408 271380 339460 271386
rect 339408 271322 339460 271328
rect 337476 271244 337528 271250
rect 337476 271186 337528 271192
rect 337488 264316 337516 271186
rect 338856 268728 338908 268734
rect 338856 268670 338908 268676
rect 337936 268660 337988 268666
rect 337936 268602 337988 268608
rect 337948 264316 337976 268602
rect 338396 265872 338448 265878
rect 338396 265814 338448 265820
rect 338408 264316 338436 265814
rect 338868 264316 338896 268670
rect 339420 264330 339448 271322
rect 339512 270298 339540 273158
rect 340156 270842 340184 277780
rect 341064 274508 341116 274514
rect 341064 274450 341116 274456
rect 340236 271788 340288 271794
rect 340236 271730 340288 271736
rect 340144 270836 340196 270842
rect 340144 270778 340196 270784
rect 339500 270292 339552 270298
rect 339500 270234 339552 270240
rect 339776 265940 339828 265946
rect 339776 265882 339828 265888
rect 339342 264302 339448 264330
rect 339788 264316 339816 265882
rect 340248 264330 340276 271730
rect 340328 270836 340380 270842
rect 340328 270778 340380 270784
rect 340340 270638 340368 270778
rect 340328 270632 340380 270638
rect 340328 270574 340380 270580
rect 340604 268796 340656 268802
rect 340604 268738 340656 268744
rect 340170 264302 340276 264330
rect 340616 264316 340644 268738
rect 341076 264316 341104 274450
rect 341352 272746 341380 277780
rect 341340 272740 341392 272746
rect 341340 272682 341392 272688
rect 342168 271516 342220 271522
rect 342168 271458 342220 271464
rect 341524 268864 341576 268870
rect 341524 268806 341576 268812
rect 341536 264316 341564 268806
rect 342180 264330 342208 271458
rect 342456 270230 342484 277780
rect 342536 274576 342588 274582
rect 342536 274518 342588 274524
rect 342444 270224 342496 270230
rect 342444 270166 342496 270172
rect 342548 264330 342576 274518
rect 342812 272536 342864 272542
rect 342812 272478 342864 272484
rect 342010 264302 342208 264330
rect 342470 264302 342576 264330
rect 342824 264316 342852 272478
rect 343652 271726 343680 277780
rect 343732 275936 343784 275942
rect 343732 275878 343784 275884
rect 343640 271720 343692 271726
rect 343640 271662 343692 271668
rect 343272 269680 343324 269686
rect 343272 269622 343324 269628
rect 343284 264316 343312 269622
rect 343744 264316 343772 275878
rect 344848 273222 344876 277780
rect 345112 276004 345164 276010
rect 345112 275946 345164 275952
rect 344836 273216 344888 273222
rect 344836 273158 344888 273164
rect 344008 273012 344060 273018
rect 344008 272954 344060 272960
rect 344020 270502 344048 272954
rect 344928 272740 344980 272746
rect 344928 272682 344980 272688
rect 344008 270496 344060 270502
rect 344008 270438 344060 270444
rect 344192 267912 344244 267918
rect 344192 267854 344244 267860
rect 344204 264316 344232 267854
rect 344940 264330 344968 272682
rect 344678 264302 344968 264330
rect 345124 264316 345152 275946
rect 346044 272338 346072 277780
rect 346032 272332 346084 272338
rect 346032 272274 346084 272280
rect 346860 270496 346912 270502
rect 346860 270438 346912 270444
rect 345480 270020 345532 270026
rect 345480 269962 345532 269968
rect 345492 264316 345520 269962
rect 345940 269000 345992 269006
rect 345940 268942 345992 268948
rect 345952 264316 345980 268942
rect 346400 266008 346452 266014
rect 346400 265950 346452 265956
rect 346412 264316 346440 265950
rect 346872 264316 346900 270438
rect 347240 270162 347268 277780
rect 348436 272882 348464 277780
rect 349068 275868 349120 275874
rect 349068 275810 349120 275816
rect 348424 272876 348476 272882
rect 348424 272818 348476 272824
rect 348240 271584 348292 271590
rect 348240 271526 348292 271532
rect 347596 271448 347648 271454
rect 347596 271390 347648 271396
rect 347228 270156 347280 270162
rect 347228 270098 347280 270104
rect 347608 264330 347636 271390
rect 347780 266076 347832 266082
rect 347780 266018 347832 266024
rect 347346 264302 347636 264330
rect 347792 264316 347820 266018
rect 348252 264316 348280 271526
rect 348608 270428 348660 270434
rect 348608 270370 348660 270376
rect 348620 264316 348648 270370
rect 349080 264316 349108 275810
rect 349528 270360 349580 270366
rect 349528 270302 349580 270308
rect 349540 264316 349568 270302
rect 349632 270094 349660 277780
rect 350356 275800 350408 275806
rect 350356 275742 350408 275748
rect 350264 271652 350316 271658
rect 350264 271594 350316 271600
rect 349620 270088 349672 270094
rect 349620 270030 349672 270036
rect 350276 264330 350304 271594
rect 350014 264302 350304 264330
rect 350368 264330 350396 275742
rect 350736 267170 350764 277780
rect 351828 274100 351880 274106
rect 351828 274042 351880 274048
rect 351840 273562 351868 274042
rect 351828 273556 351880 273562
rect 351828 273498 351880 273504
rect 351932 272678 351960 277780
rect 353128 272814 353156 277780
rect 353116 272808 353168 272814
rect 353116 272750 353168 272756
rect 351920 272672 351972 272678
rect 351920 272614 351972 272620
rect 353024 272672 353076 272678
rect 353024 272614 353076 272620
rect 351828 272332 351880 272338
rect 351828 272274 351880 272280
rect 351840 271794 351868 272274
rect 351828 271788 351880 271794
rect 351828 271730 351880 271736
rect 352380 271720 352432 271726
rect 352380 271662 352432 271668
rect 352104 271584 352156 271590
rect 351932 271532 352104 271538
rect 351932 271526 352156 271532
rect 351932 271510 352144 271526
rect 351932 271454 351960 271510
rect 351920 271448 351972 271454
rect 351920 271390 351972 271396
rect 352012 270632 352064 270638
rect 352012 270574 352064 270580
rect 351276 270292 351328 270298
rect 351276 270234 351328 270240
rect 350908 270156 350960 270162
rect 350908 270098 350960 270104
rect 350724 267164 350776 267170
rect 350724 267106 350776 267112
rect 350368 264302 350474 264330
rect 350920 264316 350948 270098
rect 351288 264316 351316 270234
rect 351736 270020 351788 270026
rect 351736 269962 351788 269968
rect 351748 267850 351776 269962
rect 351828 269068 351880 269074
rect 351828 269010 351880 269016
rect 351840 268326 351868 269010
rect 351920 268932 351972 268938
rect 351920 268874 351972 268880
rect 351828 268320 351880 268326
rect 351828 268262 351880 268268
rect 351932 268190 351960 268874
rect 351920 268184 351972 268190
rect 351920 268126 351972 268132
rect 352024 267986 352052 270574
rect 352196 270224 352248 270230
rect 352196 270166 352248 270172
rect 352104 268932 352156 268938
rect 352104 268874 352156 268880
rect 352012 267980 352064 267986
rect 352012 267922 352064 267928
rect 352116 267918 352144 268874
rect 352104 267912 352156 267918
rect 352104 267854 352156 267860
rect 351736 267844 351788 267850
rect 351736 267786 351788 267792
rect 351736 266144 351788 266150
rect 351736 266086 351788 266092
rect 351748 264316 351776 266086
rect 352208 264316 352236 270166
rect 352392 270162 352420 271662
rect 352380 270156 352432 270162
rect 352380 270098 352432 270104
rect 352288 269680 352340 269686
rect 352288 269622 352340 269628
rect 352300 269006 352328 269622
rect 352288 269000 352340 269006
rect 352288 268942 352340 268948
rect 353036 264330 353064 272614
rect 353576 270156 353628 270162
rect 353576 270098 353628 270104
rect 353116 266212 353168 266218
rect 353116 266154 353168 266160
rect 352682 264302 353064 264330
rect 353128 264316 353156 266154
rect 353588 264316 353616 270098
rect 353942 268288 353998 268297
rect 353942 268223 353998 268232
rect 353956 264316 353984 268223
rect 354324 267102 354352 277780
rect 354404 275732 354456 275738
rect 354404 275674 354456 275680
rect 354312 267096 354364 267102
rect 354312 267038 354364 267044
rect 354416 264316 354444 275674
rect 355324 273148 355376 273154
rect 355324 273090 355376 273096
rect 354864 272876 354916 272882
rect 354864 272818 354916 272824
rect 354876 264316 354904 272818
rect 355336 264316 355364 273090
rect 355520 272610 355548 277780
rect 355784 275664 355836 275670
rect 355784 275606 355836 275612
rect 355508 272604 355560 272610
rect 355508 272546 355560 272552
rect 355796 264316 355824 275606
rect 356716 272474 356744 277780
rect 356704 272468 356756 272474
rect 356704 272410 356756 272416
rect 355968 271448 356020 271454
rect 355968 271390 356020 271396
rect 355980 270094 356008 271390
rect 357440 270564 357492 270570
rect 357440 270506 357492 270512
rect 355968 270088 356020 270094
rect 355968 270030 356020 270036
rect 356244 270088 356296 270094
rect 356244 270030 356296 270036
rect 356256 264316 356284 270030
rect 356610 268424 356666 268433
rect 356610 268359 356666 268368
rect 356624 264316 356652 268359
rect 357452 268054 357480 270506
rect 357440 268048 357492 268054
rect 357440 267990 357492 267996
rect 357532 268048 357584 268054
rect 357532 267990 357584 267996
rect 357072 266280 357124 266286
rect 357072 266222 357124 266228
rect 357084 264316 357112 266222
rect 357544 264316 357572 267990
rect 357912 267034 357940 277780
rect 358452 275596 358504 275602
rect 358452 275538 358504 275544
rect 357992 272944 358044 272950
rect 357992 272886 358044 272892
rect 357900 267028 357952 267034
rect 357900 266970 357952 266976
rect 358004 264316 358032 272886
rect 358464 264316 358492 275538
rect 358820 273080 358872 273086
rect 358820 273022 358872 273028
rect 358728 268048 358780 268054
rect 358832 268036 358860 273022
rect 359016 272270 359044 277780
rect 360212 272406 360240 277780
rect 361120 275528 361172 275534
rect 361120 275470 361172 275476
rect 360660 272808 360712 272814
rect 360660 272750 360712 272756
rect 360568 272468 360620 272474
rect 360568 272410 360620 272416
rect 360200 272400 360252 272406
rect 360200 272342 360252 272348
rect 359004 272264 359056 272270
rect 359004 272206 359056 272212
rect 358910 268696 358966 268705
rect 358910 268631 358966 268640
rect 358780 268008 358860 268036
rect 358728 267990 358780 267996
rect 358924 264316 358952 268631
rect 359370 268560 359426 268569
rect 359370 268495 359426 268504
rect 359384 264316 359412 268495
rect 359740 267708 359792 267714
rect 359740 267650 359792 267656
rect 359752 264316 359780 267650
rect 360580 264330 360608 272410
rect 360226 264302 360608 264330
rect 360672 264316 360700 272750
rect 361132 264316 361160 275470
rect 361408 266966 361436 277780
rect 362604 273018 362632 277780
rect 362776 273216 362828 273222
rect 362776 273158 362828 273164
rect 362592 273012 362644 273018
rect 362592 272954 362644 272960
rect 362788 272678 362816 273158
rect 363144 273080 363196 273086
rect 362880 273028 363144 273034
rect 362880 273022 363196 273028
rect 362880 273006 363184 273022
rect 362880 272882 362908 273006
rect 362868 272876 362920 272882
rect 362868 272818 362920 272824
rect 363236 272808 363288 272814
rect 363236 272750 363288 272756
rect 362776 272672 362828 272678
rect 362776 272614 362828 272620
rect 363144 272672 363196 272678
rect 363144 272614 363196 272620
rect 361580 269680 361632 269686
rect 361580 269622 361632 269628
rect 361396 266960 361448 266966
rect 361396 266902 361448 266908
rect 361592 264316 361620 269622
rect 362038 268832 362094 268841
rect 362038 268767 362094 268776
rect 362052 264316 362080 268767
rect 362408 267640 362460 267646
rect 362408 267582 362460 267588
rect 362420 264316 362448 267582
rect 363156 264330 363184 272614
rect 363248 272474 363276 272750
rect 363236 272468 363288 272474
rect 363236 272410 363288 272416
rect 363326 271416 363382 271425
rect 363326 271351 363382 271360
rect 362894 264302 363184 264330
rect 363340 264316 363368 271351
rect 363800 270026 363828 277780
rect 364064 275460 364116 275466
rect 364064 275402 364116 275408
rect 363788 270020 363840 270026
rect 363788 269962 363840 269968
rect 364076 264330 364104 275402
rect 364708 270020 364760 270026
rect 364708 269962 364760 269968
rect 364246 268968 364302 268977
rect 364246 268903 364302 268912
rect 363814 264302 364104 264330
rect 364260 264316 364288 268903
rect 364720 264316 364748 269962
rect 364996 266898 365024 277780
rect 365994 271688 366050 271697
rect 365994 271623 366050 271632
rect 365534 271552 365590 271561
rect 365534 271487 365590 271496
rect 365076 267572 365128 267578
rect 365076 267514 365128 267520
rect 364984 266892 365036 266898
rect 364984 266834 365036 266840
rect 365088 264316 365116 267514
rect 365548 264316 365576 271487
rect 366008 264316 366036 271623
rect 366100 269958 366128 277780
rect 366456 275392 366508 275398
rect 366456 275334 366508 275340
rect 366088 269952 366140 269958
rect 366088 269894 366140 269900
rect 366468 264316 366496 275334
rect 367296 272202 367324 277780
rect 368204 272604 368256 272610
rect 368204 272546 368256 272552
rect 367284 272196 367336 272202
rect 367284 272138 367336 272144
rect 366914 270464 366970 270473
rect 366914 270399 366970 270408
rect 366928 264316 366956 270399
rect 367376 269952 367428 269958
rect 367376 269894 367428 269900
rect 367388 264316 367416 269894
rect 367744 267504 367796 267510
rect 367744 267446 367796 267452
rect 367756 264316 367784 267446
rect 368216 264316 368244 272546
rect 368492 266830 368520 277780
rect 369124 275324 369176 275330
rect 369124 275266 369176 275272
rect 368662 273184 368718 273193
rect 368662 273119 368718 273128
rect 368480 266824 368532 266830
rect 368480 266766 368532 266772
rect 368676 264316 368704 273119
rect 369136 264316 369164 275266
rect 369582 270328 369638 270337
rect 369582 270263 369638 270272
rect 369596 264316 369624 270263
rect 369688 269890 369716 277780
rect 369676 269884 369728 269890
rect 369676 269826 369728 269832
rect 370044 269884 370096 269890
rect 370044 269826 370096 269832
rect 370056 264316 370084 269826
rect 370884 269822 370912 277780
rect 371792 275256 371844 275262
rect 371792 275198 371844 275204
rect 371238 273048 371294 273057
rect 371238 272983 371294 272992
rect 370872 269816 370924 269822
rect 370872 269758 370924 269764
rect 370504 267436 370556 267442
rect 370504 267378 370556 267384
rect 370516 264316 370544 267378
rect 371252 264330 371280 272983
rect 371330 272912 371386 272921
rect 371330 272847 371386 272856
rect 370898 264302 371280 264330
rect 371344 264316 371372 272847
rect 371804 264316 371832 275198
rect 372080 266762 372108 277780
rect 373172 272468 373224 272474
rect 373172 272410 373224 272416
rect 372250 270192 372306 270201
rect 372250 270127 372306 270136
rect 372068 266756 372120 266762
rect 372068 266698 372120 266704
rect 372264 264316 372292 270127
rect 372712 268048 372764 268054
rect 372712 267990 372764 267996
rect 372724 264316 372752 267990
rect 373184 264316 373212 272410
rect 373276 269822 373304 277780
rect 373998 272776 374054 272785
rect 373998 272711 374054 272720
rect 373264 269816 373316 269822
rect 373264 269758 373316 269764
rect 373540 267368 373592 267374
rect 373540 267310 373592 267316
rect 373552 264316 373580 267310
rect 374012 264316 374040 272711
rect 374380 272134 374408 277780
rect 374920 275188 374972 275194
rect 374920 275130 374972 275136
rect 374368 272128 374420 272134
rect 374368 272070 374420 272076
rect 374460 267300 374512 267306
rect 374460 267242 374512 267248
rect 374472 264316 374500 267242
rect 374932 264316 374960 275130
rect 375380 269748 375432 269754
rect 375380 269690 375432 269696
rect 375392 264316 375420 269690
rect 375576 266694 375604 277780
rect 376668 272400 376720 272406
rect 376668 272342 376720 272348
rect 376208 267232 376260 267238
rect 376208 267174 376260 267180
rect 375840 267164 375892 267170
rect 375840 267106 375892 267112
rect 375564 266688 375616 266694
rect 375564 266630 375616 266636
rect 375852 264316 375880 267106
rect 376220 264316 376248 267174
rect 376680 264316 376708 272342
rect 376772 267782 376800 277780
rect 377588 275120 377640 275126
rect 377588 275062 377640 275068
rect 376760 267776 376812 267782
rect 376760 267718 376812 267724
rect 377128 267096 377180 267102
rect 377128 267038 377180 267044
rect 377140 264316 377168 267038
rect 377600 264316 377628 275062
rect 377968 270706 377996 277780
rect 377956 270700 378008 270706
rect 377956 270642 378008 270648
rect 378046 270056 378102 270065
rect 378046 269991 378102 270000
rect 378060 264316 378088 269991
rect 378508 267028 378560 267034
rect 378508 266970 378560 266976
rect 378520 264316 378548 266970
rect 378876 266960 378928 266966
rect 378876 266902 378928 266908
rect 378888 264316 378916 266902
rect 379164 266626 379192 277780
rect 380256 275052 380308 275058
rect 380256 274994 380308 275000
rect 379334 272640 379390 272649
rect 379334 272575 379390 272584
rect 379152 266620 379204 266626
rect 379152 266562 379204 266568
rect 379348 264316 379376 272575
rect 379796 266892 379848 266898
rect 379796 266834 379848 266840
rect 379808 264316 379836 266834
rect 380268 264316 380296 274994
rect 380360 269618 380388 277780
rect 381556 272066 381584 277780
rect 382004 272264 382056 272270
rect 382004 272206 382056 272212
rect 381544 272060 381596 272066
rect 381544 272002 381596 272008
rect 380348 269612 380400 269618
rect 380348 269554 380400 269560
rect 380716 269612 380768 269618
rect 380716 269554 380768 269560
rect 380728 264316 380756 269554
rect 381636 266824 381688 266830
rect 381636 266766 381688 266772
rect 381176 266756 381228 266762
rect 381176 266698 381228 266704
rect 381188 264316 381216 266698
rect 381648 264316 381676 266766
rect 382016 264316 382044 272206
rect 382464 270020 382516 270026
rect 382464 269962 382516 269968
rect 382476 269906 382504 269962
rect 382292 269878 382504 269906
rect 382292 269686 382320 269878
rect 382464 269748 382516 269754
rect 382464 269690 382516 269696
rect 382280 269680 382332 269686
rect 382280 269622 382332 269628
rect 382476 268054 382504 269690
rect 382464 268048 382516 268054
rect 382464 267990 382516 267996
rect 382464 266688 382516 266694
rect 382464 266630 382516 266636
rect 382188 266348 382240 266354
rect 382188 266290 382240 266296
rect 382200 265810 382228 266290
rect 382096 265804 382148 265810
rect 382096 265746 382148 265752
rect 382188 265804 382240 265810
rect 382188 265746 382240 265752
rect 382108 265690 382136 265746
rect 382108 265674 382320 265690
rect 382108 265668 382332 265674
rect 382108 265662 382280 265668
rect 382280 265610 382332 265616
rect 382476 264316 382504 266630
rect 382660 266558 382688 277780
rect 382924 274984 382976 274990
rect 382924 274926 382976 274932
rect 382648 266552 382700 266558
rect 382648 266494 382700 266500
rect 382936 264316 382964 274926
rect 383382 269920 383438 269929
rect 383382 269855 383438 269864
rect 383396 264316 383424 269855
rect 383856 269550 383884 277780
rect 384672 272196 384724 272202
rect 384672 272138 384724 272144
rect 383844 269544 383896 269550
rect 383844 269486 383896 269492
rect 384304 266620 384356 266626
rect 384304 266562 384356 266568
rect 383844 266552 383896 266558
rect 383844 266494 383896 266500
rect 383856 264316 383884 266494
rect 384316 264316 384344 266562
rect 384684 264316 384712 272138
rect 385052 270570 385080 277780
rect 385592 274916 385644 274922
rect 385592 274858 385644 274864
rect 385040 270564 385092 270570
rect 385040 270506 385092 270512
rect 385130 266112 385186 266121
rect 385130 266047 385186 266056
rect 385144 264316 385172 266047
rect 385604 264316 385632 274858
rect 386052 269544 386104 269550
rect 386052 269486 386104 269492
rect 386064 264316 386092 269486
rect 386248 266490 386276 277780
rect 387340 272128 387392 272134
rect 387340 272070 387392 272076
rect 386970 267608 387026 267617
rect 386970 267543 387026 267552
rect 386236 266484 386288 266490
rect 386236 266426 386288 266432
rect 386510 266248 386566 266257
rect 386510 266183 386566 266192
rect 386524 264316 386552 266183
rect 386984 264316 387012 267543
rect 387352 264316 387380 272070
rect 387444 269482 387472 277780
rect 388258 275904 388314 275913
rect 388258 275839 388314 275848
rect 387432 269476 387484 269482
rect 387432 269418 387484 269424
rect 387798 267744 387854 267753
rect 387798 267679 387854 267688
rect 387812 264316 387840 267679
rect 388272 264316 388300 275839
rect 388640 271998 388668 277780
rect 388628 271992 388680 271998
rect 388628 271934 388680 271940
rect 388720 269476 388772 269482
rect 388720 269418 388772 269424
rect 388732 264316 388760 269418
rect 389638 267472 389694 267481
rect 389638 267407 389694 267416
rect 389180 266484 389232 266490
rect 389180 266426 389232 266432
rect 389192 264316 389220 266426
rect 389652 264316 389680 267407
rect 389744 265266 389772 277780
rect 390940 269414 390968 277780
rect 391294 275768 391350 275777
rect 391294 275703 391350 275712
rect 390928 269408 390980 269414
rect 390928 269350 390980 269356
rect 390008 268048 390060 268054
rect 390008 267990 390060 267996
rect 389732 265260 389784 265266
rect 389732 265202 389784 265208
rect 390020 264316 390048 267990
rect 390466 267336 390522 267345
rect 390466 267271 390522 267280
rect 390480 264316 390508 267271
rect 391308 264330 391336 275703
rect 391386 269784 391442 269793
rect 391386 269719 391442 269728
rect 390954 264302 391336 264330
rect 391400 264316 391428 269719
rect 392136 269346 392164 277780
rect 392766 272504 392822 272513
rect 392766 272439 392822 272448
rect 392124 269340 392176 269346
rect 392124 269282 392176 269288
rect 391846 267200 391902 267209
rect 391846 267135 391902 267144
rect 391860 264316 391888 267135
rect 392308 266416 392360 266422
rect 392308 266358 392360 266364
rect 392320 264316 392348 266358
rect 392780 264316 392808 272439
rect 393134 267064 393190 267073
rect 393134 266999 393190 267008
rect 393148 264316 393176 266999
rect 393332 266354 393360 277780
rect 393594 275632 393650 275641
rect 393594 275567 393650 275576
rect 393320 266348 393372 266354
rect 393320 266290 393372 266296
rect 393608 264316 393636 275567
rect 394528 270638 394556 277780
rect 394608 272060 394660 272066
rect 394608 272002 394660 272008
rect 394516 270632 394568 270638
rect 394516 270574 394568 270580
rect 394056 269408 394108 269414
rect 394056 269350 394108 269356
rect 394068 264316 394096 269350
rect 394620 268054 394648 272002
rect 395436 271992 395488 271998
rect 395436 271934 395488 271940
rect 394608 268048 394660 268054
rect 394608 267990 394660 267996
rect 394514 266928 394570 266937
rect 394514 266863 394570 266872
rect 394528 264316 394556 266863
rect 394976 266348 395028 266354
rect 394976 266290 395028 266296
rect 394988 264316 395016 266290
rect 395448 264316 395476 271934
rect 395724 270774 395752 277780
rect 396262 275496 396318 275505
rect 396262 275431 396318 275440
rect 395712 270768 395764 270774
rect 395712 270710 395764 270716
rect 395802 266792 395858 266801
rect 395802 266727 395858 266736
rect 395816 264316 395844 266727
rect 396276 264316 396304 275431
rect 396724 269340 396776 269346
rect 396724 269282 396776 269288
rect 396736 264316 396764 269282
rect 396920 265810 396948 277780
rect 397182 266656 397238 266665
rect 397182 266591 397238 266600
rect 396908 265804 396960 265810
rect 396908 265746 396960 265752
rect 397196 264316 397224 266591
rect 397644 265804 397696 265810
rect 397644 265746 397696 265752
rect 397656 264316 397684 265746
rect 398024 265674 398052 277780
rect 398930 275360 398986 275369
rect 398930 275295 398986 275304
rect 398102 272368 398158 272377
rect 398102 272303 398158 272312
rect 398012 265668 398064 265674
rect 398012 265610 398064 265616
rect 398116 264316 398144 272303
rect 398470 266520 398526 266529
rect 398470 266455 398526 266464
rect 398484 264316 398512 266455
rect 398944 264316 398972 275295
rect 399220 269278 399248 277780
rect 399208 269272 399260 269278
rect 399208 269214 399260 269220
rect 399392 269272 399444 269278
rect 399392 269214 399444 269220
rect 399404 264316 399432 269214
rect 399850 266384 399906 266393
rect 399850 266319 399906 266328
rect 399864 264316 399892 266319
rect 400312 265668 400364 265674
rect 400312 265610 400364 265616
rect 400324 264316 400352 265610
rect 400416 265334 400444 277780
rect 401612 274854 401640 277780
rect 401690 275224 401746 275233
rect 401690 275159 401746 275168
rect 401600 274848 401652 274854
rect 401600 274790 401652 274796
rect 401140 273488 401192 273494
rect 401140 273430 401192 273436
rect 400772 268048 400824 268054
rect 400772 267990 400824 267996
rect 400404 265328 400456 265334
rect 400404 265270 400456 265276
rect 400784 264316 400812 267990
rect 401152 264316 401180 273430
rect 401704 264330 401732 275159
rect 402702 274952 402758 274961
rect 402702 274887 402758 274896
rect 402058 269648 402114 269657
rect 402058 269583 402114 269592
rect 401626 264302 401732 264330
rect 402072 264316 402100 269583
rect 402716 264330 402744 274887
rect 402808 271930 402836 277780
rect 403900 274848 403952 274854
rect 403900 274790 403952 274796
rect 403438 272232 403494 272241
rect 403438 272167 403494 272176
rect 402796 271924 402848 271930
rect 402796 271866 402848 271872
rect 402888 271924 402940 271930
rect 402888 271866 402940 271872
rect 402900 268054 402928 271866
rect 402888 268048 402940 268054
rect 402888 267990 402940 267996
rect 402980 265328 403032 265334
rect 402980 265270 403032 265276
rect 402546 264302 402744 264330
rect 402992 264316 403020 265270
rect 403452 264316 403480 272167
rect 403912 264316 403940 274790
rect 404004 265198 404032 277780
rect 404266 275088 404322 275097
rect 404266 275023 404322 275032
rect 403992 265192 404044 265198
rect 403992 265134 404044 265140
rect 404280 264316 404308 275023
rect 405200 274786 405228 277780
rect 405462 274816 405518 274825
rect 405188 274780 405240 274786
rect 405462 274751 405518 274760
rect 405188 274722 405240 274728
rect 404726 269512 404782 269521
rect 404726 269447 404782 269456
rect 404740 264316 404768 269447
rect 405476 264330 405504 274751
rect 406304 269210 406332 277780
rect 406568 274780 406620 274786
rect 406568 274722 406620 274728
rect 406292 269204 406344 269210
rect 406292 269146 406344 269152
rect 406108 268048 406160 268054
rect 406108 267990 406160 267996
rect 405646 265976 405702 265985
rect 405646 265911 405702 265920
rect 405214 264302 405504 264330
rect 405660 264316 405688 265911
rect 406120 264316 406148 267990
rect 406580 264316 406608 274722
rect 407500 274718 407528 277780
rect 407488 274712 407540 274718
rect 406934 274680 406990 274689
rect 407488 274654 407540 274660
rect 406934 274615 406990 274624
rect 406948 264316 406976 274615
rect 408222 274544 408278 274553
rect 408222 274479 408278 274488
rect 407394 269376 407450 269385
rect 407394 269311 407450 269320
rect 407408 264316 407436 269311
rect 408236 264330 408264 274479
rect 408314 265840 408370 265849
rect 408314 265775 408370 265784
rect 407882 264302 408264 264330
rect 408328 264316 408356 265775
rect 408696 265402 408724 277780
rect 409236 274712 409288 274718
rect 409236 274654 409288 274660
rect 408774 272096 408830 272105
rect 408774 272031 408830 272040
rect 408684 265396 408736 265402
rect 408684 265338 408736 265344
rect 408788 264316 408816 272031
rect 409248 264316 409276 274654
rect 409892 271862 409920 277780
rect 411088 274650 411116 277780
rect 411444 274848 411496 274854
rect 411444 274790 411496 274796
rect 411076 274644 411128 274650
rect 411076 274586 411128 274592
rect 411456 273494 411484 274790
rect 411444 273488 411496 273494
rect 411444 273430 411496 273436
rect 410522 271960 410578 271969
rect 410522 271895 410578 271904
rect 409880 271856 409932 271862
rect 409880 271798 409932 271804
rect 409602 269240 409658 269249
rect 409602 269175 409658 269184
rect 409616 264316 409644 269175
rect 410062 269104 410118 269113
rect 410062 269039 410118 269048
rect 410076 264316 410104 269039
rect 410536 264316 410564 271895
rect 410890 271824 410946 271833
rect 410890 271759 410946 271768
rect 410904 264330 410932 271759
rect 411812 270564 411864 270570
rect 411812 270506 411864 270512
rect 411444 269204 411496 269210
rect 411444 269146 411496 269152
rect 410904 264302 411010 264330
rect 411456 264316 411484 269146
rect 411824 269142 411852 270506
rect 411812 269136 411864 269142
rect 411812 269078 411864 269084
rect 411904 269136 411956 269142
rect 411904 269078 411956 269084
rect 411916 264316 411944 269078
rect 412284 265470 412312 277780
rect 413112 277766 413402 277794
rect 412824 271856 412876 271862
rect 412824 271798 412876 271804
rect 412836 268054 412864 271798
rect 413112 270570 413140 277766
rect 414584 273562 414612 277780
rect 414572 273556 414624 273562
rect 414572 273498 414624 273504
rect 413100 270564 413152 270570
rect 413100 270506 413152 270512
rect 412824 268048 412876 268054
rect 412824 267990 412876 267996
rect 415780 265538 415808 277780
rect 416976 270842 417004 277780
rect 418172 273766 418200 277780
rect 418160 273760 418212 273766
rect 418160 273702 418212 273708
rect 416964 270836 417016 270842
rect 416964 270778 417016 270784
rect 419368 265606 419396 277780
rect 420564 268122 420592 277780
rect 421668 273562 421696 277780
rect 422864 273698 422892 277780
rect 422852 273692 422904 273698
rect 422852 273634 422904 273640
rect 421656 273556 421708 273562
rect 421656 273498 421708 273504
rect 424060 270910 424088 277780
rect 425256 273970 425284 277780
rect 425244 273964 425296 273970
rect 425244 273906 425296 273912
rect 424048 270904 424100 270910
rect 424048 270846 424100 270852
rect 426452 268258 426480 277780
rect 427084 274304 427136 274310
rect 427084 274246 427136 274252
rect 427096 273834 427124 274246
rect 427084 273828 427136 273834
rect 427084 273770 427136 273776
rect 426440 268252 426492 268258
rect 426440 268194 426492 268200
rect 427648 268190 427676 277780
rect 428844 273902 428872 277780
rect 428832 273896 428884 273902
rect 428832 273838 428884 273844
rect 427636 268184 427688 268190
rect 427636 268126 427688 268132
rect 420552 268116 420604 268122
rect 420552 268058 420604 268064
rect 429948 265742 429976 277780
rect 431144 270978 431172 277780
rect 432340 274106 432368 277780
rect 432328 274100 432380 274106
rect 432328 274042 432380 274048
rect 431132 270972 431184 270978
rect 431132 270914 431184 270920
rect 433536 268326 433564 277780
rect 434732 271046 434760 277780
rect 435928 274038 435956 277780
rect 437032 274174 437060 277780
rect 437020 274168 437072 274174
rect 437020 274110 437072 274116
rect 435916 274032 435968 274038
rect 435916 273974 435968 273980
rect 434720 271040 434772 271046
rect 434720 270982 434772 270988
rect 438228 268394 438256 277780
rect 439424 274242 439452 277780
rect 439412 274236 439464 274242
rect 439412 274178 439464 274184
rect 440620 268462 440648 277780
rect 441816 271182 441844 277780
rect 443012 273834 443040 277780
rect 443000 273828 443052 273834
rect 443000 273770 443052 273776
rect 441804 271176 441856 271182
rect 441804 271118 441856 271124
rect 444208 271114 444236 277780
rect 444196 271108 444248 271114
rect 444196 271050 444248 271056
rect 445312 268530 445340 277780
rect 446508 274378 446536 277780
rect 446496 274372 446548 274378
rect 446496 274314 446548 274320
rect 447704 268598 447732 277780
rect 448900 271318 448928 277780
rect 450096 274446 450124 277780
rect 450084 274440 450136 274446
rect 450084 274382 450136 274388
rect 448888 271312 448940 271318
rect 448888 271254 448940 271260
rect 451292 271250 451320 277780
rect 451280 271244 451332 271250
rect 451280 271186 451332 271192
rect 452488 268666 452516 277780
rect 452476 268660 452528 268666
rect 452476 268602 452528 268608
rect 447692 268592 447744 268598
rect 447692 268534 447744 268540
rect 445300 268524 445352 268530
rect 445300 268466 445352 268472
rect 440608 268456 440660 268462
rect 440608 268398 440660 268404
rect 438216 268388 438268 268394
rect 438216 268330 438268 268336
rect 433524 268320 433576 268326
rect 433524 268262 433576 268268
rect 453592 265878 453620 277780
rect 454788 268734 454816 277780
rect 455984 271386 456012 277780
rect 455972 271380 456024 271386
rect 455972 271322 456024 271328
rect 454776 268728 454828 268734
rect 454776 268670 454828 268676
rect 457180 265946 457208 277780
rect 458376 272338 458404 277780
rect 458364 272332 458416 272338
rect 458364 272274 458416 272280
rect 459468 272332 459520 272338
rect 459468 272274 459520 272280
rect 457168 265940 457220 265946
rect 457168 265882 457220 265888
rect 453580 265872 453632 265878
rect 459480 265849 459508 272274
rect 459572 268802 459600 277780
rect 460676 274514 460704 277780
rect 460664 274508 460716 274514
rect 460664 274450 460716 274456
rect 461872 268870 461900 277780
rect 463068 271522 463096 277780
rect 464264 274582 464292 277780
rect 464252 274576 464304 274582
rect 464252 274518 464304 274524
rect 465460 272542 465488 277780
rect 465448 272536 465500 272542
rect 465448 272478 465500 272484
rect 466276 272536 466328 272542
rect 466276 272478 466328 272484
rect 463056 271516 463108 271522
rect 463056 271458 463108 271464
rect 461860 268864 461912 268870
rect 461860 268806 461912 268812
rect 459560 268796 459612 268802
rect 459560 268738 459612 268744
rect 466288 265985 466316 272478
rect 466656 269006 466684 277780
rect 467852 275942 467880 277780
rect 467840 275936 467892 275942
rect 467840 275878 467892 275884
rect 466644 269000 466696 269006
rect 466644 268942 466696 268948
rect 468956 268938 468984 277780
rect 470152 272746 470180 277780
rect 471348 276010 471376 277780
rect 471336 276004 471388 276010
rect 471336 275946 471388 275952
rect 470140 272740 470192 272746
rect 470140 272682 470192 272688
rect 471980 272740 472032 272746
rect 471980 272682 472032 272688
rect 468944 268932 468996 268938
rect 468944 268874 468996 268880
rect 466274 265976 466330 265985
rect 466274 265911 466330 265920
rect 453580 265814 453632 265820
rect 459466 265840 459522 265849
rect 459466 265775 459522 265784
rect 429936 265736 429988 265742
rect 429936 265678 429988 265684
rect 419356 265600 419408 265606
rect 419356 265542 419408 265548
rect 415768 265532 415820 265538
rect 415768 265474 415820 265480
rect 412272 265464 412324 265470
rect 412272 265406 412324 265412
rect 471992 265334 472020 272682
rect 472544 271454 472572 277780
rect 472532 271448 472584 271454
rect 472532 271390 472584 271396
rect 473740 269074 473768 277780
rect 473728 269068 473780 269074
rect 473728 269010 473780 269016
rect 474936 266014 474964 277780
rect 476132 270502 476160 277780
rect 477236 271590 477264 277780
rect 477224 271584 477276 271590
rect 477224 271526 477276 271532
rect 476120 270496 476172 270502
rect 476120 270438 476172 270444
rect 478432 266082 478460 277780
rect 479628 271658 479656 277780
rect 479616 271652 479668 271658
rect 479616 271594 479668 271600
rect 480824 270434 480852 277780
rect 482020 275874 482048 277780
rect 482008 275868 482060 275874
rect 482008 275810 482060 275816
rect 480812 270428 480864 270434
rect 480812 270370 480864 270376
rect 483216 270366 483244 277780
rect 484320 271794 484348 277780
rect 485516 275806 485544 277780
rect 485504 275800 485556 275806
rect 485504 275742 485556 275748
rect 484308 271788 484360 271794
rect 484308 271730 484360 271736
rect 486712 271726 486740 277780
rect 486700 271720 486752 271726
rect 486700 271662 486752 271668
rect 483204 270360 483256 270366
rect 483204 270302 483256 270308
rect 487908 270298 487936 277780
rect 487896 270292 487948 270298
rect 487896 270234 487948 270240
rect 489104 266150 489132 277780
rect 490300 270230 490328 277780
rect 491496 273222 491524 277780
rect 491484 273216 491536 273222
rect 491484 273158 491536 273164
rect 490288 270224 490340 270230
rect 490288 270166 490340 270172
rect 492600 266218 492628 277780
rect 493796 270162 493824 277780
rect 493784 270156 493836 270162
rect 493784 270098 493836 270104
rect 494992 268297 495020 277780
rect 496188 275738 496216 277780
rect 496176 275732 496228 275738
rect 496176 275674 496228 275680
rect 497384 273086 497412 277780
rect 498580 273154 498608 277780
rect 499776 275670 499804 277780
rect 499764 275664 499816 275670
rect 499764 275606 499816 275612
rect 498568 273148 498620 273154
rect 498568 273090 498620 273096
rect 497372 273080 497424 273086
rect 497372 273022 497424 273028
rect 498844 273080 498896 273086
rect 498844 273022 498896 273028
rect 494978 268288 495034 268297
rect 494978 268223 495034 268232
rect 492588 266212 492640 266218
rect 492588 266154 492640 266160
rect 489092 266144 489144 266150
rect 489092 266086 489144 266092
rect 478420 266076 478472 266082
rect 478420 266018 478472 266024
rect 474924 266008 474976 266014
rect 474924 265950 474976 265956
rect 498856 265674 498884 273022
rect 500880 270094 500908 277780
rect 500868 270088 500920 270094
rect 500868 270030 500920 270036
rect 502076 268433 502104 277780
rect 502062 268424 502118 268433
rect 502062 268359 502118 268368
rect 503272 266286 503300 277780
rect 504468 273018 504496 277780
rect 504456 273012 504508 273018
rect 504456 272954 504508 272960
rect 505664 272950 505692 277780
rect 506860 275602 506888 277780
rect 506848 275596 506900 275602
rect 506848 275538 506900 275544
rect 505652 272944 505704 272950
rect 505652 272886 505704 272892
rect 507964 268705 507992 277780
rect 507950 268696 508006 268705
rect 507950 268631 508006 268640
rect 509160 268569 509188 277780
rect 509146 268560 509202 268569
rect 509146 268495 509202 268504
rect 510356 267714 510384 277780
rect 511552 272814 511580 277780
rect 512748 272882 512776 277780
rect 513944 275534 513972 277780
rect 513932 275528 513984 275534
rect 513932 275470 513984 275476
rect 512736 272876 512788 272882
rect 512736 272818 512788 272824
rect 511540 272808 511592 272814
rect 511540 272750 511592 272756
rect 511632 272808 511684 272814
rect 511632 272750 511684 272756
rect 510344 267708 510396 267714
rect 510344 267650 510396 267656
rect 503260 266280 503312 266286
rect 503260 266222 503312 266228
rect 511644 265810 511672 272750
rect 515140 270026 515168 277780
rect 515128 270020 515180 270026
rect 515128 269962 515180 269968
rect 516244 268841 516272 277780
rect 516230 268832 516286 268841
rect 516230 268767 516286 268776
rect 517440 267646 517468 277780
rect 518636 272678 518664 277780
rect 518624 272672 518676 272678
rect 518624 272614 518676 272620
rect 519832 271425 519860 277780
rect 521028 275466 521056 277780
rect 521016 275460 521068 275466
rect 521016 275402 521068 275408
rect 519818 271416 519874 271425
rect 519818 271351 519874 271360
rect 522224 268977 522252 277780
rect 523420 269958 523448 277780
rect 523408 269952 523460 269958
rect 523408 269894 523460 269900
rect 522210 268968 522266 268977
rect 522210 268903 522266 268912
rect 517428 267640 517480 267646
rect 517428 267582 517480 267588
rect 524524 267578 524552 277780
rect 525720 271561 525748 277780
rect 526916 271697 526944 277780
rect 528112 275398 528140 277780
rect 528100 275392 528152 275398
rect 528100 275334 528152 275340
rect 526902 271688 526958 271697
rect 526902 271623 526958 271632
rect 525706 271552 525762 271561
rect 525706 271487 525762 271496
rect 529308 270473 529336 277780
rect 529294 270464 529350 270473
rect 529294 270399 529350 270408
rect 530504 269890 530532 277780
rect 530492 269884 530544 269890
rect 530492 269826 530544 269832
rect 524512 267572 524564 267578
rect 524512 267514 524564 267520
rect 531608 267510 531636 277780
rect 532804 272610 532832 277780
rect 534000 273193 534028 277780
rect 535196 275330 535224 277780
rect 535184 275324 535236 275330
rect 535184 275266 535236 275272
rect 533986 273184 534042 273193
rect 533986 273119 534042 273128
rect 532792 272604 532844 272610
rect 532792 272546 532844 272552
rect 536392 270337 536420 277780
rect 536378 270328 536434 270337
rect 536378 270263 536434 270272
rect 537588 269822 537616 277780
rect 537576 269816 537628 269822
rect 537576 269758 537628 269764
rect 531596 267504 531648 267510
rect 531596 267446 531648 267452
rect 538784 267442 538812 277780
rect 539888 273057 539916 277780
rect 539874 273048 539930 273057
rect 539874 272983 539930 272992
rect 541084 272921 541112 277780
rect 542280 275262 542308 277780
rect 542268 275256 542320 275262
rect 542268 275198 542320 275204
rect 541070 272912 541126 272921
rect 541070 272847 541126 272856
rect 543476 270201 543504 277780
rect 543462 270192 543518 270201
rect 543462 270127 543518 270136
rect 544672 269754 544700 277780
rect 545868 272474 545896 277780
rect 545856 272468 545908 272474
rect 545856 272410 545908 272416
rect 544660 269748 544712 269754
rect 544660 269690 544712 269696
rect 538772 267436 538824 267442
rect 538772 267378 538824 267384
rect 547064 267374 547092 277780
rect 548168 272785 548196 277780
rect 548154 272776 548210 272785
rect 548154 272711 548210 272720
rect 547052 267368 547104 267374
rect 547052 267310 547104 267316
rect 549364 267306 549392 277780
rect 550560 275194 550588 277780
rect 550548 275188 550600 275194
rect 550548 275130 550600 275136
rect 551756 269686 551784 277780
rect 551744 269680 551796 269686
rect 551744 269622 551796 269628
rect 549352 267300 549404 267306
rect 549352 267242 549404 267248
rect 552952 267170 552980 277780
rect 554148 267238 554176 277780
rect 555252 272406 555280 277780
rect 555240 272400 555292 272406
rect 555240 272342 555292 272348
rect 554136 267232 554188 267238
rect 554136 267174 554188 267180
rect 552940 267164 552992 267170
rect 552940 267106 552992 267112
rect 556448 267102 556476 277780
rect 557644 275126 557672 277780
rect 557632 275120 557684 275126
rect 557632 275062 557684 275068
rect 558840 270065 558868 277780
rect 558826 270056 558882 270065
rect 558826 269991 558882 270000
rect 556436 267096 556488 267102
rect 556436 267038 556488 267044
rect 560036 267034 560064 277780
rect 560024 267028 560076 267034
rect 560024 266970 560076 266976
rect 561232 266966 561260 277780
rect 562428 272649 562456 277780
rect 562414 272640 562470 272649
rect 562414 272575 562470 272584
rect 561220 266960 561272 266966
rect 561220 266902 561272 266908
rect 563532 266898 563560 277780
rect 564728 275058 564756 277780
rect 564716 275052 564768 275058
rect 564716 274994 564768 275000
rect 565924 269618 565952 277780
rect 565912 269612 565964 269618
rect 565912 269554 565964 269560
rect 563520 266892 563572 266898
rect 563520 266834 563572 266840
rect 567120 266762 567148 277780
rect 568316 266830 568344 277780
rect 569512 272270 569540 277780
rect 569500 272264 569552 272270
rect 569500 272206 569552 272212
rect 568304 266824 568356 266830
rect 568304 266766 568356 266772
rect 567108 266756 567160 266762
rect 567108 266698 567160 266704
rect 570708 266694 570736 277780
rect 571812 274990 571840 277780
rect 571800 274984 571852 274990
rect 571800 274926 571852 274932
rect 573008 269929 573036 277780
rect 572994 269920 573050 269929
rect 572994 269855 573050 269864
rect 570696 266688 570748 266694
rect 570696 266630 570748 266636
rect 574204 266558 574232 277780
rect 575400 266626 575428 277780
rect 576596 272202 576624 277780
rect 576584 272196 576636 272202
rect 576584 272138 576636 272144
rect 575388 266620 575440 266626
rect 575388 266562 575440 266568
rect 574192 266552 574244 266558
rect 574192 266494 574244 266500
rect 577792 266121 577820 277780
rect 578896 274922 578924 277780
rect 578884 274916 578936 274922
rect 578884 274858 578936 274864
rect 580092 269550 580120 277780
rect 580080 269544 580132 269550
rect 580080 269486 580132 269492
rect 581288 266257 581316 277780
rect 582484 267617 582512 277780
rect 583680 272134 583708 277780
rect 583668 272128 583720 272134
rect 583668 272070 583720 272076
rect 584876 267753 584904 277780
rect 586072 275913 586100 277780
rect 586058 275904 586114 275913
rect 586058 275839 586114 275848
rect 587176 269482 587204 277780
rect 587164 269476 587216 269482
rect 587164 269418 587216 269424
rect 584862 267744 584918 267753
rect 584862 267679 584918 267688
rect 582470 267608 582526 267617
rect 582470 267543 582526 267552
rect 588372 266490 588400 277780
rect 589568 267481 589596 277780
rect 590764 272066 590792 277780
rect 590752 272060 590804 272066
rect 590752 272002 590804 272008
rect 589554 267472 589610 267481
rect 589554 267407 589610 267416
rect 591960 267345 591988 277780
rect 593156 275777 593184 277780
rect 593142 275768 593198 275777
rect 593142 275703 593198 275712
rect 594352 269793 594380 277780
rect 594338 269784 594394 269793
rect 594338 269719 594394 269728
rect 591946 267336 592002 267345
rect 591946 267271 592002 267280
rect 595456 267209 595484 277780
rect 595442 267200 595498 267209
rect 595442 267135 595498 267144
rect 588360 266484 588412 266490
rect 588360 266426 588412 266432
rect 596652 266422 596680 277780
rect 597848 272513 597876 277780
rect 597834 272504 597890 272513
rect 597834 272439 597890 272448
rect 599044 267073 599072 277780
rect 600240 275641 600268 277780
rect 600226 275632 600282 275641
rect 600226 275567 600282 275576
rect 601436 269414 601464 277780
rect 601424 269408 601476 269414
rect 601424 269350 601476 269356
rect 599030 267064 599086 267073
rect 599030 266999 599086 267008
rect 602540 266937 602568 277780
rect 602526 266928 602582 266937
rect 602526 266863 602582 266872
rect 596640 266416 596692 266422
rect 596640 266358 596692 266364
rect 603736 266354 603764 277780
rect 604932 271998 604960 277780
rect 604920 271992 604972 271998
rect 604920 271934 604972 271940
rect 606128 266801 606156 277780
rect 607324 275505 607352 277780
rect 607310 275496 607366 275505
rect 607310 275431 607366 275440
rect 608520 269346 608548 277780
rect 608508 269340 608560 269346
rect 608508 269282 608560 269288
rect 606114 266792 606170 266801
rect 606114 266727 606170 266736
rect 609716 266665 609744 277780
rect 610820 272814 610848 277780
rect 610808 272808 610860 272814
rect 610808 272750 610860 272756
rect 612016 272377 612044 277780
rect 612002 272368 612058 272377
rect 612002 272303 612058 272312
rect 609702 266656 609758 266665
rect 609702 266591 609758 266600
rect 613212 266529 613240 277780
rect 614408 275369 614436 277780
rect 614394 275360 614450 275369
rect 614394 275295 614450 275304
rect 615604 269278 615632 277780
rect 615592 269272 615644 269278
rect 615592 269214 615644 269220
rect 613198 266520 613254 266529
rect 613198 266455 613254 266464
rect 616800 266393 616828 277780
rect 617996 273086 618024 277780
rect 617984 273080 618036 273086
rect 617984 273022 618036 273028
rect 619100 271930 619128 277780
rect 620296 274854 620324 277780
rect 621492 275233 621520 277780
rect 621478 275224 621534 275233
rect 621478 275159 621534 275168
rect 620284 274848 620336 274854
rect 620284 274790 620336 274796
rect 619088 271924 619140 271930
rect 619088 271866 619140 271872
rect 622688 269657 622716 277780
rect 623884 274961 623912 277780
rect 623870 274952 623926 274961
rect 623870 274887 623926 274896
rect 625080 272746 625108 277780
rect 625068 272740 625120 272746
rect 625068 272682 625120 272688
rect 626184 272241 626212 277780
rect 627380 274786 627408 277780
rect 628576 275097 628604 277780
rect 628562 275088 628618 275097
rect 628562 275023 628618 275032
rect 627368 274780 627420 274786
rect 627368 274722 627420 274728
rect 626170 272232 626226 272241
rect 626170 272167 626226 272176
rect 622674 269648 622730 269657
rect 622674 269583 622730 269592
rect 629772 269521 629800 277780
rect 630968 274825 630996 277780
rect 630954 274816 631010 274825
rect 630954 274751 631010 274760
rect 632164 272542 632192 277780
rect 632152 272536 632204 272542
rect 632152 272478 632204 272484
rect 633360 271862 633388 277780
rect 634464 274718 634492 277780
rect 634452 274712 634504 274718
rect 635660 274689 635688 277780
rect 634452 274654 634504 274660
rect 635646 274680 635702 274689
rect 635646 274615 635702 274624
rect 633348 271856 633400 271862
rect 633348 271798 633400 271804
rect 629758 269512 629814 269521
rect 629758 269447 629814 269456
rect 636856 269385 636884 277780
rect 638052 274553 638080 277780
rect 638038 274544 638094 274553
rect 638038 274479 638094 274488
rect 639248 272338 639276 277780
rect 639236 272332 639288 272338
rect 639236 272274 639288 272280
rect 640444 272105 640472 277780
rect 641640 274650 641668 277780
rect 641628 274644 641680 274650
rect 641628 274586 641680 274592
rect 640430 272096 640486 272105
rect 640430 272031 640486 272040
rect 636842 269376 636898 269385
rect 636842 269311 636898 269320
rect 642744 269249 642772 277780
rect 642730 269240 642786 269249
rect 642730 269175 642786 269184
rect 643940 269113 643968 277780
rect 645136 271969 645164 277780
rect 645122 271960 645178 271969
rect 645122 271895 645178 271904
rect 646332 271833 646360 277780
rect 646318 271824 646374 271833
rect 646318 271759 646374 271768
rect 647528 269210 647556 277780
rect 647516 269204 647568 269210
rect 647516 269146 647568 269152
rect 648724 269142 648752 277780
rect 648712 269136 648764 269142
rect 643926 269104 643982 269113
rect 648712 269078 648764 269084
rect 643926 269039 643982 269048
rect 616786 266384 616842 266393
rect 603724 266348 603776 266354
rect 616786 266319 616842 266328
rect 603724 266290 603776 266296
rect 581274 266248 581330 266257
rect 581274 266183 581330 266192
rect 577778 266112 577834 266121
rect 577778 266047 577834 266056
rect 511632 265804 511684 265810
rect 511632 265746 511684 265752
rect 498844 265668 498896 265674
rect 498844 265610 498896 265616
rect 471980 265328 472032 265334
rect 471980 265270 472032 265276
rect 416778 262304 416834 262313
rect 416778 262239 416780 262248
rect 416832 262239 416834 262248
rect 571708 262268 571760 262274
rect 416780 262210 416832 262216
rect 571708 262210 571760 262216
rect 416778 259176 416834 259185
rect 416778 259111 416834 259120
rect 184938 258632 184994 258641
rect 184938 258567 184994 258576
rect 184952 256766 184980 258567
rect 416792 256766 416820 259111
rect 184940 256760 184992 256766
rect 184940 256702 184992 256708
rect 416780 256760 416832 256766
rect 416780 256702 416832 256708
rect 416778 255912 416834 255921
rect 416778 255847 416834 255856
rect 416792 253978 416820 255847
rect 416780 253972 416832 253978
rect 416780 253914 416832 253920
rect 571524 253972 571576 253978
rect 571524 253914 571576 253920
rect 416778 252784 416834 252793
rect 416778 252719 416834 252728
rect 416792 251258 416820 252719
rect 416780 251252 416832 251258
rect 416780 251194 416832 251200
rect 416778 249520 416834 249529
rect 416778 249455 416834 249464
rect 416792 248470 416820 249455
rect 416780 248464 416832 248470
rect 416780 248406 416832 248412
rect 184938 248024 184994 248033
rect 184938 247959 184994 247968
rect 184952 245682 184980 247959
rect 416778 246392 416834 246401
rect 416778 246327 416834 246336
rect 416792 245682 416820 246327
rect 184940 245676 184992 245682
rect 184940 245618 184992 245624
rect 416780 245676 416832 245682
rect 416780 245618 416832 245624
rect 418066 243128 418122 243137
rect 418066 243063 418122 243072
rect 184940 237448 184992 237454
rect 184938 237416 184940 237425
rect 184992 237416 184994 237425
rect 184938 237351 184994 237360
rect 156144 229084 156196 229090
rect 156144 229026 156196 229032
rect 152832 229016 152884 229022
rect 93030 228984 93086 228993
rect 152832 228958 152884 228964
rect 93030 228919 93086 228928
rect 84658 228848 84714 228857
rect 84658 228783 84714 228792
rect 82726 228440 82782 228449
rect 82726 228375 82782 228384
rect 76286 228304 76342 228313
rect 76286 228239 76342 228248
rect 71226 228168 71282 228177
rect 71226 228103 71282 228112
rect 69478 228032 69534 228041
rect 65340 227996 65392 228002
rect 69478 227967 69534 227976
rect 65340 227938 65392 227944
rect 62762 227896 62818 227905
rect 62762 227831 62818 227840
rect 60280 223236 60332 223242
rect 60280 223178 60332 223184
rect 60292 217410 60320 223178
rect 61106 222320 61162 222329
rect 61106 222255 61162 222264
rect 61936 222284 61988 222290
rect 61120 217410 61148 222255
rect 61936 222226 61988 222232
rect 61948 217410 61976 222226
rect 62776 217410 62804 227831
rect 64512 227792 64564 227798
rect 64512 227734 64564 227740
rect 63406 225176 63462 225185
rect 63406 225111 63462 225120
rect 63420 217410 63448 225111
rect 64524 217410 64552 227734
rect 65352 217410 65380 227938
rect 66994 225312 67050 225321
rect 66994 225247 67050 225256
rect 66168 222352 66220 222358
rect 66168 222294 66220 222300
rect 66180 217410 66208 222294
rect 67008 217410 67036 225247
rect 68652 222488 68704 222494
rect 67822 222456 67878 222465
rect 68652 222430 68704 222436
rect 67822 222391 67878 222400
rect 67836 217410 67864 222391
rect 68664 217410 68692 222430
rect 69492 217410 69520 227967
rect 70398 225448 70454 225457
rect 70398 225383 70454 225392
rect 70412 217410 70440 225383
rect 71240 217410 71268 228103
rect 72056 227860 72108 227866
rect 72056 227802 72108 227808
rect 72068 217410 72096 227802
rect 73712 224936 73764 224942
rect 73712 224878 73764 224884
rect 72882 222728 72938 222737
rect 72882 222663 72938 222672
rect 72896 217410 72924 222663
rect 73724 217410 73752 224878
rect 74446 222592 74502 222601
rect 74446 222527 74502 222536
rect 75368 222556 75420 222562
rect 74460 217410 74488 222527
rect 75368 222498 75420 222504
rect 75380 217410 75408 222498
rect 76300 217410 76328 228239
rect 78772 228064 78824 228070
rect 78772 228006 78824 228012
rect 77944 227928 77996 227934
rect 77944 227870 77996 227876
rect 77114 225584 77170 225593
rect 77114 225519 77170 225528
rect 77128 217410 77156 225519
rect 77956 217410 77984 227870
rect 78784 217410 78812 228006
rect 80426 225856 80482 225865
rect 80426 225791 80482 225800
rect 79598 222864 79654 222873
rect 79598 222799 79654 222808
rect 79612 217410 79640 222799
rect 80440 217410 80468 225791
rect 81254 223000 81310 223009
rect 81254 222935 81310 222944
rect 81268 217410 81296 222935
rect 82176 222692 82228 222698
rect 82176 222634 82228 222640
rect 82188 217410 82216 222634
rect 82740 217410 82768 228375
rect 83830 225720 83886 225729
rect 83830 225655 83886 225664
rect 83844 217410 83872 225655
rect 84672 217410 84700 228783
rect 86314 228712 86370 228721
rect 86314 228647 86370 228656
rect 85488 222624 85540 222630
rect 85488 222566 85540 222572
rect 85500 217410 85528 222566
rect 86328 217410 86356 228647
rect 88062 228576 88118 228585
rect 88062 228511 88118 228520
rect 87144 223440 87196 223446
rect 87144 223382 87196 223388
rect 87156 217410 87184 223382
rect 88076 217410 88104 228511
rect 92202 225992 92258 226001
rect 92202 225927 92258 225936
rect 90548 225276 90600 225282
rect 90548 225218 90600 225224
rect 88892 225004 88944 225010
rect 88892 224946 88944 224952
rect 88904 217410 88932 224946
rect 89718 223136 89774 223145
rect 89718 223071 89774 223080
rect 89732 217410 89760 223071
rect 90560 217410 90588 225218
rect 91376 222760 91428 222766
rect 91376 222702 91428 222708
rect 91388 217410 91416 222702
rect 92216 217410 92244 225927
rect 93044 217410 93072 228919
rect 150256 228880 150308 228886
rect 150256 228822 150308 228828
rect 146024 228812 146076 228818
rect 146024 228754 146076 228760
rect 143448 228676 143500 228682
rect 143448 228618 143500 228624
rect 138480 228608 138532 228614
rect 138480 228550 138532 228556
rect 136824 228472 136876 228478
rect 136824 228414 136876 228420
rect 131764 228404 131816 228410
rect 131764 228346 131816 228352
rect 125048 228336 125100 228342
rect 125048 228278 125100 228284
rect 123392 228200 123444 228206
rect 123392 228142 123444 228148
rect 108212 228132 108264 228138
rect 108212 228074 108264 228080
rect 94778 227488 94834 227497
rect 94778 227423 94834 227432
rect 93768 222080 93820 222086
rect 93768 222022 93820 222028
rect 93780 217410 93808 222022
rect 94792 217410 94820 227423
rect 101494 227352 101550 227361
rect 101494 227287 101550 227296
rect 99838 227216 99894 227225
rect 99838 227151 99894 227160
rect 98918 226264 98974 226273
rect 98918 226199 98974 226208
rect 95608 225072 95660 225078
rect 95608 225014 95660 225020
rect 95620 217410 95648 225014
rect 97262 224768 97318 224777
rect 97262 224703 97318 224712
rect 96434 223272 96490 223281
rect 96434 223207 96490 223216
rect 96448 217410 96476 223207
rect 97276 217410 97304 224703
rect 98090 223408 98146 223417
rect 98090 223343 98146 223352
rect 98104 217410 98132 223343
rect 98932 217410 98960 226199
rect 99852 217410 99880 227151
rect 100668 225208 100720 225214
rect 100668 225150 100720 225156
rect 100680 217410 100708 225150
rect 101508 217410 101536 227287
rect 106554 227080 106610 227089
rect 106554 227015 106610 227024
rect 102046 226128 102102 226137
rect 102046 226063 102102 226072
rect 102060 217410 102088 226063
rect 105728 225344 105780 225350
rect 105728 225286 105780 225292
rect 103980 225140 104032 225146
rect 103980 225082 104032 225088
rect 103150 222048 103206 222057
rect 103150 221983 103206 221992
rect 103164 217410 103192 221983
rect 103992 217410 104020 225082
rect 104806 223544 104862 223553
rect 104806 223479 104862 223488
rect 104820 217410 104848 223479
rect 105740 217410 105768 225286
rect 106568 217410 106596 227015
rect 107384 225412 107436 225418
rect 107384 225354 107436 225360
rect 107396 217410 107424 225354
rect 108224 217410 108252 228074
rect 113086 226944 113142 226953
rect 113086 226879 113142 226888
rect 109038 224632 109094 224641
rect 109038 224567 109094 224576
rect 109052 217410 109080 224567
rect 112442 224496 112498 224505
rect 112442 224431 112498 224440
rect 110694 224224 110750 224233
rect 110694 224159 110750 224168
rect 109866 221912 109922 221921
rect 109866 221847 109922 221856
rect 109880 217410 109908 221847
rect 110708 217410 110736 224159
rect 111614 221776 111670 221785
rect 111614 221711 111670 221720
rect 111628 217410 111656 221711
rect 112456 217410 112484 224431
rect 113100 217410 113128 226879
rect 114926 226808 114982 226817
rect 114926 226743 114982 226752
rect 114100 225548 114152 225554
rect 114100 225490 114152 225496
rect 114112 217410 114140 225490
rect 114940 217410 114968 226743
rect 119160 225684 119212 225690
rect 119160 225626 119212 225632
rect 117504 225480 117556 225486
rect 117504 225422 117556 225428
rect 115754 224360 115810 224369
rect 115754 224295 115810 224304
rect 115768 217410 115796 224295
rect 116584 222828 116636 222834
rect 116584 222770 116636 222776
rect 116596 217410 116624 222770
rect 117516 217410 117544 225422
rect 118330 221504 118386 221513
rect 118330 221439 118386 221448
rect 118344 217410 118372 221439
rect 119172 217410 119200 225626
rect 120814 224088 120870 224097
rect 120814 224023 120870 224032
rect 119988 222896 120040 222902
rect 119988 222838 120040 222844
rect 120000 217410 120028 222838
rect 120828 217410 120856 224023
rect 121366 221640 121422 221649
rect 121366 221575 121422 221584
rect 121380 217410 121408 221575
rect 122472 219904 122524 219910
rect 122472 219846 122524 219852
rect 122484 217410 122512 219846
rect 123404 217410 123432 228142
rect 124128 225616 124180 225622
rect 124128 225558 124180 225564
rect 124140 217410 124168 225558
rect 125060 217410 125088 228278
rect 130108 228268 130160 228274
rect 130108 228210 130160 228216
rect 127532 225752 127584 225758
rect 127532 225694 127584 225700
rect 126704 222964 126756 222970
rect 126704 222906 126756 222912
rect 125876 219972 125928 219978
rect 125876 219914 125928 219920
rect 125888 217410 125916 219914
rect 126716 217410 126744 222906
rect 127544 217410 127572 225694
rect 128360 223032 128412 223038
rect 128360 222974 128412 222980
rect 128372 217410 128400 222974
rect 129280 220040 129332 220046
rect 129280 219982 129332 219988
rect 129292 217410 129320 219982
rect 130120 217410 130148 228210
rect 130936 225820 130988 225826
rect 130936 225762 130988 225768
rect 130948 217410 130976 225762
rect 131776 217410 131804 228346
rect 134248 225888 134300 225894
rect 134248 225830 134300 225836
rect 133420 223100 133472 223106
rect 133420 223042 133472 223048
rect 132408 220108 132460 220114
rect 132408 220050 132460 220056
rect 132420 217410 132448 220050
rect 133432 217410 133460 223042
rect 134260 217410 134288 225830
rect 135168 223168 135220 223174
rect 135168 223110 135220 223116
rect 135180 217410 135208 223110
rect 135996 220176 136048 220182
rect 135996 220118 136048 220124
rect 136008 217410 136036 220118
rect 136836 217410 136864 228414
rect 137652 225956 137704 225962
rect 137652 225898 137704 225904
rect 137664 217410 137692 225898
rect 138492 217410 138520 228550
rect 141056 226024 141108 226030
rect 141056 225966 141108 225972
rect 139308 224120 139360 224126
rect 139308 224062 139360 224068
rect 139320 223242 139348 224062
rect 140136 223576 140188 223582
rect 140136 223518 140188 223524
rect 139308 223236 139360 223242
rect 139308 223178 139360 223184
rect 139308 220312 139360 220318
rect 139308 220254 139360 220260
rect 139320 217410 139348 220254
rect 140148 217410 140176 223518
rect 141068 217410 141096 225966
rect 141884 223236 141936 223242
rect 141884 223178 141936 223184
rect 141896 217410 141924 223178
rect 142712 220244 142764 220250
rect 142712 220186 142764 220192
rect 142724 217410 142752 220186
rect 143460 217410 143488 228618
rect 145196 228540 145248 228546
rect 145196 228482 145248 228488
rect 144368 226160 144420 226166
rect 144368 226102 144420 226108
rect 144380 217410 144408 226102
rect 145208 217410 145236 228482
rect 146036 217410 146064 228754
rect 147772 226092 147824 226098
rect 147772 226034 147824 226040
rect 146944 223372 146996 223378
rect 146944 223314 146996 223320
rect 146956 217410 146984 223314
rect 147784 217410 147812 226034
rect 148600 223304 148652 223310
rect 148600 223246 148652 223252
rect 148612 217410 148640 223246
rect 149428 221196 149480 221202
rect 149428 221138 149480 221144
rect 149440 217410 149468 221138
rect 150268 217410 150296 228822
rect 151728 228744 151780 228750
rect 151728 228686 151780 228692
rect 151084 226296 151136 226302
rect 151084 226238 151136 226244
rect 151096 217410 151124 226238
rect 151740 217410 151768 228686
rect 152844 217410 152872 228958
rect 154488 226228 154540 226234
rect 154488 226170 154540 226176
rect 153660 223508 153712 223514
rect 153660 223450 153712 223456
rect 153672 217410 153700 223450
rect 154500 217410 154528 226170
rect 155868 224052 155920 224058
rect 155868 223994 155920 224000
rect 155316 222148 155368 222154
rect 155316 222090 155368 222096
rect 155328 217410 155356 222090
rect 155880 222086 155908 223994
rect 155868 222080 155920 222086
rect 155868 222022 155920 222028
rect 156156 217410 156184 229026
rect 156972 228948 157024 228954
rect 156972 228890 157024 228896
rect 156984 217410 157012 228890
rect 158720 227656 158772 227662
rect 158720 227598 158772 227604
rect 157800 224800 157852 224806
rect 157800 224742 157852 224748
rect 157812 217410 157840 224742
rect 158732 217410 158760 227598
rect 165436 227588 165488 227594
rect 165436 227530 165488 227536
rect 162768 227520 162820 227526
rect 162768 227462 162820 227468
rect 161204 224868 161256 224874
rect 161204 224810 161256 224816
rect 160376 222012 160428 222018
rect 160376 221954 160428 221960
rect 159548 221536 159600 221542
rect 159548 221478 159600 221484
rect 159560 217410 159588 221478
rect 160388 217410 160416 221954
rect 161216 217410 161244 224810
rect 162032 220924 162084 220930
rect 162032 220866 162084 220872
rect 162044 217410 162072 220866
rect 162780 217410 162808 227462
rect 163688 227452 163740 227458
rect 163688 227394 163740 227400
rect 163700 217410 163728 227394
rect 164608 224664 164660 224670
rect 164608 224606 164660 224612
rect 164620 217410 164648 224606
rect 165448 217410 165476 227530
rect 167092 227384 167144 227390
rect 167092 227326 167144 227332
rect 166264 221468 166316 221474
rect 166264 221410 166316 221416
rect 166276 217410 166304 221410
rect 167104 217410 167132 227326
rect 172152 227316 172204 227322
rect 172152 227258 172204 227264
rect 169576 227248 169628 227254
rect 169576 227190 169628 227196
rect 167920 224732 167972 224738
rect 167920 224674 167972 224680
rect 167932 217410 167960 224674
rect 168748 221876 168800 221882
rect 168748 221818 168800 221824
rect 168760 217410 168788 221818
rect 169588 217410 169616 227190
rect 170956 224596 171008 224602
rect 170956 224538 171008 224544
rect 170496 221944 170548 221950
rect 170496 221886 170548 221892
rect 170508 217410 170536 221886
rect 59984 217382 60320 217410
rect 60812 217382 61148 217410
rect 61640 217382 61976 217410
rect 62468 217382 62804 217410
rect 63296 217382 63448 217410
rect 64216 217382 64552 217410
rect 65044 217382 65380 217410
rect 65872 217382 66208 217410
rect 66700 217382 67036 217410
rect 67528 217382 67864 217410
rect 68356 217382 68692 217410
rect 69184 217382 69520 217410
rect 70104 217382 70440 217410
rect 70932 217382 71268 217410
rect 71760 217382 72096 217410
rect 72588 217382 72924 217410
rect 73416 217382 73752 217410
rect 74244 217382 74488 217410
rect 75072 217382 75408 217410
rect 75992 217382 76328 217410
rect 76820 217382 77156 217410
rect 77648 217382 77984 217410
rect 78476 217382 78812 217410
rect 79304 217382 79640 217410
rect 80132 217382 80468 217410
rect 80960 217382 81296 217410
rect 81880 217382 82216 217410
rect 82708 217382 82768 217410
rect 83536 217382 83872 217410
rect 84364 217382 84700 217410
rect 85192 217382 85528 217410
rect 86020 217382 86356 217410
rect 86848 217382 87184 217410
rect 87768 217382 88104 217410
rect 88596 217382 88932 217410
rect 89424 217382 89760 217410
rect 90252 217382 90588 217410
rect 91080 217382 91416 217410
rect 91908 217382 92244 217410
rect 92736 217382 93072 217410
rect 93656 217382 93808 217410
rect 94484 217382 94820 217410
rect 95312 217382 95648 217410
rect 96140 217382 96476 217410
rect 96968 217382 97304 217410
rect 97796 217382 98132 217410
rect 98624 217382 98960 217410
rect 99544 217382 99880 217410
rect 100372 217382 100708 217410
rect 101200 217382 101536 217410
rect 102028 217382 102088 217410
rect 102856 217382 103192 217410
rect 103684 217382 104020 217410
rect 104512 217382 104848 217410
rect 105432 217382 105768 217410
rect 106260 217382 106596 217410
rect 107088 217382 107424 217410
rect 107916 217382 108252 217410
rect 108744 217382 109080 217410
rect 109572 217382 109908 217410
rect 110400 217382 110736 217410
rect 111320 217382 111656 217410
rect 112148 217382 112484 217410
rect 112976 217382 113128 217410
rect 113804 217382 114140 217410
rect 114632 217382 114968 217410
rect 115460 217382 115796 217410
rect 116288 217382 116624 217410
rect 117208 217382 117544 217410
rect 118036 217382 118372 217410
rect 118864 217382 119200 217410
rect 119692 217382 120028 217410
rect 120520 217382 120856 217410
rect 121348 217382 121408 217410
rect 122176 217382 122512 217410
rect 123096 217382 123432 217410
rect 123924 217382 124168 217410
rect 124752 217382 125088 217410
rect 125580 217382 125916 217410
rect 126408 217382 126744 217410
rect 127236 217382 127572 217410
rect 128064 217382 128400 217410
rect 128984 217382 129320 217410
rect 129812 217382 130148 217410
rect 130640 217382 130976 217410
rect 131468 217382 131804 217410
rect 132296 217382 132448 217410
rect 133124 217382 133460 217410
rect 133952 217382 134288 217410
rect 134872 217382 135208 217410
rect 135700 217382 136036 217410
rect 136528 217382 136864 217410
rect 137356 217382 137692 217410
rect 138184 217382 138520 217410
rect 139012 217382 139348 217410
rect 139840 217382 140176 217410
rect 140760 217382 141096 217410
rect 141588 217382 141924 217410
rect 142416 217382 142752 217410
rect 143244 217382 143488 217410
rect 144072 217382 144408 217410
rect 144900 217382 145236 217410
rect 145728 217382 146064 217410
rect 146648 217382 146984 217410
rect 147476 217382 147812 217410
rect 148304 217382 148640 217410
rect 149132 217382 149468 217410
rect 149960 217382 150296 217410
rect 150788 217382 151124 217410
rect 151616 217382 151768 217410
rect 152536 217382 152872 217410
rect 153364 217382 153700 217410
rect 154192 217382 154528 217410
rect 155020 217382 155356 217410
rect 155848 217382 156184 217410
rect 156676 217382 157012 217410
rect 157504 217382 157840 217410
rect 158424 217382 158760 217410
rect 159252 217382 159588 217410
rect 160080 217382 160416 217410
rect 160908 217382 161244 217410
rect 161736 217382 162072 217410
rect 162564 217382 162808 217410
rect 163392 217382 163728 217410
rect 164312 217382 164648 217410
rect 165140 217382 165476 217410
rect 165968 217382 166304 217410
rect 166796 217382 167132 217410
rect 167624 217382 167960 217410
rect 168452 217382 168788 217410
rect 169280 217382 169616 217410
rect 170200 217382 170536 217410
rect 170968 217410 170996 224538
rect 171048 223712 171100 223718
rect 171048 223654 171100 223660
rect 171060 223446 171088 223654
rect 171048 223440 171100 223446
rect 171048 223382 171100 223388
rect 172164 217410 172192 227258
rect 173624 227180 173676 227186
rect 173624 227122 173676 227128
rect 172980 221332 173032 221338
rect 172980 221274 173032 221280
rect 172992 217410 173020 221274
rect 173636 217410 173664 227122
rect 178868 227112 178920 227118
rect 178868 227054 178920 227060
rect 176384 227044 176436 227050
rect 176384 226986 176436 226992
rect 174636 224528 174688 224534
rect 174636 224470 174688 224476
rect 174648 217410 174676 224470
rect 175464 221808 175516 221814
rect 175464 221750 175516 221756
rect 175476 217410 175504 221750
rect 176396 217410 176424 226986
rect 178040 224392 178092 224398
rect 178040 224334 178092 224340
rect 177212 223440 177264 223446
rect 177212 223382 177264 223388
rect 177224 217410 177252 223382
rect 178052 217410 178080 224334
rect 178880 217410 178908 227054
rect 180524 226976 180576 226982
rect 180524 226918 180576 226924
rect 179696 221128 179748 221134
rect 179696 221070 179748 221076
rect 179708 217410 179736 221070
rect 180536 217410 180564 226918
rect 190368 226908 190420 226914
rect 190368 226850 190420 226856
rect 185584 226840 185636 226846
rect 185584 226782 185636 226788
rect 181352 224460 181404 224466
rect 181352 224402 181404 224408
rect 181364 217410 181392 224402
rect 184756 224324 184808 224330
rect 184756 224266 184808 224272
rect 182180 223644 182232 223650
rect 182180 223586 182232 223592
rect 182192 222426 182220 223586
rect 182180 222420 182232 222426
rect 182180 222362 182232 222368
rect 182088 221740 182140 221746
rect 182088 221682 182140 221688
rect 182100 217410 182128 221682
rect 183928 221672 183980 221678
rect 183928 221614 183980 221620
rect 183100 221604 183152 221610
rect 183100 221546 183152 221552
rect 183112 217410 183140 221546
rect 183940 217410 183968 221614
rect 184768 217410 184796 224266
rect 185596 217410 185624 226782
rect 186412 226772 186464 226778
rect 186412 226714 186464 226720
rect 186424 217410 186452 226714
rect 188160 224256 188212 224262
rect 188160 224198 188212 224204
rect 187240 221400 187292 221406
rect 187240 221342 187292 221348
rect 187252 217410 187280 221342
rect 188172 217410 188200 224198
rect 189724 223848 189776 223854
rect 189724 223790 189776 223796
rect 188988 222420 189040 222426
rect 188988 222362 189040 222368
rect 189000 217410 189028 222362
rect 189736 221202 189764 223790
rect 189724 221196 189776 221202
rect 189724 221138 189776 221144
rect 189816 221196 189868 221202
rect 189816 221138 189868 221144
rect 189828 217410 189856 221138
rect 190380 217410 190408 226850
rect 191472 224188 191524 224194
rect 191472 224130 191524 224136
rect 191484 217410 191512 224130
rect 192312 223650 192340 231676
rect 192588 225049 192616 231676
rect 192956 227730 192984 231676
rect 192944 227724 192996 227730
rect 192944 227666 192996 227672
rect 193036 227724 193088 227730
rect 193036 227666 193088 227672
rect 192944 226704 192996 226710
rect 192944 226646 192996 226652
rect 192574 225040 192630 225049
rect 192574 224975 192630 224984
rect 192300 223644 192352 223650
rect 192300 223586 192352 223592
rect 192300 221264 192352 221270
rect 192300 221206 192352 221212
rect 192312 217410 192340 221206
rect 192956 217410 192984 226646
rect 193048 221270 193076 227666
rect 193324 222193 193352 231676
rect 193692 224913 193720 231676
rect 193784 231662 194074 231690
rect 193678 224904 193734 224913
rect 193678 224839 193734 224848
rect 193310 222184 193366 222193
rect 193310 222119 193366 222128
rect 193036 221264 193088 221270
rect 193036 221206 193088 221212
rect 193784 219842 193812 231662
rect 194428 227633 194456 231676
rect 194796 227769 194824 231676
rect 194888 231662 195178 231690
rect 194782 227760 194838 227769
rect 194782 227695 194838 227704
rect 194414 227624 194470 227633
rect 194414 227559 194470 227568
rect 194888 224126 194916 231662
rect 194876 224120 194928 224126
rect 194876 224062 194928 224068
rect 194968 224120 195020 224126
rect 194968 224062 195020 224068
rect 194048 220856 194100 220862
rect 194048 220798 194100 220804
rect 193772 219836 193824 219842
rect 193772 219778 193824 219784
rect 194060 217410 194088 220798
rect 194980 217410 195008 224062
rect 195440 222290 195468 231676
rect 195428 222284 195480 222290
rect 195428 222226 195480 222232
rect 195704 222284 195756 222290
rect 195704 222226 195756 222232
rect 195716 217410 195744 222226
rect 195808 222222 195836 231676
rect 196176 222329 196204 231676
rect 196544 225185 196572 231676
rect 196912 228002 196940 231676
rect 196900 227996 196952 228002
rect 196900 227938 196952 227944
rect 197280 227905 197308 231676
rect 197266 227896 197322 227905
rect 197266 227831 197322 227840
rect 197648 227798 197676 231676
rect 197636 227792 197688 227798
rect 197636 227734 197688 227740
rect 197728 227792 197780 227798
rect 197728 227734 197780 227740
rect 197740 226334 197768 227734
rect 197464 226306 197768 226334
rect 197912 226364 197964 226370
rect 197912 226306 197964 226312
rect 196530 225176 196586 225185
rect 196530 225111 196586 225120
rect 196162 222320 196218 222329
rect 196162 222255 196218 222264
rect 195796 222216 195848 222222
rect 195796 222158 195848 222164
rect 196532 220992 196584 220998
rect 196532 220934 196584 220940
rect 196544 217410 196572 220934
rect 197464 217410 197492 226306
rect 197924 225282 197952 226306
rect 198016 225321 198044 231676
rect 198002 225312 198058 225321
rect 197912 225276 197964 225282
rect 198002 225247 198058 225256
rect 198188 225276 198240 225282
rect 197912 225218 197964 225224
rect 198188 225218 198240 225224
rect 198200 217410 198228 225218
rect 198292 222494 198320 231676
rect 198280 222488 198332 222494
rect 198280 222430 198332 222436
rect 198660 222358 198688 231676
rect 198752 231662 199042 231690
rect 198752 222465 198780 231662
rect 199016 227996 199068 228002
rect 199016 227938 199068 227944
rect 198738 222456 198794 222465
rect 198738 222391 198794 222400
rect 198648 222352 198700 222358
rect 198648 222294 198700 222300
rect 199028 217410 199056 227938
rect 199396 225457 199424 231676
rect 199764 227866 199792 231676
rect 200132 228041 200160 231676
rect 200500 228177 200528 231676
rect 200486 228168 200542 228177
rect 200486 228103 200542 228112
rect 200118 228032 200174 228041
rect 200118 227967 200174 227976
rect 199752 227860 199804 227866
rect 199752 227802 199804 227808
rect 199382 225448 199438 225457
rect 199382 225383 199438 225392
rect 200868 224942 200896 231676
rect 200856 224936 200908 224942
rect 200856 224878 200908 224884
rect 201144 222562 201172 231676
rect 201408 224936 201460 224942
rect 201408 224878 201460 224884
rect 201132 222556 201184 222562
rect 201132 222498 201184 222504
rect 200764 222352 200816 222358
rect 200764 222294 200816 222300
rect 199936 221196 199988 221202
rect 199936 221138 199988 221144
rect 199948 217410 199976 221138
rect 200776 217410 200804 222294
rect 201420 217410 201448 224878
rect 201512 222737 201540 231676
rect 201498 222728 201554 222737
rect 201498 222663 201554 222672
rect 201880 222601 201908 231676
rect 202248 225593 202276 231676
rect 202616 228070 202644 231676
rect 202984 228313 203012 231676
rect 203076 231662 203366 231690
rect 202970 228304 203026 228313
rect 202970 228239 203026 228248
rect 202604 228064 202656 228070
rect 202604 228006 202656 228012
rect 203076 227934 203104 231662
rect 203064 227928 203116 227934
rect 203064 227870 203116 227876
rect 203248 227928 203300 227934
rect 203248 227870 203300 227876
rect 202234 225584 202290 225593
rect 202234 225519 202290 225528
rect 201866 222592 201922 222601
rect 201866 222527 201922 222536
rect 202420 222488 202472 222494
rect 202420 222430 202472 222436
rect 202432 217410 202460 222430
rect 203260 217410 203288 227870
rect 203720 225865 203748 231676
rect 203706 225856 203762 225865
rect 203706 225791 203762 225800
rect 203996 222698 204024 231676
rect 204272 231662 204378 231690
rect 204076 227860 204128 227866
rect 204076 227802 204128 227808
rect 203984 222692 204036 222698
rect 203984 222634 204036 222640
rect 204088 217410 204116 227802
rect 204272 226334 204300 231662
rect 204272 226306 204392 226334
rect 204260 223916 204312 223922
rect 204260 223858 204312 223864
rect 204272 220998 204300 223858
rect 204364 222873 204392 226306
rect 204732 223009 204760 231676
rect 205100 225729 205128 231676
rect 205086 225720 205142 225729
rect 205086 225655 205142 225664
rect 204904 223984 204956 223990
rect 204904 223926 204956 223932
rect 204718 223000 204774 223009
rect 204718 222935 204774 222944
rect 204350 222864 204406 222873
rect 204350 222799 204406 222808
rect 204260 220992 204312 220998
rect 204260 220934 204312 220940
rect 204916 217410 204944 223926
rect 205468 222630 205496 231676
rect 205836 228449 205864 231676
rect 206204 228857 206232 231676
rect 206190 228848 206246 228857
rect 206190 228783 206246 228792
rect 205822 228440 205878 228449
rect 205822 228375 205878 228384
rect 206572 223718 206600 231676
rect 206848 225010 206876 231676
rect 207216 228721 207244 231676
rect 207202 228712 207258 228721
rect 207202 228647 207258 228656
rect 207584 228585 207612 231676
rect 207570 228576 207626 228585
rect 207570 228511 207626 228520
rect 207952 226370 207980 231676
rect 207940 226364 207992 226370
rect 207940 226306 207992 226312
rect 208320 226001 208348 231676
rect 208306 225992 208362 226001
rect 208306 225927 208362 225936
rect 206836 225004 206888 225010
rect 206836 224946 206888 224952
rect 208308 225004 208360 225010
rect 208308 224946 208360 224952
rect 206560 223712 206612 223718
rect 206560 223654 206612 223660
rect 205456 222624 205508 222630
rect 205456 222566 205508 222572
rect 205824 222556 205876 222562
rect 205824 222498 205876 222504
rect 205836 217410 205864 222498
rect 207480 222216 207532 222222
rect 207480 222158 207532 222164
rect 206652 221060 206704 221066
rect 206652 221002 206704 221008
rect 206664 217410 206692 221002
rect 207492 217410 207520 222158
rect 208320 217410 208348 224946
rect 208688 223145 208716 231676
rect 208674 223136 208730 223145
rect 208674 223071 208730 223080
rect 209056 222766 209084 231676
rect 209424 223786 209452 231676
rect 209516 231662 209714 231690
rect 209516 225078 209544 231662
rect 210068 228993 210096 231676
rect 210054 228984 210110 228993
rect 210054 228919 210110 228928
rect 209688 228064 209740 228070
rect 209688 228006 209740 228012
rect 209504 225072 209556 225078
rect 209504 225014 209556 225020
rect 209596 224052 209648 224058
rect 209596 223994 209648 224000
rect 209412 223780 209464 223786
rect 209412 223722 209464 223728
rect 209044 222760 209096 222766
rect 209044 222702 209096 222708
rect 209136 222624 209188 222630
rect 209136 222566 209188 222572
rect 209148 217410 209176 222566
rect 209608 221542 209636 223994
rect 209596 221536 209648 221542
rect 209596 221478 209648 221484
rect 209700 217410 209728 228006
rect 210436 227497 210464 231676
rect 210528 231662 210818 231690
rect 210422 227488 210478 227497
rect 210422 227423 210478 227432
rect 210528 224777 210556 231662
rect 210790 227760 210846 227769
rect 210790 227695 210846 227704
rect 210514 224768 210570 224777
rect 210514 224703 210570 224712
rect 210804 217410 210832 227695
rect 211172 226273 211200 231676
rect 211158 226264 211214 226273
rect 211158 226199 211214 226208
rect 211540 223281 211568 231676
rect 211712 225072 211764 225078
rect 211712 225014 211764 225020
rect 211526 223272 211582 223281
rect 211526 223207 211582 223216
rect 211724 217410 211752 225014
rect 211908 223417 211936 231676
rect 212276 225214 212304 231676
rect 212354 227624 212410 227633
rect 212354 227559 212410 227568
rect 212264 225208 212316 225214
rect 212264 225150 212316 225156
rect 211894 223408 211950 223417
rect 211894 223343 211950 223352
rect 212368 217410 212396 227559
rect 212552 226137 212580 231676
rect 212920 227225 212948 231676
rect 213288 227361 213316 231676
rect 213274 227352 213330 227361
rect 213274 227287 213330 227296
rect 212906 227216 212962 227225
rect 212906 227151 212962 227160
rect 212538 226128 212594 226137
rect 212538 226063 212594 226072
rect 213656 225146 213684 231676
rect 214024 225350 214052 231676
rect 214012 225344 214064 225350
rect 214012 225286 214064 225292
rect 213644 225140 213696 225146
rect 213644 225082 213696 225088
rect 213092 223780 213144 223786
rect 213092 223722 213144 223728
rect 213104 221338 213132 223722
rect 214392 222057 214420 231676
rect 214484 231662 214774 231690
rect 214484 223553 214512 231662
rect 215128 225418 215156 231676
rect 215116 225412 215168 225418
rect 215116 225354 215168 225360
rect 215024 225140 215076 225146
rect 215024 225082 215076 225088
rect 214470 223544 214526 223553
rect 214470 223479 214526 223488
rect 214378 222048 214434 222057
rect 214378 221983 214434 221992
rect 214196 221536 214248 221542
rect 214196 221478 214248 221484
rect 213092 221332 213144 221338
rect 213092 221274 213144 221280
rect 213368 220992 213420 220998
rect 213368 220934 213420 220940
rect 213380 217410 213408 220934
rect 214208 217410 214236 221478
rect 215036 217410 215064 225082
rect 215404 224641 215432 231676
rect 215772 227089 215800 231676
rect 216140 228138 216168 231676
rect 216128 228132 216180 228138
rect 216128 228074 216180 228080
rect 215758 227080 215814 227089
rect 215758 227015 215814 227024
rect 215390 224632 215446 224641
rect 215390 224567 215446 224576
rect 216508 224233 216536 231676
rect 216680 228132 216732 228138
rect 216680 228074 216732 228080
rect 216494 224224 216550 224233
rect 216494 224159 216550 224168
rect 215208 223712 215260 223718
rect 215208 223654 215260 223660
rect 215220 221474 215248 223654
rect 215852 222692 215904 222698
rect 215852 222634 215904 222640
rect 215208 221468 215260 221474
rect 215208 221410 215260 221416
rect 215864 217410 215892 222634
rect 216692 217410 216720 228074
rect 216876 224505 216904 231676
rect 216862 224496 216918 224505
rect 216862 224431 216918 224440
rect 217244 221921 217272 231676
rect 217336 231662 217626 231690
rect 217230 221912 217286 221921
rect 217230 221847 217286 221856
rect 217336 221785 217364 231662
rect 217598 227896 217654 227905
rect 217598 227831 217654 227840
rect 217322 221776 217378 221785
rect 217322 221711 217378 221720
rect 217612 217410 217640 227831
rect 217980 225554 218008 231676
rect 217968 225548 218020 225554
rect 217968 225490 218020 225496
rect 218060 225548 218112 225554
rect 218060 225490 218112 225496
rect 218072 225434 218100 225490
rect 217980 225406 218100 225434
rect 217980 221134 218008 225406
rect 218256 224369 218284 231676
rect 218624 226953 218652 231676
rect 218610 226944 218666 226953
rect 218610 226879 218666 226888
rect 218992 226817 219020 231676
rect 219254 228032 219310 228041
rect 219254 227967 219310 227976
rect 218978 226808 219034 226817
rect 218978 226743 219034 226752
rect 218428 225412 218480 225418
rect 218428 225354 218480 225360
rect 218242 224360 218298 224369
rect 218242 224295 218298 224304
rect 217968 221128 218020 221134
rect 217968 221070 218020 221076
rect 218440 217410 218468 225354
rect 219268 217410 219296 227967
rect 219360 225486 219388 231676
rect 219728 225690 219756 231676
rect 219716 225684 219768 225690
rect 219716 225626 219768 225632
rect 219348 225480 219400 225486
rect 219348 225422 219400 225428
rect 220096 222834 220124 231676
rect 220084 222828 220136 222834
rect 220084 222770 220136 222776
rect 220464 221513 220492 231676
rect 220726 228168 220782 228177
rect 220726 228103 220782 228112
rect 220450 221504 220506 221513
rect 220084 221468 220136 221474
rect 220450 221439 220506 221448
rect 220084 221410 220136 221416
rect 220096 217410 220124 221410
rect 220740 217410 220768 228103
rect 220832 224097 220860 231676
rect 220818 224088 220874 224097
rect 220818 224023 220874 224032
rect 221108 219910 221136 231676
rect 221476 222902 221504 231676
rect 221740 225344 221792 225350
rect 221740 225286 221792 225292
rect 221464 222896 221516 222902
rect 221464 222838 221516 222844
rect 221096 219904 221148 219910
rect 221096 219846 221148 219852
rect 221752 217410 221780 225286
rect 221844 221649 221872 231676
rect 222212 225622 222240 231676
rect 222304 231662 222594 231690
rect 222200 225616 222252 225622
rect 222200 225558 222252 225564
rect 221830 221640 221886 221649
rect 221830 221575 221886 221584
rect 222304 219978 222332 231662
rect 222948 228206 222976 231676
rect 223316 228342 223344 231676
rect 223304 228336 223356 228342
rect 223304 228278 223356 228284
rect 223488 228336 223540 228342
rect 223488 228278 223540 228284
rect 222936 228200 222988 228206
rect 222936 228142 222988 228148
rect 222568 222828 222620 222834
rect 222568 222770 222620 222776
rect 222292 219972 222344 219978
rect 222292 219914 222344 219920
rect 222580 217410 222608 222770
rect 223500 217410 223528 228278
rect 223684 225758 223712 231676
rect 223672 225752 223724 225758
rect 223672 225694 223724 225700
rect 223960 220046 223988 231676
rect 224052 231662 224342 231690
rect 224052 222970 224080 231662
rect 224696 223038 224724 231676
rect 225064 225826 225092 231676
rect 225052 225820 225104 225826
rect 225052 225762 225104 225768
rect 225144 225208 225196 225214
rect 225144 225150 225196 225156
rect 224684 223032 224736 223038
rect 224684 222974 224736 222980
rect 224040 222964 224092 222970
rect 224040 222906 224092 222912
rect 224316 222896 224368 222902
rect 224316 222838 224368 222844
rect 223948 220040 224000 220046
rect 223948 219982 224000 219988
rect 224328 217410 224356 222838
rect 225156 217410 225184 225150
rect 225432 220114 225460 231676
rect 225800 228274 225828 231676
rect 226168 228410 226196 231676
rect 226156 228404 226208 228410
rect 226156 228346 226208 228352
rect 225970 228304 226026 228313
rect 225788 228268 225840 228274
rect 225970 228239 226026 228248
rect 225788 228210 225840 228216
rect 225420 220108 225472 220114
rect 225420 220050 225472 220056
rect 225984 217410 226012 228239
rect 226536 225894 226564 231676
rect 226628 231662 226826 231690
rect 226524 225888 226576 225894
rect 226524 225830 226576 225836
rect 226628 220182 226656 231662
rect 227180 223106 227208 231676
rect 227548 223174 227576 231676
rect 227628 228404 227680 228410
rect 227628 228346 227680 228352
rect 227536 223168 227588 223174
rect 227536 223110 227588 223116
rect 227168 223100 227220 223106
rect 227168 223042 227220 223048
rect 226800 221060 226852 221066
rect 226800 221002 226852 221008
rect 226616 220176 226668 220182
rect 226616 220118 226668 220124
rect 226812 217410 226840 221002
rect 227640 217410 227668 228346
rect 227916 225962 227944 231676
rect 227904 225956 227956 225962
rect 227904 225898 227956 225904
rect 228284 220318 228312 231676
rect 228652 228478 228680 231676
rect 229020 228614 229048 231676
rect 229112 231662 229402 231690
rect 229008 228608 229060 228614
rect 229008 228550 229060 228556
rect 228640 228472 228692 228478
rect 228640 228414 228692 228420
rect 229112 226030 229140 231662
rect 229376 228268 229428 228274
rect 229376 228210 229428 228216
rect 229100 226024 229152 226030
rect 229100 225966 229152 225972
rect 228456 225480 228508 225486
rect 228456 225422 228508 225428
rect 228272 220312 228324 220318
rect 228272 220254 228324 220260
rect 228468 217410 228496 225422
rect 229388 217410 229416 228210
rect 229664 220250 229692 231676
rect 230032 223650 230060 231676
rect 230112 225752 230164 225758
rect 230112 225694 230164 225700
rect 230020 223644 230072 223650
rect 230020 223586 230072 223592
rect 230124 221270 230152 225694
rect 230296 225684 230348 225690
rect 230296 225626 230348 225632
rect 230308 221406 230336 225626
rect 230400 223242 230428 231676
rect 230768 226166 230796 231676
rect 231136 228818 231164 231676
rect 231124 228812 231176 228818
rect 231124 228754 231176 228760
rect 231504 228682 231532 231676
rect 231492 228676 231544 228682
rect 231492 228618 231544 228624
rect 231872 228546 231900 231676
rect 231860 228540 231912 228546
rect 231860 228482 231912 228488
rect 231676 228200 231728 228206
rect 231676 228142 231728 228148
rect 230756 226160 230808 226166
rect 230756 226102 230808 226108
rect 230388 223236 230440 223242
rect 230388 223178 230440 223184
rect 231032 223100 231084 223106
rect 231032 223042 231084 223048
rect 230296 221400 230348 221406
rect 230296 221342 230348 221348
rect 230112 221264 230164 221270
rect 230112 221206 230164 221212
rect 230204 221264 230256 221270
rect 230204 221206 230256 221212
rect 229652 220244 229704 220250
rect 229652 220186 229704 220192
rect 230216 217410 230244 221206
rect 231044 217410 231072 223042
rect 231688 217410 231716 228142
rect 232240 226098 232268 231676
rect 232228 226092 232280 226098
rect 232228 226034 232280 226040
rect 232516 223854 232544 231676
rect 232504 223848 232556 223854
rect 232504 223790 232556 223796
rect 232884 223378 232912 231676
rect 232872 223372 232924 223378
rect 232872 223314 232924 223320
rect 233252 223310 233280 231676
rect 233620 226302 233648 231676
rect 233988 229022 234016 231676
rect 233976 229016 234028 229022
rect 233976 228958 234028 228964
rect 234356 228886 234384 231676
rect 234344 228880 234396 228886
rect 234344 228822 234396 228828
rect 234724 228750 234752 231676
rect 234712 228744 234764 228750
rect 234712 228686 234764 228692
rect 234068 226840 234120 226846
rect 233896 226788 234068 226794
rect 233896 226782 234120 226788
rect 233896 226778 234108 226782
rect 233884 226772 234108 226778
rect 233936 226766 234108 226772
rect 233884 226714 233936 226720
rect 233608 226296 233660 226302
rect 233608 226238 233660 226244
rect 235092 226234 235120 231676
rect 235368 229090 235396 231676
rect 235356 229084 235408 229090
rect 235356 229026 235408 229032
rect 235264 228472 235316 228478
rect 235264 228414 235316 228420
rect 235538 228440 235594 228449
rect 235080 226228 235132 226234
rect 235080 226170 235132 226176
rect 234528 225616 234580 225622
rect 234528 225558 234580 225564
rect 233240 223304 233292 223310
rect 233240 223246 233292 223252
rect 232688 222964 232740 222970
rect 232688 222906 232740 222912
rect 232596 222080 232648 222086
rect 232596 222022 232648 222028
rect 232608 221814 232636 222022
rect 232596 221808 232648 221814
rect 232596 221750 232648 221756
rect 232700 217410 232728 222906
rect 234344 221808 234396 221814
rect 234344 221750 234396 221756
rect 233516 221332 233568 221338
rect 233516 221274 233568 221280
rect 233528 217410 233556 221274
rect 234356 217410 234384 221750
rect 234540 221202 234568 225558
rect 234528 221196 234580 221202
rect 234528 221138 234580 221144
rect 235276 217410 235304 228414
rect 235538 228375 235594 228384
rect 235552 221406 235580 228375
rect 235736 223514 235764 231676
rect 235828 231662 236118 231690
rect 235724 223508 235776 223514
rect 235724 223450 235776 223456
rect 235828 222154 235856 231662
rect 236472 224806 236500 231676
rect 236460 224800 236512 224806
rect 236460 224742 236512 224748
rect 236840 224058 236868 231676
rect 237208 228954 237236 231676
rect 237196 228948 237248 228954
rect 237196 228890 237248 228896
rect 237102 228576 237158 228585
rect 237102 228511 237158 228520
rect 236828 224052 236880 224058
rect 236828 223994 236880 224000
rect 236092 223032 236144 223038
rect 236092 222974 236144 222980
rect 235816 222148 235868 222154
rect 235816 222090 235868 222096
rect 235644 221610 235948 221626
rect 235632 221604 235960 221610
rect 235684 221598 235908 221604
rect 235632 221546 235684 221552
rect 235908 221546 235960 221552
rect 235540 221400 235592 221406
rect 235540 221342 235592 221348
rect 236104 217410 236132 222974
rect 236920 221400 236972 221406
rect 236920 221342 236972 221348
rect 236932 217410 236960 221342
rect 237116 220998 237144 228511
rect 237576 227662 237604 231676
rect 237564 227656 237616 227662
rect 237564 227598 237616 227604
rect 237288 226636 237340 226642
rect 237288 226578 237340 226584
rect 237300 221134 237328 226578
rect 237944 224874 237972 231676
rect 238220 227526 238248 231676
rect 238312 231662 238602 231690
rect 238208 227520 238260 227526
rect 238208 227462 238260 227468
rect 237932 224868 237984 224874
rect 237932 224810 237984 224816
rect 238312 222086 238340 231662
rect 238576 228540 238628 228546
rect 238576 228482 238628 228488
rect 238300 222080 238352 222086
rect 238300 222022 238352 222028
rect 237748 222012 237800 222018
rect 237748 221954 237800 221960
rect 237288 221128 237340 221134
rect 237288 221070 237340 221076
rect 237104 220992 237156 220998
rect 237104 220934 237156 220940
rect 237760 217410 237788 221954
rect 238588 217410 238616 228482
rect 238956 220930 238984 231676
rect 239220 228948 239272 228954
rect 239220 228890 239272 228896
rect 239232 221270 239260 228890
rect 239324 224670 239352 231676
rect 239312 224664 239364 224670
rect 239312 224606 239364 224612
rect 239692 223718 239720 231676
rect 239956 229016 240008 229022
rect 239956 228958 240008 228964
rect 239864 228676 239916 228682
rect 239864 228618 239916 228624
rect 239680 223712 239732 223718
rect 239680 223654 239732 223660
rect 239404 221740 239456 221746
rect 239404 221682 239456 221688
rect 239220 221264 239272 221270
rect 239220 221206 239272 221212
rect 238944 220924 238996 220930
rect 238944 220866 238996 220872
rect 239416 217410 239444 221682
rect 239876 221338 239904 228618
rect 239864 221332 239916 221338
rect 239864 221274 239916 221280
rect 239968 221066 239996 228958
rect 240060 227458 240088 231676
rect 240140 228608 240192 228614
rect 240140 228550 240192 228556
rect 240048 227452 240100 227458
rect 240048 227394 240100 227400
rect 240152 222578 240180 228550
rect 240428 227594 240456 231676
rect 240692 228880 240744 228886
rect 240692 228822 240744 228828
rect 240416 227588 240468 227594
rect 240416 227530 240468 227536
rect 240060 222550 240180 222578
rect 239956 221060 240008 221066
rect 239956 221002 240008 221008
rect 240060 217410 240088 222550
rect 240704 221406 240732 228822
rect 240796 224738 240824 231676
rect 241072 227254 241100 231676
rect 241440 227390 241468 231676
rect 241428 227384 241480 227390
rect 241428 227326 241480 227332
rect 241060 227248 241112 227254
rect 241060 227190 241112 227196
rect 240784 224732 240836 224738
rect 240784 224674 240836 224680
rect 241808 221882 241836 231676
rect 241980 228744 242032 228750
rect 241980 228686 242032 228692
rect 241796 221876 241848 221882
rect 241796 221818 241848 221824
rect 240968 221672 241020 221678
rect 240968 221614 241020 221620
rect 240980 221542 241008 221614
rect 241152 221604 241204 221610
rect 241152 221546 241204 221552
rect 240968 221536 241020 221542
rect 240968 221478 241020 221484
rect 240692 221400 240744 221406
rect 240692 221342 240744 221348
rect 241164 217410 241192 221546
rect 241992 217410 242020 228686
rect 242176 224602 242204 231676
rect 242164 224596 242216 224602
rect 242164 224538 242216 224544
rect 242544 223786 242572 231676
rect 242532 223780 242584 223786
rect 242532 223722 242584 223728
rect 242808 223168 242860 223174
rect 242808 223110 242860 223116
rect 242820 217410 242848 223110
rect 242912 221950 242940 231676
rect 243280 227322 243308 231676
rect 243372 231662 243662 231690
rect 243268 227316 243320 227322
rect 243268 227258 243320 227264
rect 243372 224534 243400 231662
rect 243636 227656 243688 227662
rect 243636 227598 243688 227604
rect 243360 224528 243412 224534
rect 243360 224470 243412 224476
rect 242900 221944 242952 221950
rect 242900 221886 242952 221892
rect 243648 217410 243676 227598
rect 243924 227050 243952 231676
rect 244292 227186 244320 231676
rect 244280 227180 244332 227186
rect 244280 227122 244332 227128
rect 243912 227044 243964 227050
rect 243912 226986 243964 226992
rect 243728 222352 243780 222358
rect 243728 222294 243780 222300
rect 243740 222086 243768 222294
rect 244660 222154 244688 231676
rect 245028 224398 245056 231676
rect 245292 228812 245344 228818
rect 245292 228754 245344 228760
rect 245016 224392 245068 224398
rect 245016 224334 245068 224340
rect 244648 222148 244700 222154
rect 244648 222090 244700 222096
rect 243728 222080 243780 222086
rect 243728 222022 243780 222028
rect 244464 221876 244516 221882
rect 244464 221818 244516 221824
rect 244476 217410 244504 221818
rect 245304 217410 245332 228754
rect 245396 225554 245424 231676
rect 245384 225548 245436 225554
rect 245384 225490 245436 225496
rect 245764 223446 245792 231676
rect 246132 227118 246160 231676
rect 246120 227112 246172 227118
rect 246120 227054 246172 227060
rect 246304 226500 246356 226506
rect 246304 226442 246356 226448
rect 245752 223440 245804 223446
rect 245752 223382 245804 223388
rect 246316 222222 246344 226442
rect 246500 224466 246528 231676
rect 246592 231662 246790 231690
rect 246488 224460 246540 224466
rect 246488 224402 246540 224408
rect 246304 222216 246356 222222
rect 246304 222158 246356 222164
rect 246592 221678 246620 231662
rect 247040 229084 247092 229090
rect 247040 229026 247092 229032
rect 246946 228848 247002 228857
rect 246946 228783 247002 228792
rect 246672 223304 246724 223310
rect 246672 223246 246724 223252
rect 246684 222494 246712 223246
rect 246764 223100 246816 223106
rect 246764 223042 246816 223048
rect 246776 222902 246804 223042
rect 246764 222896 246816 222902
rect 246764 222838 246816 222844
rect 246856 222896 246908 222902
rect 246856 222838 246908 222844
rect 246868 222698 246896 222838
rect 246856 222692 246908 222698
rect 246856 222634 246908 222640
rect 246672 222488 246724 222494
rect 246672 222430 246724 222436
rect 246580 221672 246632 221678
rect 246580 221614 246632 221620
rect 246960 221406 246988 228783
rect 246948 221400 247000 221406
rect 246948 221342 247000 221348
rect 246120 221196 246172 221202
rect 246120 221138 246172 221144
rect 246132 217410 246160 221138
rect 247052 217410 247080 229026
rect 247144 226982 247172 231676
rect 247132 226976 247184 226982
rect 247132 226918 247184 226924
rect 247512 221542 247540 231676
rect 247880 224330 247908 231676
rect 248248 226846 248276 231676
rect 248630 231662 248828 231690
rect 248512 227316 248564 227322
rect 248512 227258 248564 227264
rect 248420 227044 248472 227050
rect 248420 226986 248472 226992
rect 248236 226840 248288 226846
rect 248236 226782 248288 226788
rect 247868 224324 247920 224330
rect 247868 224266 247920 224272
rect 248432 223106 248460 226986
rect 248524 223242 248552 227258
rect 248604 227180 248656 227186
rect 248604 227122 248656 227128
rect 248512 223236 248564 223242
rect 248512 223178 248564 223184
rect 248420 223100 248472 223106
rect 248420 223042 248472 223048
rect 247868 222420 247920 222426
rect 247868 222362 247920 222368
rect 247500 221536 247552 221542
rect 247500 221478 247552 221484
rect 247880 217410 247908 222362
rect 248616 221814 248644 227122
rect 248696 226840 248748 226846
rect 248696 226782 248748 226788
rect 248604 221808 248656 221814
rect 248604 221750 248656 221756
rect 248708 217410 248736 226782
rect 248800 221474 248828 231662
rect 248984 226710 249012 231676
rect 248972 226704 249024 226710
rect 248972 226646 249024 226652
rect 249352 224262 249380 231676
rect 249628 225758 249656 231676
rect 249616 225752 249668 225758
rect 249616 225694 249668 225700
rect 249996 225690 250024 231676
rect 250088 231662 250378 231690
rect 249984 225684 250036 225690
rect 249984 225626 250036 225632
rect 249340 224256 249392 224262
rect 249340 224198 249392 224204
rect 249524 222488 249576 222494
rect 249524 222430 249576 222436
rect 248788 221468 248840 221474
rect 248788 221410 248840 221416
rect 249536 217410 249564 222430
rect 250088 222358 250116 231662
rect 250352 227588 250404 227594
rect 250352 227530 250404 227536
rect 250076 222352 250128 222358
rect 250076 222294 250128 222300
rect 250364 217410 250392 227530
rect 250732 224194 250760 231676
rect 251100 226574 251128 231676
rect 251272 227384 251324 227390
rect 251272 227326 251324 227332
rect 251180 227248 251232 227254
rect 251180 227190 251232 227196
rect 251088 226568 251140 226574
rect 251088 226510 251140 226516
rect 250720 224188 250772 224194
rect 250720 224130 250772 224136
rect 251088 222148 251140 222154
rect 251088 222090 251140 222096
rect 251100 217410 251128 222090
rect 251192 221610 251220 227190
rect 251284 222018 251312 227326
rect 251468 226914 251496 231676
rect 251836 227730 251864 231676
rect 251824 227724 251876 227730
rect 251824 227666 251876 227672
rect 252008 227724 252060 227730
rect 252008 227666 252060 227672
rect 251456 226908 251508 226914
rect 251456 226850 251508 226856
rect 251272 222012 251324 222018
rect 251272 221954 251324 221960
rect 251180 221604 251232 221610
rect 251180 221546 251232 221552
rect 252020 217410 252048 227666
rect 252204 224126 252232 231676
rect 252192 224120 252244 224126
rect 252192 224062 252244 224068
rect 252480 223922 252508 231676
rect 252468 223916 252520 223922
rect 252468 223858 252520 223864
rect 252848 220862 252876 231676
rect 253216 222290 253244 231676
rect 253584 225282 253612 231676
rect 253664 227520 253716 227526
rect 253664 227462 253716 227468
rect 253572 225276 253624 225282
rect 253572 225218 253624 225224
rect 253204 222284 253256 222290
rect 253204 222226 253256 222232
rect 252928 221128 252980 221134
rect 252928 221070 252980 221076
rect 252836 220856 252888 220862
rect 252836 220798 252888 220804
rect 252940 217410 252968 221070
rect 253676 217410 253704 227462
rect 253952 226522 253980 231676
rect 254044 231662 254334 231690
rect 254412 231662 254702 231690
rect 254044 227798 254072 231662
rect 254412 228154 254440 231662
rect 254320 228126 254440 228154
rect 254320 228002 254348 228126
rect 254308 227996 254360 228002
rect 254308 227938 254360 227944
rect 254400 227996 254452 228002
rect 254400 227938 254452 227944
rect 254032 227792 254084 227798
rect 254032 227734 254084 227740
rect 254216 227792 254268 227798
rect 254216 227734 254268 227740
rect 254124 227112 254176 227118
rect 254124 227054 254176 227060
rect 253860 226494 253980 226522
rect 254032 226568 254084 226574
rect 254032 226510 254084 226516
rect 253860 225622 253888 226494
rect 253940 226364 253992 226370
rect 253940 226306 253992 226312
rect 253848 225616 253900 225622
rect 253848 225558 253900 225564
rect 253952 222970 253980 226306
rect 254044 223038 254072 226510
rect 254032 223032 254084 223038
rect 254032 222974 254084 222980
rect 253940 222964 253992 222970
rect 253940 222906 253992 222912
rect 254136 221882 254164 227054
rect 254228 222154 254256 227734
rect 254308 226976 254360 226982
rect 254308 226918 254360 226924
rect 254216 222148 254268 222154
rect 254216 222090 254268 222096
rect 254124 221876 254176 221882
rect 254124 221818 254176 221824
rect 254320 221746 254348 226918
rect 254412 222426 254440 227938
rect 255056 224942 255084 231676
rect 255332 227934 255360 231676
rect 255320 227928 255372 227934
rect 255320 227870 255372 227876
rect 255044 224936 255096 224942
rect 255044 224878 255096 224884
rect 254400 222420 254452 222426
rect 254400 222362 254452 222368
rect 254584 222420 254636 222426
rect 254584 222362 254636 222368
rect 254308 221740 254360 221746
rect 254308 221682 254360 221688
rect 254596 217410 254624 222362
rect 255700 222086 255728 231676
rect 256068 223310 256096 231676
rect 256436 223990 256464 231676
rect 256698 228984 256754 228993
rect 256698 228919 256754 228928
rect 256424 223984 256476 223990
rect 256424 223926 256476 223932
rect 256056 223304 256108 223310
rect 256056 223246 256108 223252
rect 256712 222902 256740 228919
rect 256804 226642 256832 231676
rect 257172 227866 257200 231676
rect 257252 227928 257304 227934
rect 257252 227870 257304 227876
rect 257160 227860 257212 227866
rect 257160 227802 257212 227808
rect 256792 226636 256844 226642
rect 256792 226578 256844 226584
rect 256700 222896 256752 222902
rect 256700 222838 256752 222844
rect 257068 222896 257120 222902
rect 257068 222838 257120 222844
rect 255688 222080 255740 222086
rect 255688 222022 255740 222028
rect 255412 221808 255464 221814
rect 255412 221750 255464 221756
rect 255424 217410 255452 221750
rect 256240 221400 256292 221406
rect 256240 221342 256292 221348
rect 256252 217410 256280 221342
rect 257080 217410 257108 222838
rect 257264 221134 257292 227870
rect 257344 227452 257396 227458
rect 257344 227394 257396 227400
rect 257356 222834 257384 227394
rect 257344 222828 257396 222834
rect 257344 222770 257396 222776
rect 257540 222630 257568 231676
rect 257804 226908 257856 226914
rect 257804 226850 257856 226856
rect 257528 222624 257580 222630
rect 257528 222566 257580 222572
rect 257816 221202 257844 226850
rect 257908 225010 257936 231676
rect 258184 228070 258212 231676
rect 258172 228064 258224 228070
rect 258172 228006 258224 228012
rect 258448 226772 258500 226778
rect 258448 226714 258500 226720
rect 257896 225004 257948 225010
rect 257896 224946 257948 224952
rect 258460 223174 258488 226714
rect 258552 226506 258580 231676
rect 258540 226500 258592 226506
rect 258540 226442 258592 226448
rect 258448 223168 258500 223174
rect 258448 223110 258500 223116
rect 258920 222766 258948 231676
rect 259288 225078 259316 231676
rect 259656 228585 259684 231676
rect 259642 228576 259698 228585
rect 259642 228511 259698 228520
rect 259368 228064 259420 228070
rect 259368 228006 259420 228012
rect 259276 225072 259328 225078
rect 259276 225014 259328 225020
rect 258908 222760 258960 222766
rect 258908 222702 258960 222708
rect 259380 222494 259408 228006
rect 260024 227769 260052 231676
rect 260010 227760 260066 227769
rect 260010 227695 260066 227704
rect 260392 227633 260420 231676
rect 260378 227624 260434 227633
rect 260378 227559 260434 227568
rect 260760 225146 260788 231676
rect 261036 228138 261064 231676
rect 261404 228857 261432 231676
rect 261772 228993 261800 231676
rect 261758 228984 261814 228993
rect 261758 228919 261814 228928
rect 261390 228848 261446 228857
rect 261390 228783 261446 228792
rect 261024 228132 261076 228138
rect 261024 228074 261076 228080
rect 261484 227860 261536 227866
rect 261484 227802 261536 227808
rect 260748 225140 260800 225146
rect 260748 225082 260800 225088
rect 261300 222828 261352 222834
rect 261300 222770 261352 222776
rect 260472 222692 260524 222698
rect 260472 222634 260524 222640
rect 259368 222488 259420 222494
rect 259368 222430 259420 222436
rect 259368 222352 259420 222358
rect 259368 222294 259420 222300
rect 257896 222216 257948 222222
rect 257896 222158 257948 222164
rect 257804 221196 257856 221202
rect 257804 221138 257856 221144
rect 257252 221128 257304 221134
rect 257252 221070 257304 221076
rect 257908 217410 257936 222158
rect 258816 221740 258868 221746
rect 258816 221682 258868 221688
rect 258828 217410 258856 221682
rect 259380 217410 259408 222294
rect 260484 217410 260512 222634
rect 261312 217410 261340 222770
rect 261496 221406 261524 227802
rect 262140 225418 262168 231676
rect 262508 228449 262536 231676
rect 262494 228440 262550 228449
rect 262494 228375 262550 228384
rect 262876 227905 262904 231676
rect 263244 228041 263272 231676
rect 263230 228032 263286 228041
rect 263230 227967 263286 227976
rect 262862 227896 262918 227905
rect 262862 227831 262918 227840
rect 262128 225412 262180 225418
rect 262128 225354 262180 225360
rect 263612 225350 263640 231676
rect 263888 228342 263916 231676
rect 263876 228336 263928 228342
rect 263876 228278 263928 228284
rect 264256 228177 264284 231676
rect 264242 228168 264298 228177
rect 264242 228103 264298 228112
rect 264624 227458 264652 231676
rect 264612 227452 264664 227458
rect 264612 227394 264664 227400
rect 264704 227452 264756 227458
rect 264704 227394 264756 227400
rect 264716 226846 264744 227394
rect 264704 226840 264756 226846
rect 264704 226782 264756 226788
rect 263600 225344 263652 225350
rect 263600 225286 263652 225292
rect 264992 225214 265020 231676
rect 265360 229022 265388 231676
rect 265348 229016 265400 229022
rect 265348 228958 265400 228964
rect 265728 227050 265756 231676
rect 266096 228313 266124 231676
rect 266082 228304 266138 228313
rect 266082 228239 266138 228248
rect 265716 227044 265768 227050
rect 265716 226986 265768 226992
rect 266464 225486 266492 231676
rect 266740 228954 266768 231676
rect 266728 228948 266780 228954
rect 266728 228890 266780 228896
rect 267108 228410 267136 231676
rect 267096 228404 267148 228410
rect 267096 228346 267148 228352
rect 267476 228274 267504 231676
rect 267464 228268 267516 228274
rect 267464 228210 267516 228216
rect 267844 228206 267872 231676
rect 268212 228682 268240 231676
rect 268200 228676 268252 228682
rect 268200 228618 268252 228624
rect 267832 228200 267884 228206
rect 267832 228142 267884 228148
rect 268580 227322 268608 231676
rect 268568 227316 268620 227322
rect 268568 227258 268620 227264
rect 268948 226370 268976 231676
rect 269316 228478 269344 231676
rect 269592 228886 269620 231676
rect 269580 228880 269632 228886
rect 269580 228822 269632 228828
rect 269304 228472 269356 228478
rect 269304 228414 269356 228420
rect 269960 227186 269988 231676
rect 269948 227180 270000 227186
rect 269948 227122 270000 227128
rect 270328 226574 270356 231676
rect 270696 228546 270724 231676
rect 271064 228614 271092 231676
rect 271052 228608 271104 228614
rect 271052 228550 271104 228556
rect 270684 228540 270736 228546
rect 270684 228482 270736 228488
rect 271432 227390 271460 231676
rect 271420 227384 271472 227390
rect 271420 227326 271472 227332
rect 271800 226982 271828 231676
rect 272168 228750 272196 231676
rect 272156 228744 272208 228750
rect 272156 228686 272208 228692
rect 272444 227662 272472 231676
rect 272432 227656 272484 227662
rect 272432 227598 272484 227604
rect 272812 227254 272840 231676
rect 272800 227248 272852 227254
rect 272800 227190 272852 227196
rect 271788 226976 271840 226982
rect 271788 226918 271840 226924
rect 273180 226778 273208 231676
rect 273548 228818 273576 231676
rect 273916 229090 273944 231676
rect 273904 229084 273956 229090
rect 273904 229026 273956 229032
rect 273536 228812 273588 228818
rect 273536 228754 273588 228760
rect 274284 227118 274312 231676
rect 274272 227112 274324 227118
rect 274272 227054 274324 227060
rect 274652 226914 274680 231676
rect 275020 227458 275048 231676
rect 275296 227594 275324 231676
rect 275664 228002 275692 231676
rect 276032 228070 276060 231676
rect 276020 228064 276072 228070
rect 276020 228006 276072 228012
rect 275652 227996 275704 228002
rect 275652 227938 275704 227944
rect 276400 227730 276428 231676
rect 276388 227724 276440 227730
rect 276388 227666 276440 227672
rect 275284 227588 275336 227594
rect 275284 227530 275336 227536
rect 276768 227526 276796 231676
rect 277136 227798 277164 231676
rect 277504 227934 277532 231676
rect 277492 227928 277544 227934
rect 277492 227870 277544 227876
rect 277124 227792 277176 227798
rect 277124 227734 277176 227740
rect 276756 227520 276808 227526
rect 276756 227462 276808 227468
rect 275008 227452 275060 227458
rect 275008 227394 275060 227400
rect 274640 226908 274692 226914
rect 274640 226850 274692 226856
rect 273168 226772 273220 226778
rect 273168 226714 273220 226720
rect 270316 226568 270368 226574
rect 270316 226510 270368 226516
rect 268936 226364 268988 226370
rect 268936 226306 268988 226312
rect 266452 225480 266504 225486
rect 266452 225422 266504 225428
rect 264980 225208 265032 225214
rect 264980 225150 265032 225156
rect 269672 223304 269724 223310
rect 269672 223246 269724 223252
rect 263784 223032 263836 223038
rect 263784 222974 263836 222980
rect 262956 222760 263008 222766
rect 262956 222702 263008 222708
rect 262128 222624 262180 222630
rect 262128 222566 262180 222572
rect 261484 221400 261536 221406
rect 261484 221342 261536 221348
rect 262140 217410 262168 222566
rect 262968 217410 262996 222702
rect 263796 217410 263824 222974
rect 266360 222964 266412 222970
rect 266360 222906 266412 222912
rect 264612 222556 264664 222562
rect 264612 222498 264664 222504
rect 264624 217410 264652 222498
rect 265532 221128 265584 221134
rect 265532 221070 265584 221076
rect 265544 217410 265572 221070
rect 266372 217410 266400 222906
rect 268844 221604 268896 221610
rect 268844 221546 268896 221552
rect 267188 221400 267240 221406
rect 267188 221342 267240 221348
rect 267200 217410 267228 221342
rect 268016 220992 268068 220998
rect 268016 220934 268068 220940
rect 268028 217410 268056 220934
rect 268856 217410 268884 221546
rect 269684 217410 269712 223246
rect 271420 223100 271472 223106
rect 271420 223042 271472 223048
rect 270408 221536 270460 221542
rect 270408 221478 270460 221484
rect 270420 217410 270448 221478
rect 271432 217410 271460 223042
rect 272248 222488 272300 222494
rect 272248 222430 272300 222436
rect 272260 217410 272288 222430
rect 273076 222148 273128 222154
rect 273076 222090 273128 222096
rect 273088 217410 273116 222090
rect 274732 221876 274784 221882
rect 274732 221818 274784 221824
rect 273904 221672 273956 221678
rect 273904 221614 273956 221620
rect 273916 217410 273944 221614
rect 274744 217410 274772 221818
rect 277872 221814 277900 231676
rect 278148 222902 278176 231676
rect 278136 222896 278188 222902
rect 278136 222838 278188 222844
rect 278516 222426 278544 231676
rect 278884 227866 278912 231676
rect 278872 227860 278924 227866
rect 278872 227802 278924 227808
rect 278688 223576 278740 223582
rect 278688 223518 278740 223524
rect 278504 222420 278556 222426
rect 278504 222362 278556 222368
rect 277860 221808 277912 221814
rect 277860 221750 277912 221756
rect 275560 221468 275612 221474
rect 275560 221410 275612 221416
rect 275572 217410 275600 221410
rect 277308 221264 277360 221270
rect 277308 221206 277360 221212
rect 276480 220924 276532 220930
rect 276480 220866 276532 220872
rect 276492 217410 276520 220866
rect 277320 217410 277348 221206
rect 278136 221060 278188 221066
rect 278136 221002 278188 221008
rect 278148 217410 278176 221002
rect 278700 217410 278728 223518
rect 279252 221746 279280 231676
rect 279620 222698 279648 231676
rect 279608 222692 279660 222698
rect 279608 222634 279660 222640
rect 279988 222222 280016 231676
rect 280356 222358 280384 231676
rect 280724 222630 280752 231676
rect 281000 223038 281028 231676
rect 280988 223032 281040 223038
rect 280988 222974 281040 222980
rect 281368 222834 281396 231676
rect 281356 222828 281408 222834
rect 281356 222770 281408 222776
rect 281736 222766 281764 231676
rect 281724 222760 281776 222766
rect 281724 222702 281776 222708
rect 280712 222624 280764 222630
rect 280712 222566 280764 222572
rect 280344 222352 280396 222358
rect 280344 222294 280396 222300
rect 279976 222216 280028 222222
rect 279976 222158 280028 222164
rect 281448 222216 281500 222222
rect 281448 222158 281500 222164
rect 279240 221740 279292 221746
rect 279240 221682 279292 221688
rect 280620 221332 280672 221338
rect 280620 221274 280672 221280
rect 279792 221196 279844 221202
rect 279792 221138 279844 221144
rect 279804 217410 279832 221138
rect 280632 217410 280660 221274
rect 281460 217410 281488 222158
rect 282104 221134 282132 231676
rect 282472 221406 282500 231676
rect 282840 222562 282868 231676
rect 283208 222970 283236 231676
rect 283196 222964 283248 222970
rect 283196 222906 283248 222912
rect 282828 222556 282880 222562
rect 282828 222498 282880 222504
rect 283196 222556 283248 222562
rect 283196 222498 283248 222504
rect 282460 221400 282512 221406
rect 282460 221342 282512 221348
rect 282092 221128 282144 221134
rect 282092 221070 282144 221076
rect 282368 221128 282420 221134
rect 282368 221070 282420 221076
rect 282380 217410 282408 221070
rect 283208 217410 283236 222498
rect 283576 221610 283604 231676
rect 283564 221604 283616 221610
rect 283564 221546 283616 221552
rect 283852 221542 283880 231676
rect 283932 221740 283984 221746
rect 283932 221682 283984 221688
rect 283840 221536 283892 221542
rect 283840 221478 283892 221484
rect 283944 217410 283972 221682
rect 284220 220998 284248 231676
rect 284588 223310 284616 231676
rect 284576 223304 284628 223310
rect 284576 223246 284628 223252
rect 284956 222630 284984 231676
rect 284944 222624 284996 222630
rect 284944 222566 284996 222572
rect 285324 221814 285352 231676
rect 285692 223106 285720 231676
rect 285680 223100 285732 223106
rect 285680 223042 285732 223048
rect 286060 222154 286088 231676
rect 286048 222148 286100 222154
rect 286048 222090 286100 222096
rect 285312 221808 285364 221814
rect 285312 221750 285364 221756
rect 284852 221536 284904 221542
rect 284852 221478 284904 221484
rect 284208 220992 284260 220998
rect 284208 220934 284260 220940
rect 284864 217410 284892 221478
rect 286428 221474 286456 231676
rect 286416 221468 286468 221474
rect 286416 221410 286468 221416
rect 286508 221468 286560 221474
rect 286508 221410 286560 221416
rect 285680 220992 285732 220998
rect 285680 220934 285732 220940
rect 285692 217410 285720 220934
rect 286520 217410 286548 221410
rect 286704 221270 286732 231676
rect 287072 221882 287100 231676
rect 287060 221876 287112 221882
rect 287060 221818 287112 221824
rect 287152 221876 287204 221882
rect 287152 221818 287204 221824
rect 287060 221672 287112 221678
rect 287060 221614 287112 221620
rect 286692 221264 286744 221270
rect 286692 221206 286744 221212
rect 287072 221066 287100 221614
rect 287164 221134 287192 221818
rect 287152 221128 287204 221134
rect 287152 221070 287204 221076
rect 287060 221060 287112 221066
rect 287060 221002 287112 221008
rect 287336 221060 287388 221066
rect 287336 221002 287388 221008
rect 287348 217410 287376 221002
rect 287440 220930 287468 231676
rect 287808 223582 287836 231676
rect 287796 223576 287848 223582
rect 287796 223518 287848 223524
rect 288176 221338 288204 231676
rect 288544 221678 288572 231676
rect 288532 221672 288584 221678
rect 288532 221614 288584 221620
rect 288164 221332 288216 221338
rect 288164 221274 288216 221280
rect 288912 221202 288940 231676
rect 289280 221882 289308 231676
rect 289268 221876 289320 221882
rect 289268 221818 289320 221824
rect 289556 221746 289584 231676
rect 289924 222222 289952 231676
rect 290292 222562 290320 231676
rect 290280 222556 290332 222562
rect 290280 222498 290332 222504
rect 289912 222216 289964 222222
rect 289912 222158 289964 222164
rect 289544 221740 289596 221746
rect 289544 221682 289596 221688
rect 289084 221400 289136 221406
rect 289084 221342 289136 221348
rect 288900 221196 288952 221202
rect 288900 221138 288952 221144
rect 288256 221128 288308 221134
rect 288256 221070 288308 221076
rect 287428 220924 287480 220930
rect 287428 220866 287480 220872
rect 288268 217410 288296 221070
rect 289096 217410 289124 221342
rect 289728 221332 289780 221338
rect 289728 221274 289780 221280
rect 289740 217410 289768 221274
rect 290660 220998 290688 231676
rect 290740 229016 290792 229022
rect 290740 228958 290792 228964
rect 290648 220992 290700 220998
rect 290648 220934 290700 220940
rect 290752 217410 290780 228958
rect 291028 221066 291056 231676
rect 291396 221542 291424 231676
rect 291384 221536 291436 221542
rect 291384 221478 291436 221484
rect 291764 221474 291792 231676
rect 291752 221468 291804 221474
rect 291752 221410 291804 221416
rect 292132 221406 292160 231676
rect 292408 229022 292436 231676
rect 292396 229016 292448 229022
rect 292396 228958 292448 228964
rect 292120 221400 292172 221406
rect 292120 221342 292172 221348
rect 292396 221400 292448 221406
rect 292396 221342 292448 221348
rect 291016 221060 291068 221066
rect 291016 221002 291068 221008
rect 291568 220992 291620 220998
rect 291568 220934 291620 220940
rect 291580 217410 291608 220934
rect 292408 217410 292436 221342
rect 292776 221134 292804 231676
rect 293144 221338 293172 231676
rect 293224 229016 293276 229022
rect 293224 228958 293276 228964
rect 293132 221332 293184 221338
rect 293132 221274 293184 221280
rect 292764 221128 292816 221134
rect 292764 221070 292816 221076
rect 293236 217410 293264 228958
rect 293512 221406 293540 231676
rect 293500 221400 293552 221406
rect 293500 221342 293552 221348
rect 293880 217410 293908 231676
rect 294248 220998 294276 231676
rect 294616 229022 294644 231676
rect 294998 231662 295196 231690
rect 294604 229016 294656 229022
rect 294604 228958 294656 228964
rect 295168 226334 295196 231662
rect 295260 227322 295288 231676
rect 295248 227316 295300 227322
rect 295248 227258 295300 227264
rect 295168 226306 295380 226334
rect 294972 221332 295024 221338
rect 294972 221274 295024 221280
rect 294236 220992 294288 220998
rect 294236 220934 294288 220940
rect 294984 217410 295012 221274
rect 170968 217382 171028 217410
rect 171856 217382 172192 217410
rect 172684 217382 173020 217410
rect 173512 217382 173664 217410
rect 174340 217382 174676 217410
rect 175168 217382 175504 217410
rect 176088 217382 176424 217410
rect 176916 217382 177252 217410
rect 177744 217382 178080 217410
rect 178572 217382 178908 217410
rect 179400 217382 179736 217410
rect 180228 217382 180564 217410
rect 181056 217382 181392 217410
rect 181976 217382 182128 217410
rect 182804 217382 183140 217410
rect 183632 217382 183968 217410
rect 184460 217382 184796 217410
rect 185288 217382 185624 217410
rect 186116 217382 186452 217410
rect 186944 217382 187280 217410
rect 187864 217382 188200 217410
rect 188692 217382 189028 217410
rect 189520 217382 189856 217410
rect 190348 217382 190408 217410
rect 191176 217382 191512 217410
rect 192004 217382 192340 217410
rect 192832 217382 192984 217410
rect 193752 217382 194088 217410
rect 194580 217382 195008 217410
rect 195408 217382 195744 217410
rect 196236 217382 196572 217410
rect 197064 217382 197492 217410
rect 197892 217382 198228 217410
rect 198720 217382 199056 217410
rect 199640 217382 199976 217410
rect 200468 217382 200804 217410
rect 201296 217382 201448 217410
rect 202124 217382 202460 217410
rect 202952 217382 203288 217410
rect 203780 217382 204116 217410
rect 204608 217382 204944 217410
rect 205528 217382 205864 217410
rect 206356 217382 206692 217410
rect 207184 217382 207520 217410
rect 208012 217382 208348 217410
rect 208840 217382 209176 217410
rect 209668 217382 209728 217410
rect 210496 217382 210832 217410
rect 211416 217382 211752 217410
rect 212244 217382 212396 217410
rect 213072 217382 213408 217410
rect 213900 217382 214236 217410
rect 214728 217382 215064 217410
rect 215556 217382 215892 217410
rect 216384 217382 216720 217410
rect 217304 217382 217640 217410
rect 218132 217382 218468 217410
rect 218960 217382 219296 217410
rect 219788 217382 220124 217410
rect 220616 217382 220768 217410
rect 221444 217382 221780 217410
rect 222272 217382 222608 217410
rect 223192 217382 223528 217410
rect 224020 217382 224356 217410
rect 224848 217382 225184 217410
rect 225676 217382 226012 217410
rect 226504 217382 226840 217410
rect 227332 217382 227668 217410
rect 228160 217382 228496 217410
rect 229080 217382 229416 217410
rect 229908 217382 230244 217410
rect 230736 217382 231072 217410
rect 231564 217382 231716 217410
rect 232392 217382 232728 217410
rect 233220 217382 233556 217410
rect 234048 217382 234384 217410
rect 234968 217382 235304 217410
rect 235796 217382 236132 217410
rect 236624 217382 236960 217410
rect 237452 217382 237788 217410
rect 238280 217382 238616 217410
rect 239108 217382 239444 217410
rect 239936 217382 240088 217410
rect 240856 217382 241192 217410
rect 241684 217382 242020 217410
rect 242512 217382 242848 217410
rect 243340 217382 243676 217410
rect 244168 217382 244504 217410
rect 244996 217382 245332 217410
rect 245824 217382 246160 217410
rect 246744 217382 247080 217410
rect 247572 217382 247908 217410
rect 248400 217382 248736 217410
rect 249228 217382 249564 217410
rect 250056 217382 250392 217410
rect 250884 217382 251128 217410
rect 251712 217382 252048 217410
rect 252632 217382 252968 217410
rect 253460 217382 253704 217410
rect 254288 217382 254624 217410
rect 255116 217382 255452 217410
rect 255944 217382 256280 217410
rect 256772 217382 257108 217410
rect 257600 217382 257936 217410
rect 258520 217382 258856 217410
rect 259348 217382 259408 217410
rect 260176 217382 260512 217410
rect 261004 217382 261340 217410
rect 261832 217382 262168 217410
rect 262660 217382 262996 217410
rect 263488 217382 263824 217410
rect 264408 217382 264652 217410
rect 265236 217382 265572 217410
rect 266064 217382 266400 217410
rect 266892 217382 267228 217410
rect 267720 217382 268056 217410
rect 268548 217382 268884 217410
rect 269376 217382 269712 217410
rect 270296 217382 270448 217410
rect 271124 217382 271460 217410
rect 271952 217382 272288 217410
rect 272780 217382 273116 217410
rect 273608 217382 273944 217410
rect 274436 217382 274772 217410
rect 275264 217382 275600 217410
rect 276184 217382 276520 217410
rect 277012 217382 277348 217410
rect 277840 217382 278176 217410
rect 278668 217382 278728 217410
rect 279496 217382 279832 217410
rect 280324 217382 280660 217410
rect 281152 217382 281488 217410
rect 282072 217382 282408 217410
rect 282900 217382 283236 217410
rect 283728 217382 283972 217410
rect 284556 217382 284892 217410
rect 285384 217382 285720 217410
rect 286212 217382 286548 217410
rect 287040 217382 287376 217410
rect 287960 217382 288296 217410
rect 288788 217382 289124 217410
rect 289616 217382 289768 217410
rect 290444 217382 290780 217410
rect 291272 217382 291608 217410
rect 292100 217382 292436 217410
rect 292928 217382 293264 217410
rect 293848 217382 293908 217410
rect 294676 217382 295012 217410
rect 295352 217410 295380 226306
rect 295628 221338 295656 231676
rect 295616 221332 295668 221338
rect 295616 221274 295668 221280
rect 295996 217410 296024 231676
rect 296364 229090 296392 231676
rect 296352 229084 296404 229090
rect 296352 229026 296404 229032
rect 296732 226642 296760 231676
rect 297114 231662 297404 231690
rect 296812 227316 296864 227322
rect 296812 227258 296864 227264
rect 296720 226636 296772 226642
rect 296720 226578 296772 226584
rect 296824 217410 296852 227258
rect 297376 226334 297404 231662
rect 297468 229022 297496 231676
rect 297456 229016 297508 229022
rect 297456 228958 297508 228964
rect 297836 228954 297864 231676
rect 297824 228948 297876 228954
rect 297824 228890 297876 228896
rect 298112 226710 298140 231676
rect 298494 231662 298784 231690
rect 298468 229084 298520 229090
rect 298468 229026 298520 229032
rect 298100 226704 298152 226710
rect 298100 226646 298152 226652
rect 297376 226306 297588 226334
rect 297560 217410 297588 226306
rect 298480 217410 298508 229026
rect 298756 227322 298784 231662
rect 298848 228750 298876 231676
rect 298836 228744 298888 228750
rect 298836 228686 298888 228692
rect 298744 227316 298796 227322
rect 298744 227258 298796 227264
rect 299216 226778 299244 231676
rect 299388 229016 299440 229022
rect 299388 228958 299440 228964
rect 299204 226772 299256 226778
rect 299204 226714 299256 226720
rect 299400 217410 299428 228958
rect 299584 226846 299612 231676
rect 299572 226840 299624 226846
rect 299572 226782 299624 226788
rect 299952 226370 299980 231676
rect 300320 226642 300348 231676
rect 300688 226914 300716 231676
rect 300964 228206 300992 231676
rect 300952 228200 301004 228206
rect 300952 228142 301004 228148
rect 301044 227316 301096 227322
rect 301044 227258 301096 227264
rect 300676 226908 300728 226914
rect 300676 226850 300728 226856
rect 300216 226636 300268 226642
rect 300216 226578 300268 226584
rect 300308 226636 300360 226642
rect 300308 226578 300360 226584
rect 299940 226364 299992 226370
rect 299940 226306 299992 226312
rect 300228 217410 300256 226578
rect 301056 217410 301084 227258
rect 301332 226574 301360 231676
rect 301700 227934 301728 231676
rect 301872 228948 301924 228954
rect 301872 228890 301924 228896
rect 301688 227928 301740 227934
rect 301688 227870 301740 227876
rect 301320 226568 301372 226574
rect 301320 226510 301372 226516
rect 301884 217410 301912 228890
rect 302068 227254 302096 231676
rect 302436 227322 302464 231676
rect 302700 228744 302752 228750
rect 302700 228686 302752 228692
rect 302424 227316 302476 227322
rect 302424 227258 302476 227264
rect 302056 227248 302108 227254
rect 302056 227190 302108 227196
rect 302712 217410 302740 228686
rect 302804 228002 302832 231676
rect 302792 227996 302844 228002
rect 302792 227938 302844 227944
rect 303172 227526 303200 231676
rect 303540 228546 303568 231676
rect 303528 228540 303580 228546
rect 303528 228482 303580 228488
rect 303816 227866 303844 231676
rect 304184 229022 304212 231676
rect 304552 229090 304580 231676
rect 304540 229084 304592 229090
rect 304540 229026 304592 229032
rect 304172 229016 304224 229022
rect 304172 228958 304224 228964
rect 303804 227860 303856 227866
rect 303804 227802 303856 227808
rect 304920 227798 304948 231676
rect 304908 227792 304960 227798
rect 304908 227734 304960 227740
rect 305288 227662 305316 231676
rect 305656 228954 305684 231676
rect 305644 228948 305696 228954
rect 305644 228890 305696 228896
rect 306024 228478 306052 231676
rect 306012 228472 306064 228478
rect 306012 228414 306064 228420
rect 305276 227656 305328 227662
rect 305276 227598 305328 227604
rect 303160 227520 303212 227526
rect 303160 227462 303212 227468
rect 306392 226778 306420 231676
rect 306668 228682 306696 231676
rect 306656 228676 306708 228682
rect 306656 228618 306708 228624
rect 307036 227594 307064 231676
rect 307404 228750 307432 231676
rect 307392 228744 307444 228750
rect 307392 228686 307444 228692
rect 307772 228342 307800 231676
rect 308140 228614 308168 231676
rect 308508 228886 308536 231676
rect 308496 228880 308548 228886
rect 308496 228822 308548 228828
rect 308128 228608 308180 228614
rect 308128 228550 308180 228556
rect 307760 228336 307812 228342
rect 307760 228278 307812 228284
rect 308876 228138 308904 231676
rect 309244 228274 309272 231676
rect 309520 228410 309548 231676
rect 309508 228404 309560 228410
rect 309508 228346 309560 228352
rect 309232 228268 309284 228274
rect 309232 228210 309284 228216
rect 308864 228132 308916 228138
rect 308864 228074 308916 228080
rect 309416 227928 309468 227934
rect 309416 227870 309468 227876
rect 307024 227588 307076 227594
rect 307024 227530 307076 227536
rect 308588 226908 308640 226914
rect 308588 226850 308640 226856
rect 306932 226840 306984 226846
rect 306932 226782 306984 226788
rect 305276 226772 305328 226778
rect 305276 226714 305328 226720
rect 306380 226772 306432 226778
rect 306380 226714 306432 226720
rect 303620 226704 303672 226710
rect 303620 226646 303672 226652
rect 303632 217410 303660 226646
rect 304356 226364 304408 226370
rect 304356 226306 304408 226312
rect 304368 217410 304396 226306
rect 305288 217410 305316 226714
rect 306380 226636 306432 226642
rect 306380 226578 306432 226584
rect 306392 217410 306420 226578
rect 306944 217410 306972 226782
rect 307760 226568 307812 226574
rect 307760 226510 307812 226516
rect 307772 217410 307800 226510
rect 308600 217410 308628 226850
rect 309428 217410 309456 227870
rect 309888 226370 309916 231676
rect 310270 231662 310560 231690
rect 310532 228206 310560 231662
rect 310624 228818 310652 231676
rect 310612 228812 310664 228818
rect 310612 228754 310664 228760
rect 310244 228200 310296 228206
rect 310244 228142 310296 228148
rect 310520 228200 310572 228206
rect 310520 228142 310572 228148
rect 309876 226364 309928 226370
rect 309876 226306 309928 226312
rect 310256 217410 310284 228142
rect 310992 222358 311020 231676
rect 311360 228002 311388 231676
rect 311728 228070 311756 231676
rect 311716 228064 311768 228070
rect 311716 228006 311768 228012
rect 311164 227996 311216 228002
rect 311164 227938 311216 227944
rect 311348 227996 311400 228002
rect 311348 227938 311400 227944
rect 310980 222352 311032 222358
rect 310980 222294 311032 222300
rect 311176 217410 311204 227938
rect 312096 227730 312124 231676
rect 312084 227724 312136 227730
rect 312084 227666 312136 227672
rect 311992 227248 312044 227254
rect 311992 227190 312044 227196
rect 312004 217410 312032 227190
rect 312372 221202 312400 231676
rect 312740 227934 312768 231676
rect 312728 227928 312780 227934
rect 312728 227870 312780 227876
rect 312820 227520 312872 227526
rect 312820 227462 312872 227468
rect 312360 221196 312412 221202
rect 312360 221138 312412 221144
rect 312832 217410 312860 227462
rect 313108 222222 313136 231676
rect 313476 225078 313504 231676
rect 313648 227316 313700 227322
rect 313648 227258 313700 227264
rect 313464 225072 313516 225078
rect 313464 225014 313516 225020
rect 313096 222216 313148 222222
rect 313096 222158 313148 222164
rect 313660 217410 313688 227258
rect 313844 221610 313872 231676
rect 314212 222290 314240 231676
rect 314200 222284 314252 222290
rect 314200 222226 314252 222232
rect 313832 221604 313884 221610
rect 313832 221546 313884 221552
rect 314580 221406 314608 231676
rect 314660 229016 314712 229022
rect 314660 228958 314712 228964
rect 314568 221400 314620 221406
rect 314568 221342 314620 221348
rect 314672 217410 314700 228958
rect 314948 224942 314976 231676
rect 314936 224936 314988 224942
rect 314936 224878 314988 224884
rect 315224 221474 315252 231676
rect 315304 228540 315356 228546
rect 315304 228482 315356 228488
rect 315212 221468 315264 221474
rect 315212 221410 315264 221416
rect 315316 217410 315344 228482
rect 315592 221270 315620 231676
rect 315960 221338 315988 231676
rect 316132 229084 316184 229090
rect 316132 229026 316184 229032
rect 315948 221332 316000 221338
rect 315948 221274 316000 221280
rect 315580 221264 315632 221270
rect 315580 221206 315632 221212
rect 316144 217410 316172 229026
rect 316328 225010 316356 231676
rect 316316 225004 316368 225010
rect 316316 224946 316368 224952
rect 316696 221678 316724 231676
rect 316684 221672 316736 221678
rect 316684 221614 316736 221620
rect 317064 221542 317092 231676
rect 317432 228546 317460 231676
rect 317420 228540 317472 228546
rect 317420 228482 317472 228488
rect 317420 227860 317472 227866
rect 317420 227802 317472 227808
rect 317052 221536 317104 221542
rect 317052 221478 317104 221484
rect 317432 217410 317460 227802
rect 317800 225214 317828 231676
rect 317880 228948 317932 228954
rect 317880 228890 317932 228896
rect 317788 225208 317840 225214
rect 317788 225150 317840 225156
rect 295352 217382 295504 217410
rect 295996 217382 296332 217410
rect 296824 217382 297160 217410
rect 297560 217382 297988 217410
rect 298480 217382 298816 217410
rect 299400 217382 299736 217410
rect 300228 217382 300564 217410
rect 301056 217382 301392 217410
rect 301884 217382 302220 217410
rect 302712 217382 303048 217410
rect 303632 217382 303876 217410
rect 304368 217382 304704 217410
rect 305288 217382 305624 217410
rect 306392 217382 306452 217410
rect 306944 217382 307280 217410
rect 307772 217382 308108 217410
rect 308600 217382 308936 217410
rect 309428 217382 309764 217410
rect 310256 217382 310592 217410
rect 311176 217382 311512 217410
rect 312004 217382 312340 217410
rect 312832 217382 313168 217410
rect 313660 217382 313996 217410
rect 314672 217382 314824 217410
rect 315316 217382 315652 217410
rect 316144 217382 316480 217410
rect 317400 217382 317460 217410
rect 317892 217410 317920 228890
rect 318076 221882 318104 231676
rect 318444 223582 318472 231676
rect 318812 227866 318840 231676
rect 318800 227860 318852 227866
rect 318800 227802 318852 227808
rect 318708 227792 318760 227798
rect 318708 227734 318760 227740
rect 318432 223576 318484 223582
rect 318432 223518 318484 223524
rect 318064 221876 318116 221882
rect 318064 221818 318116 221824
rect 318720 217410 318748 227734
rect 319180 225146 319208 231676
rect 319562 231662 319852 231690
rect 319536 228472 319588 228478
rect 319536 228414 319588 228420
rect 319168 225140 319220 225146
rect 319168 225082 319220 225088
rect 319548 217410 319576 228414
rect 319824 221950 319852 231662
rect 319812 221944 319864 221950
rect 319812 221886 319864 221892
rect 319916 221746 319944 231676
rect 320284 228954 320312 231676
rect 320272 228948 320324 228954
rect 320272 228890 320324 228896
rect 320652 227662 320680 231676
rect 320364 227656 320416 227662
rect 320364 227598 320416 227604
rect 320640 227656 320692 227662
rect 320640 227598 320692 227604
rect 319904 221740 319956 221746
rect 319904 221682 319956 221688
rect 320376 217410 320404 227598
rect 320928 222086 320956 231676
rect 321192 227588 321244 227594
rect 321192 227530 321244 227536
rect 320916 222080 320968 222086
rect 320916 222022 320968 222028
rect 321204 217410 321232 227530
rect 321296 221814 321324 231676
rect 321664 222154 321692 231676
rect 322032 227050 322060 231676
rect 322020 227044 322072 227050
rect 322020 226986 322072 226992
rect 322020 226772 322072 226778
rect 322020 226714 322072 226720
rect 321652 222148 321704 222154
rect 321652 222090 321704 222096
rect 321284 221808 321336 221814
rect 321284 221750 321336 221756
rect 322032 217410 322060 226714
rect 322400 223514 322428 231676
rect 322388 223508 322440 223514
rect 322388 223450 322440 223456
rect 322768 222018 322796 231676
rect 322940 228744 322992 228750
rect 322940 228686 322992 228692
rect 322756 222012 322808 222018
rect 322756 221954 322808 221960
rect 322952 217410 322980 228686
rect 323136 227390 323164 231676
rect 323124 227384 323176 227390
rect 323124 227326 323176 227332
rect 323504 226846 323532 231676
rect 323794 231662 324084 231690
rect 323768 228676 323820 228682
rect 323768 228618 323820 228624
rect 323492 226840 323544 226846
rect 323492 226782 323544 226788
rect 323780 217410 323808 228618
rect 324056 223038 324084 231662
rect 324148 223310 324176 231676
rect 324516 227526 324544 231676
rect 324596 228880 324648 228886
rect 324596 228822 324648 228828
rect 324504 227520 324556 227526
rect 324504 227462 324556 227468
rect 324136 223304 324188 223310
rect 324136 223246 324188 223252
rect 324044 223032 324096 223038
rect 324044 222974 324096 222980
rect 324608 217410 324636 228822
rect 324884 228478 324912 231676
rect 324872 228472 324924 228478
rect 324872 228414 324924 228420
rect 325252 222494 325280 231676
rect 325620 223106 325648 231676
rect 325700 228336 325752 228342
rect 325700 228278 325752 228284
rect 325608 223100 325660 223106
rect 325608 223042 325660 223048
rect 325240 222488 325292 222494
rect 325240 222430 325292 222436
rect 325712 217410 325740 228278
rect 325988 227458 326016 231676
rect 326252 228132 326304 228138
rect 326252 228074 326304 228080
rect 325976 227452 326028 227458
rect 325976 227394 326028 227400
rect 326264 217410 326292 228074
rect 326356 223242 326384 231676
rect 326344 223236 326396 223242
rect 326344 223178 326396 223184
rect 326632 222970 326660 231676
rect 327000 223378 327028 231676
rect 327080 228608 327132 228614
rect 327080 228550 327132 228556
rect 326988 223372 327040 223378
rect 326988 223314 327040 223320
rect 326620 222964 326672 222970
rect 326620 222906 326672 222912
rect 327092 217410 327120 228550
rect 327368 222902 327396 231676
rect 327356 222896 327408 222902
rect 327356 222838 327408 222844
rect 327736 222426 327764 231676
rect 327908 226364 327960 226370
rect 327908 226306 327960 226312
rect 327724 222420 327776 222426
rect 327724 222362 327776 222368
rect 327920 217410 327948 226306
rect 328104 222766 328132 231676
rect 328472 223174 328500 231676
rect 328840 228682 328868 231676
rect 328828 228676 328880 228682
rect 328828 228618 328880 228624
rect 328828 228268 328880 228274
rect 328828 228210 328880 228216
rect 328460 223168 328512 223174
rect 328460 223110 328512 223116
rect 328092 222760 328144 222766
rect 328092 222702 328144 222708
rect 328840 217410 328868 228210
rect 329208 221066 329236 231676
rect 329484 222698 329512 231676
rect 329656 228200 329708 228206
rect 329656 228142 329708 228148
rect 329472 222692 329524 222698
rect 329472 222634 329524 222640
rect 329196 221060 329248 221066
rect 329196 221002 329248 221008
rect 329668 217410 329696 228142
rect 329852 221134 329880 231676
rect 330220 222834 330248 231676
rect 330484 228404 330536 228410
rect 330484 228346 330536 228352
rect 330208 222828 330260 222834
rect 330208 222770 330260 222776
rect 329840 221128 329892 221134
rect 329840 221070 329892 221076
rect 330496 217410 330524 228346
rect 330588 228342 330616 231676
rect 330576 228336 330628 228342
rect 330576 228278 330628 228284
rect 330956 222873 330984 231676
rect 331338 231662 331628 231690
rect 331312 227996 331364 228002
rect 331312 227938 331364 227944
rect 330942 222864 330998 222873
rect 330942 222799 330998 222808
rect 331324 217410 331352 227938
rect 331600 222630 331628 231662
rect 331692 227118 331720 231676
rect 332060 227662 332088 231676
rect 332140 228812 332192 228818
rect 332140 228754 332192 228760
rect 332048 227656 332100 227662
rect 332048 227598 332100 227604
rect 331680 227112 331732 227118
rect 331680 227054 331732 227060
rect 331588 222624 331640 222630
rect 331588 222566 331640 222572
rect 332152 217410 332180 228754
rect 332336 222601 332364 231676
rect 332704 223009 332732 231676
rect 332968 228064 333020 228070
rect 332968 228006 333020 228012
rect 332690 223000 332746 223009
rect 332690 222935 332746 222944
rect 332322 222592 332378 222601
rect 332322 222527 332378 222536
rect 332980 217410 333008 228006
rect 333072 227186 333100 231676
rect 333440 228274 333468 231676
rect 333428 228268 333480 228274
rect 333428 228210 333480 228216
rect 333060 227180 333112 227186
rect 333060 227122 333112 227128
rect 333808 222465 333836 231676
rect 333794 222456 333850 222465
rect 333794 222391 333850 222400
rect 333980 222352 334032 222358
rect 333980 222294 334032 222300
rect 333992 217410 334020 222294
rect 334176 220998 334204 231676
rect 334544 226574 334572 231676
rect 334912 228138 334940 231676
rect 334900 228132 334952 228138
rect 334900 228074 334952 228080
rect 334716 227928 334768 227934
rect 334716 227870 334768 227876
rect 334532 226568 334584 226574
rect 334532 226510 334584 226516
rect 334164 220992 334216 220998
rect 334164 220934 334216 220940
rect 334728 217410 334756 227870
rect 335188 224126 335216 231676
rect 335570 231662 335860 231690
rect 335544 227724 335596 227730
rect 335544 227666 335596 227672
rect 335176 224120 335228 224126
rect 335176 224062 335228 224068
rect 335556 217410 335584 227666
rect 335832 222737 335860 231662
rect 335818 222728 335874 222737
rect 335818 222663 335874 222672
rect 335924 222193 335952 231676
rect 336292 228070 336320 231676
rect 336660 228750 336688 231676
rect 337042 231662 337332 231690
rect 336648 228744 336700 228750
rect 336648 228686 336700 228692
rect 336280 228064 336332 228070
rect 336280 228006 336332 228012
rect 336740 222216 336792 222222
rect 335910 222184 335966 222193
rect 336740 222158 336792 222164
rect 335910 222119 335966 222128
rect 336752 217410 336780 222158
rect 337304 221202 337332 231662
rect 337396 222222 337424 231676
rect 337764 228614 337792 231676
rect 337752 228608 337804 228614
rect 337752 228550 337804 228556
rect 338040 228410 338068 231676
rect 338120 228540 338172 228546
rect 338120 228482 338172 228488
rect 338028 228404 338080 228410
rect 338028 228346 338080 228352
rect 338132 222290 338160 228482
rect 338408 227934 338436 231676
rect 338396 227928 338448 227934
rect 338396 227870 338448 227876
rect 338776 222329 338804 231676
rect 339144 228206 339172 231676
rect 339132 228200 339184 228206
rect 339132 228142 339184 228148
rect 338856 225072 338908 225078
rect 338856 225014 338908 225020
rect 338762 222320 338818 222329
rect 338028 222284 338080 222290
rect 338028 222226 338080 222232
rect 338120 222284 338172 222290
rect 338762 222255 338818 222264
rect 338120 222226 338172 222232
rect 337384 222216 337436 222222
rect 337384 222158 337436 222164
rect 337200 221196 337252 221202
rect 337200 221138 337252 221144
rect 337292 221196 337344 221202
rect 337292 221138 337344 221144
rect 317892 217382 318228 217410
rect 318720 217382 319056 217410
rect 319548 217382 319884 217410
rect 320376 217382 320712 217410
rect 321204 217382 321540 217410
rect 322032 217382 322368 217410
rect 322952 217382 323288 217410
rect 323780 217382 324116 217410
rect 324608 217382 324944 217410
rect 325712 217382 325772 217410
rect 326264 217382 326600 217410
rect 327092 217382 327428 217410
rect 327920 217382 328256 217410
rect 328840 217382 329176 217410
rect 329668 217382 330004 217410
rect 330496 217382 330832 217410
rect 331324 217382 331660 217410
rect 332152 217382 332488 217410
rect 332980 217382 333316 217410
rect 333992 217382 334144 217410
rect 334728 217382 335064 217410
rect 335556 217382 335892 217410
rect 336720 217382 336780 217410
rect 337212 217410 337240 221138
rect 338040 217410 338068 222226
rect 338868 217410 338896 225014
rect 339512 224194 339540 231676
rect 339776 227792 339828 227798
rect 339776 227734 339828 227740
rect 339500 224188 339552 224194
rect 339500 224130 339552 224136
rect 339788 222358 339816 227734
rect 339880 225486 339908 231676
rect 339868 225480 339920 225486
rect 339868 225422 339920 225428
rect 340248 224398 340276 231676
rect 340616 228886 340644 231676
rect 340604 228880 340656 228886
rect 340604 228822 340656 228828
rect 340892 228818 340920 231676
rect 340880 228812 340932 228818
rect 340880 228754 340932 228760
rect 341260 227866 341288 231676
rect 341248 227860 341300 227866
rect 341248 227802 341300 227808
rect 341628 227730 341656 231676
rect 341996 228546 342024 231676
rect 342364 228954 342392 231676
rect 342168 228948 342220 228954
rect 342168 228890 342220 228896
rect 342352 228948 342404 228954
rect 342352 228890 342404 228896
rect 341984 228540 342036 228546
rect 341984 228482 342036 228488
rect 341616 227724 341668 227730
rect 341616 227666 341668 227672
rect 340236 224392 340288 224398
rect 340236 224334 340288 224340
rect 339776 222352 339828 222358
rect 339776 222294 339828 222300
rect 340604 221604 340656 221610
rect 340604 221546 340656 221552
rect 339684 221400 339736 221406
rect 339684 221342 339736 221348
rect 339696 217410 339724 221342
rect 340616 217410 340644 221546
rect 342180 221270 342208 228890
rect 342732 228002 342760 231676
rect 342720 227996 342772 228002
rect 342720 227938 342772 227944
rect 342812 227384 342864 227390
rect 342812 227326 342864 227332
rect 342444 224936 342496 224942
rect 342444 224878 342496 224884
rect 341432 221264 341484 221270
rect 341432 221206 341484 221212
rect 342168 221264 342220 221270
rect 342168 221206 342220 221212
rect 341444 217410 341472 221206
rect 342456 217410 342484 224878
rect 342824 221406 342852 227326
rect 343100 224058 343128 231676
rect 343468 229022 343496 231676
rect 343456 229016 343508 229022
rect 343456 228958 343508 228964
rect 343744 224942 343772 231676
rect 344112 225078 344140 231676
rect 344480 225690 344508 231676
rect 344468 225684 344520 225690
rect 344468 225626 344520 225632
rect 344100 225072 344152 225078
rect 344100 225014 344152 225020
rect 343732 224936 343784 224942
rect 343732 224878 343784 224884
rect 343088 224052 343140 224058
rect 343088 223994 343140 224000
rect 343640 223440 343692 223446
rect 343468 223388 343640 223394
rect 343468 223382 343692 223388
rect 343468 223366 343680 223382
rect 343468 223310 343496 223366
rect 343456 223304 343508 223310
rect 343456 223246 343508 223252
rect 343548 223304 343600 223310
rect 343548 223246 343600 223252
rect 343560 223038 343588 223246
rect 343548 223032 343600 223038
rect 343548 222974 343600 222980
rect 343640 223032 343692 223038
rect 343640 222974 343692 222980
rect 343652 222562 343680 222974
rect 343640 222556 343692 222562
rect 343640 222498 343692 222504
rect 343732 222556 343784 222562
rect 343732 222498 343784 222504
rect 343548 222420 343600 222426
rect 343548 222362 343600 222368
rect 342812 221400 342864 221406
rect 342812 221342 342864 221348
rect 343088 221332 343140 221338
rect 343088 221274 343140 221280
rect 343100 217410 343128 221274
rect 343560 221066 343588 222362
rect 343744 221134 343772 222498
rect 343916 221468 343968 221474
rect 343916 221410 343968 221416
rect 343732 221128 343784 221134
rect 343732 221070 343784 221076
rect 343548 221060 343600 221066
rect 343548 221002 343600 221008
rect 343928 217410 343956 221410
rect 344848 219230 344876 231676
rect 345112 227452 345164 227458
rect 345112 227394 345164 227400
rect 345124 221542 345152 227394
rect 345216 226982 345244 231676
rect 345598 231662 345888 231690
rect 345388 228676 345440 228682
rect 345388 228618 345440 228624
rect 345296 227520 345348 227526
rect 345296 227462 345348 227468
rect 345204 226976 345256 226982
rect 345204 226918 345256 226924
rect 345020 221536 345072 221542
rect 345020 221478 345072 221484
rect 345112 221536 345164 221542
rect 345112 221478 345164 221484
rect 344836 219224 344888 219230
rect 344836 219166 344888 219172
rect 345032 217410 345060 221478
rect 345308 221474 345336 227462
rect 345400 221610 345428 228618
rect 345860 225010 345888 231662
rect 345952 227798 345980 231676
rect 345940 227792 345992 227798
rect 345940 227734 345992 227740
rect 345664 225004 345716 225010
rect 345664 224946 345716 224952
rect 345848 225004 345900 225010
rect 345848 224946 345900 224952
rect 345388 221604 345440 221610
rect 345388 221546 345440 221552
rect 345296 221468 345348 221474
rect 345296 221410 345348 221416
rect 345676 217410 345704 224946
rect 346320 219162 346348 231676
rect 346596 224534 346624 231676
rect 346584 224528 346636 224534
rect 346584 224470 346636 224476
rect 346964 224262 346992 231676
rect 347332 230110 347360 231676
rect 347320 230104 347372 230110
rect 347320 230046 347372 230052
rect 346952 224256 347004 224262
rect 346952 224198 347004 224204
rect 346492 222284 346544 222290
rect 346492 222226 346544 222232
rect 346308 219156 346360 219162
rect 346308 219098 346360 219104
rect 346504 217410 346532 222226
rect 346676 222216 346728 222222
rect 346676 222158 346728 222164
rect 346688 221202 346716 222158
rect 347320 221672 347372 221678
rect 347320 221614 347372 221620
rect 346676 221196 346728 221202
rect 346676 221138 346728 221144
rect 347332 217410 347360 221614
rect 347700 220794 347728 231676
rect 347780 227180 347832 227186
rect 347780 227122 347832 227128
rect 347792 223582 347820 227122
rect 347872 227112 347924 227118
rect 347872 227054 347924 227060
rect 347780 223576 347832 223582
rect 347780 223518 347832 223524
rect 347884 221270 347912 227054
rect 348068 224466 348096 231676
rect 348056 224460 348108 224466
rect 348056 224402 348108 224408
rect 348436 224330 348464 231676
rect 348804 230178 348832 231676
rect 348792 230172 348844 230178
rect 348792 230114 348844 230120
rect 348976 225208 349028 225214
rect 348976 225150 349028 225156
rect 348424 224324 348476 224330
rect 348424 224266 348476 224272
rect 348148 223644 348200 223650
rect 348148 223586 348200 223592
rect 347872 221264 347924 221270
rect 347872 221206 347924 221212
rect 347688 220788 347740 220794
rect 347688 220730 347740 220736
rect 348160 217410 348188 223586
rect 348988 217410 349016 225150
rect 349172 219366 349200 231676
rect 349448 224806 349476 231676
rect 349436 224800 349488 224806
rect 349436 224742 349488 224748
rect 349816 224602 349844 231676
rect 350184 230314 350212 231676
rect 350172 230308 350224 230314
rect 350172 230250 350224 230256
rect 349804 224596 349856 224602
rect 349804 224538 349856 224544
rect 349804 222352 349856 222358
rect 349804 222294 349856 222300
rect 349896 222352 349948 222358
rect 349896 222294 349948 222300
rect 349160 219360 349212 219366
rect 349160 219302 349212 219308
rect 349816 217410 349844 222294
rect 349908 220998 349936 222294
rect 349896 220992 349948 220998
rect 349896 220934 349948 220940
rect 350552 219298 350580 231676
rect 350920 224670 350948 231676
rect 350908 224664 350960 224670
rect 350908 224606 350960 224612
rect 350632 221876 350684 221882
rect 350632 221818 350684 221824
rect 350540 219292 350592 219298
rect 350540 219234 350592 219240
rect 350644 217410 350672 221818
rect 351288 220726 351316 231676
rect 351656 230246 351684 231676
rect 351644 230240 351696 230246
rect 351644 230182 351696 230188
rect 351920 226568 351972 226574
rect 351920 226510 351972 226516
rect 351460 221740 351512 221746
rect 351460 221682 351512 221688
rect 351276 220720 351328 220726
rect 351276 220662 351328 220668
rect 351472 217410 351500 221682
rect 351932 221678 351960 226510
rect 351920 221672 351972 221678
rect 351920 221614 351972 221620
rect 352024 220658 352052 231676
rect 352300 226234 352328 231676
rect 352288 226228 352340 226234
rect 352288 226170 352340 226176
rect 352380 225140 352432 225146
rect 352380 225082 352432 225088
rect 352012 220652 352064 220658
rect 352012 220594 352064 220600
rect 352392 217410 352420 225082
rect 352668 224738 352696 231676
rect 353036 227526 353064 231676
rect 353024 227520 353076 227526
rect 353024 227462 353076 227468
rect 352656 224732 352708 224738
rect 352656 224674 352708 224680
rect 353300 221196 353352 221202
rect 353300 221138 353352 221144
rect 353312 217410 353340 221138
rect 353404 220590 353432 231676
rect 353772 226302 353800 231676
rect 353760 226296 353812 226302
rect 353760 226238 353812 226244
rect 354140 224874 354168 231676
rect 354508 230042 354536 231676
rect 354890 231662 355088 231690
rect 354496 230036 354548 230042
rect 354496 229978 354548 229984
rect 354128 224868 354180 224874
rect 354128 224810 354180 224816
rect 354036 221944 354088 221950
rect 354036 221886 354088 221892
rect 353392 220584 353444 220590
rect 353392 220526 353444 220532
rect 354048 217410 354076 221886
rect 354864 221808 354916 221814
rect 354864 221750 354916 221756
rect 354876 217410 354904 221750
rect 355060 220454 355088 231662
rect 355152 226166 355180 231676
rect 355140 226160 355192 226166
rect 355140 226102 355192 226108
rect 355520 225554 355548 231676
rect 355888 229974 355916 231676
rect 355876 229968 355928 229974
rect 355876 229910 355928 229916
rect 356060 227588 356112 227594
rect 356060 227530 356112 227536
rect 355508 225548 355560 225554
rect 355508 225490 355560 225496
rect 355048 220448 355100 220454
rect 355048 220390 355100 220396
rect 356072 217410 356100 227530
rect 356256 220522 356284 231676
rect 356624 227594 356652 231676
rect 356612 227588 356664 227594
rect 356612 227530 356664 227536
rect 356992 225418 357020 231676
rect 357360 229906 357388 231676
rect 357348 229900 357400 229906
rect 357348 229842 357400 229848
rect 356980 225412 357032 225418
rect 356980 225354 357032 225360
rect 356520 222148 356572 222154
rect 356520 222090 356572 222096
rect 356244 220516 356296 220522
rect 356244 220458 356296 220464
rect 337212 217382 337548 217410
rect 338040 217382 338376 217410
rect 338868 217382 339204 217410
rect 339696 217382 340032 217410
rect 340616 217382 340952 217410
rect 341444 217382 341780 217410
rect 342456 217382 342608 217410
rect 343100 217382 343436 217410
rect 343928 217382 344264 217410
rect 345032 217382 345092 217410
rect 345676 217382 345920 217410
rect 346504 217382 346840 217410
rect 347332 217382 347668 217410
rect 348160 217382 348496 217410
rect 348988 217382 349324 217410
rect 349816 217382 350152 217410
rect 350644 217382 350980 217410
rect 351472 217382 351808 217410
rect 352392 217382 352728 217410
rect 353312 217382 353556 217410
rect 354048 217382 354384 217410
rect 354876 217382 355212 217410
rect 356040 217382 356100 217410
rect 356532 217410 356560 222090
rect 357348 222080 357400 222086
rect 357348 222022 357400 222028
rect 357360 217410 357388 222022
rect 357728 220318 357756 231676
rect 358004 225282 358032 231676
rect 358372 225350 358400 231676
rect 358740 227390 358768 231676
rect 359122 231662 359412 231690
rect 358728 227384 358780 227390
rect 358728 227326 358780 227332
rect 359096 227044 359148 227050
rect 359096 226986 359148 226992
rect 358360 225344 358412 225350
rect 358360 225286 358412 225292
rect 357992 225276 358044 225282
rect 357992 225218 358044 225224
rect 358268 222012 358320 222018
rect 358268 221954 358320 221960
rect 357716 220312 357768 220318
rect 357716 220254 357768 220260
rect 358280 217410 358308 221954
rect 359108 217410 359136 226986
rect 359384 220386 359412 231662
rect 359476 226098 359504 231676
rect 359844 226914 359872 231676
rect 360212 229838 360240 231676
rect 360200 229832 360252 229838
rect 360200 229774 360252 229780
rect 359832 226908 359884 226914
rect 359832 226850 359884 226856
rect 359464 226092 359516 226098
rect 359464 226034 359516 226040
rect 359924 221400 359976 221406
rect 359924 221342 359976 221348
rect 359372 220380 359424 220386
rect 359372 220322 359424 220328
rect 359936 217410 359964 221342
rect 360580 220182 360608 231676
rect 360856 225146 360884 231676
rect 361224 225214 361252 231676
rect 361592 227050 361620 231676
rect 361580 227044 361632 227050
rect 361580 226986 361632 226992
rect 361212 225208 361264 225214
rect 361212 225150 361264 225156
rect 360844 225140 360896 225146
rect 360844 225082 360896 225088
rect 360752 223508 360804 223514
rect 360752 223450 360804 223456
rect 360568 220176 360620 220182
rect 360568 220118 360620 220124
rect 360764 217410 360792 223450
rect 361764 223440 361816 223446
rect 361764 223382 361816 223388
rect 361776 217410 361804 223382
rect 361960 220250 361988 231676
rect 362328 226030 362356 231676
rect 362408 226840 362460 226846
rect 362408 226782 362460 226788
rect 362316 226024 362368 226030
rect 362316 225966 362368 225972
rect 361948 220244 362000 220250
rect 361948 220186 362000 220192
rect 362420 217410 362448 226782
rect 362696 225962 362724 231676
rect 363064 226846 363092 231676
rect 363052 226840 363104 226846
rect 363052 226782 363104 226788
rect 362684 225956 362736 225962
rect 362684 225898 362736 225904
rect 363236 221468 363288 221474
rect 363236 221410 363288 221416
rect 363248 217410 363276 221410
rect 363432 220046 363460 231676
rect 363708 225758 363736 231676
rect 364076 229770 364104 231676
rect 364064 229764 364116 229770
rect 364064 229706 364116 229712
rect 364444 227118 364472 231676
rect 364432 227112 364484 227118
rect 364432 227054 364484 227060
rect 363696 225752 363748 225758
rect 363696 225694 363748 225700
rect 364340 223304 364392 223310
rect 364340 223246 364392 223252
rect 363420 220040 363472 220046
rect 363420 219982 363472 219988
rect 364352 217410 364380 223246
rect 364812 220114 364840 231676
rect 365180 225826 365208 231676
rect 365548 229702 365576 231676
rect 365536 229696 365588 229702
rect 365536 229638 365588 229644
rect 365812 228472 365864 228478
rect 365812 228414 365864 228420
rect 365168 225820 365220 225826
rect 365168 225762 365220 225768
rect 364984 223100 365036 223106
rect 364984 223042 365036 223048
rect 364800 220108 364852 220114
rect 364800 220050 364852 220056
rect 364996 217410 365024 223042
rect 365824 217410 365852 228414
rect 365916 221406 365944 231676
rect 365904 221400 365956 221406
rect 365904 221342 365956 221348
rect 366284 219910 366312 231676
rect 366560 225622 366588 231676
rect 366928 225894 366956 231676
rect 367296 227186 367324 231676
rect 367284 227180 367336 227186
rect 367284 227122 367336 227128
rect 366916 225888 366968 225894
rect 366916 225830 366968 225836
rect 366548 225616 366600 225622
rect 366548 225558 366600 225564
rect 367468 223032 367520 223038
rect 367468 222974 367520 222980
rect 366640 221536 366692 221542
rect 366640 221478 366692 221484
rect 366272 219904 366324 219910
rect 366272 219846 366324 219852
rect 366652 217410 366680 221478
rect 367480 217410 367508 222974
rect 367664 219978 367692 231676
rect 368032 229090 368060 231676
rect 368400 229634 368428 231676
rect 368388 229628 368440 229634
rect 368388 229570 368440 229576
rect 368020 229084 368072 229090
rect 368020 229026 368072 229032
rect 368112 224052 368164 224058
rect 368112 223994 368164 224000
rect 368124 221134 368152 223994
rect 368296 223372 368348 223378
rect 368296 223314 368348 223320
rect 368112 221128 368164 221134
rect 368112 221070 368164 221076
rect 367652 219972 367704 219978
rect 367652 219914 367704 219920
rect 368308 217410 368336 223314
rect 368768 221474 368796 231676
rect 369150 231662 369348 231690
rect 369124 223236 369176 223242
rect 369124 223178 369176 223184
rect 368756 221468 368808 221474
rect 368756 221410 368808 221416
rect 369136 217410 369164 223178
rect 369320 219842 369348 231662
rect 369412 224505 369440 231676
rect 369596 231662 369794 231690
rect 369596 226710 369624 231662
rect 369768 229084 369820 229090
rect 369768 229026 369820 229032
rect 369676 227656 369728 227662
rect 369676 227598 369728 227604
rect 369584 226704 369636 226710
rect 369584 226646 369636 226652
rect 369584 225684 369636 225690
rect 369584 225626 369636 225632
rect 369398 224496 369454 224505
rect 369398 224431 369454 224440
rect 369596 221202 369624 225626
rect 369584 221196 369636 221202
rect 369584 221138 369636 221144
rect 369688 220930 369716 227598
rect 369780 225690 369808 229026
rect 370148 227254 370176 231676
rect 370516 229498 370544 231676
rect 370504 229492 370556 229498
rect 370504 229434 370556 229440
rect 370136 227248 370188 227254
rect 370136 227190 370188 227196
rect 369768 225684 369820 225690
rect 369768 225626 369820 225632
rect 370884 224641 370912 231676
rect 371252 229430 371280 231676
rect 371620 229566 371648 231676
rect 371608 229560 371660 229566
rect 371608 229502 371660 229508
rect 371240 229424 371292 229430
rect 371240 229366 371292 229372
rect 371516 226840 371568 226846
rect 371516 226782 371568 226788
rect 371240 225480 371292 225486
rect 371240 225422 371292 225428
rect 370870 224632 370926 224641
rect 370870 224567 370926 224576
rect 371148 224392 371200 224398
rect 371148 224334 371200 224340
rect 370872 222964 370924 222970
rect 370872 222906 370924 222912
rect 370044 222896 370096 222902
rect 370044 222838 370096 222844
rect 369676 220924 369728 220930
rect 369676 220866 369728 220872
rect 369308 219836 369360 219842
rect 369308 219778 369360 219784
rect 370056 217410 370084 222838
rect 370884 217410 370912 222906
rect 371160 222902 371188 224334
rect 371252 222970 371280 225422
rect 371240 222964 371292 222970
rect 371240 222906 371292 222912
rect 371148 222896 371200 222902
rect 371148 222838 371200 222844
rect 371528 221338 371556 226782
rect 371988 226778 372016 231676
rect 371976 226772 372028 226778
rect 371976 226714 372028 226720
rect 372264 226273 372292 231676
rect 372250 226264 372306 226273
rect 372250 226199 372306 226208
rect 372632 225486 372660 231676
rect 372896 227588 372948 227594
rect 372896 227530 372948 227536
rect 372620 225480 372672 225486
rect 372620 225422 372672 225428
rect 372908 224398 372936 227530
rect 373000 227458 373028 231676
rect 372988 227452 373040 227458
rect 372988 227394 373040 227400
rect 373368 226846 373396 231676
rect 373356 226840 373408 226846
rect 373356 226782 373408 226788
rect 373736 224777 373764 231676
rect 374104 229362 374132 231676
rect 374092 229356 374144 229362
rect 374092 229298 374144 229304
rect 373722 224768 373778 224777
rect 373722 224703 373778 224712
rect 372896 224392 372948 224398
rect 372896 224334 372948 224340
rect 371700 223168 371752 223174
rect 371700 223110 371752 223116
rect 371516 221332 371568 221338
rect 371516 221274 371568 221280
rect 371712 217410 371740 223110
rect 374184 222760 374236 222766
rect 374184 222702 374236 222708
rect 372620 222488 372672 222494
rect 372620 222430 372672 222436
rect 372632 217410 372660 222430
rect 373356 221604 373408 221610
rect 373356 221546 373408 221552
rect 373368 217410 373396 221546
rect 374196 217410 374224 222702
rect 374472 221542 374500 231676
rect 374840 227322 374868 231676
rect 374828 227316 374880 227322
rect 374828 227258 374880 227264
rect 375116 222057 375144 231676
rect 375380 222556 375432 222562
rect 375380 222498 375432 222504
rect 375102 222048 375158 222057
rect 375102 221983 375158 221992
rect 374460 221536 374512 221542
rect 374460 221478 374512 221484
rect 375392 217410 375420 222498
rect 375484 221610 375512 231676
rect 375852 227225 375880 231676
rect 376220 229294 376248 231676
rect 376208 229288 376260 229294
rect 376208 229230 376260 229236
rect 376588 228682 376616 231676
rect 376576 228676 376628 228682
rect 376576 228618 376628 228624
rect 375838 227216 375894 227225
rect 375838 227151 375894 227160
rect 376668 226976 376720 226982
rect 376668 226918 376720 226924
rect 376680 224058 376708 226918
rect 376668 224052 376720 224058
rect 376668 223994 376720 224000
rect 376956 223553 376984 231676
rect 376942 223544 376998 223553
rect 376942 223479 376998 223488
rect 377324 223417 377352 231676
rect 377310 223408 377366 223417
rect 377310 223343 377366 223352
rect 376760 222828 376812 222834
rect 376760 222770 376812 222776
rect 375932 222420 375984 222426
rect 375932 222362 375984 222368
rect 375472 221604 375524 221610
rect 375472 221546 375524 221552
rect 356532 217382 356868 217410
rect 357360 217382 357696 217410
rect 358280 217382 358616 217410
rect 359108 217382 359444 217410
rect 359936 217382 360272 217410
rect 360764 217382 361100 217410
rect 361776 217382 361928 217410
rect 362420 217382 362756 217410
rect 363248 217382 363584 217410
rect 364352 217382 364504 217410
rect 364996 217382 365332 217410
rect 365824 217382 366160 217410
rect 366652 217382 366988 217410
rect 367480 217382 367816 217410
rect 368308 217382 368644 217410
rect 369136 217382 369472 217410
rect 370056 217382 370392 217410
rect 370884 217382 371220 217410
rect 371712 217382 372048 217410
rect 372632 217382 372876 217410
rect 373368 217382 373704 217410
rect 374196 217382 374532 217410
rect 375360 217382 375420 217410
rect 375944 217410 375972 222362
rect 376772 217410 376800 222770
rect 377588 222692 377640 222698
rect 377588 222634 377640 222640
rect 377600 217410 377628 222634
rect 377692 221746 377720 231676
rect 377968 221882 377996 231676
rect 378140 228404 378192 228410
rect 378140 228346 378192 228352
rect 378152 222426 378180 228346
rect 378336 227361 378364 231676
rect 378322 227352 378378 227361
rect 378322 227287 378378 227296
rect 378704 226574 378732 231676
rect 379072 226982 379100 231676
rect 379244 228336 379296 228342
rect 379244 228278 379296 228284
rect 379060 226976 379112 226982
rect 379060 226918 379112 226924
rect 378692 226568 378744 226574
rect 378692 226510 378744 226516
rect 378416 222624 378468 222630
rect 378416 222566 378468 222572
rect 378140 222420 378192 222426
rect 378140 222362 378192 222368
rect 377956 221876 378008 221882
rect 377956 221818 378008 221824
rect 377680 221740 377732 221746
rect 377680 221682 377732 221688
rect 378428 217410 378456 222566
rect 379256 217410 379284 228278
rect 379440 221814 379468 231676
rect 379808 223281 379836 231676
rect 379794 223272 379850 223281
rect 379794 223207 379850 223216
rect 380176 223145 380204 231676
rect 380162 223136 380218 223145
rect 380162 223071 380218 223080
rect 380544 222018 380572 231676
rect 380820 228478 380848 231676
rect 381084 229016 381136 229022
rect 381084 228958 381136 228964
rect 380992 228744 381044 228750
rect 380992 228686 381044 228692
rect 380808 228472 380860 228478
rect 380808 228414 380860 228420
rect 381004 222562 381032 228686
rect 381096 226334 381124 228958
rect 381188 227497 381216 231676
rect 381556 228857 381584 231676
rect 381542 228848 381598 228857
rect 381542 228783 381598 228792
rect 381924 227662 381952 231676
rect 381912 227656 381964 227662
rect 381912 227598 381964 227604
rect 381174 227488 381230 227497
rect 381174 227423 381230 227432
rect 381096 226306 381216 226334
rect 381082 222864 381138 222873
rect 381082 222799 381138 222808
rect 380992 222556 381044 222562
rect 380992 222498 381044 222504
rect 380532 222012 380584 222018
rect 380532 221954 380584 221960
rect 379428 221808 379480 221814
rect 379428 221750 379480 221756
rect 380072 221264 380124 221270
rect 380072 221206 380124 221212
rect 380084 217410 380112 221206
rect 381096 217410 381124 222799
rect 381188 220998 381216 226306
rect 381818 223000 381874 223009
rect 381818 222935 381874 222944
rect 381176 220992 381228 220998
rect 381176 220934 381228 220940
rect 381832 217410 381860 222935
rect 382292 222494 382320 231676
rect 382660 222873 382688 231676
rect 382646 222864 382702 222873
rect 382646 222799 382702 222808
rect 382280 222488 382332 222494
rect 382280 222430 382332 222436
rect 383028 222154 383056 231676
rect 383396 228410 383424 231676
rect 383672 228993 383700 231676
rect 383658 228984 383714 228993
rect 383658 228919 383714 228928
rect 383752 228948 383804 228954
rect 383752 228890 383804 228896
rect 383660 228812 383712 228818
rect 383660 228754 383712 228760
rect 383384 228404 383436 228410
rect 383384 228346 383436 228352
rect 383672 223922 383700 228754
rect 383764 223990 383792 228890
rect 383844 228608 383896 228614
rect 383844 228550 383896 228556
rect 383752 223984 383804 223990
rect 383752 223926 383804 223932
rect 383660 223916 383712 223922
rect 383660 223858 383712 223864
rect 383660 223576 383712 223582
rect 383660 223518 383712 223524
rect 383016 222148 383068 222154
rect 383016 222090 383068 222096
rect 382648 220924 382700 220930
rect 382648 220866 382700 220872
rect 382660 217410 382688 220866
rect 383672 217410 383700 223518
rect 383856 221678 383884 228550
rect 384040 227594 384068 231676
rect 384028 227588 384080 227594
rect 384028 227530 384080 227536
rect 384302 222592 384358 222601
rect 384302 222527 384358 222536
rect 383752 221672 383804 221678
rect 383752 221614 383804 221620
rect 383844 221672 383896 221678
rect 383844 221614 383896 221620
rect 383764 221270 383792 221614
rect 383752 221264 383804 221270
rect 383752 221206 383804 221212
rect 384316 217410 384344 222527
rect 384408 222086 384436 231676
rect 384776 223009 384804 231676
rect 385158 231662 385448 231690
rect 385224 228880 385276 228886
rect 385224 228822 385276 228828
rect 384762 223000 384818 223009
rect 384762 222935 384818 222944
rect 385236 222358 385264 228822
rect 385132 222352 385184 222358
rect 385132 222294 385184 222300
rect 385224 222352 385276 222358
rect 385224 222294 385276 222300
rect 384396 222080 384448 222086
rect 384396 222022 384448 222028
rect 385144 217410 385172 222294
rect 385420 220862 385448 231662
rect 385512 228342 385540 231676
rect 385880 228721 385908 231676
rect 386248 229090 386276 231676
rect 386236 229084 386288 229090
rect 386236 229026 386288 229032
rect 385866 228712 385922 228721
rect 385866 228647 385922 228656
rect 385500 228336 385552 228342
rect 385500 228278 385552 228284
rect 385960 228268 386012 228274
rect 385960 228210 386012 228216
rect 385408 220856 385460 220862
rect 385408 220798 385460 220804
rect 385972 217410 386000 228210
rect 386524 223582 386552 231676
rect 386512 223576 386564 223582
rect 386512 223518 386564 223524
rect 386892 221785 386920 231676
rect 387260 223446 387288 231676
rect 387628 228274 387656 231676
rect 387996 228585 388024 231676
rect 388364 228614 388392 231676
rect 388732 228954 388760 231676
rect 388720 228948 388772 228954
rect 388720 228890 388772 228896
rect 388352 228608 388404 228614
rect 387982 228576 388038 228585
rect 388352 228550 388404 228556
rect 387982 228511 388038 228520
rect 389100 228449 389128 231676
rect 389086 228440 389142 228449
rect 389086 228375 389142 228384
rect 387616 228268 387668 228274
rect 387616 228210 387668 228216
rect 389088 228132 389140 228138
rect 389088 228074 389140 228080
rect 388996 228064 389048 228070
rect 388996 228006 389048 228012
rect 387524 226976 387576 226982
rect 387524 226918 387576 226924
rect 387248 223440 387300 223446
rect 387248 223382 387300 223388
rect 387536 221950 387564 226918
rect 388534 222728 388590 222737
rect 388534 222663 388590 222672
rect 387706 222456 387762 222465
rect 387706 222391 387762 222400
rect 387524 221944 387576 221950
rect 387524 221886 387576 221892
rect 386878 221776 386934 221785
rect 386878 221711 386934 221720
rect 386788 221264 386840 221270
rect 386788 221206 386840 221212
rect 386800 217410 386828 221206
rect 387720 217410 387748 222391
rect 388548 217410 388576 222663
rect 389008 221270 389036 228006
rect 388996 221264 389048 221270
rect 388996 221206 389048 221212
rect 389100 221082 389128 228074
rect 389376 226506 389404 231676
rect 389364 226500 389416 226506
rect 389364 226442 389416 226448
rect 389744 223378 389772 231676
rect 389732 223372 389784 223378
rect 389732 223314 389784 223320
rect 390112 222737 390140 231676
rect 390480 225729 390508 231676
rect 390848 228818 390876 231676
rect 390836 228812 390888 228818
rect 390836 228754 390888 228760
rect 391216 228313 391244 231676
rect 391202 228304 391258 228313
rect 391202 228239 391258 228248
rect 390466 225720 390522 225729
rect 390466 225655 390522 225664
rect 391584 225457 391612 231676
rect 391848 228200 391900 228206
rect 391848 228142 391900 228148
rect 391570 225448 391626 225457
rect 391570 225383 391626 225392
rect 391020 224120 391072 224126
rect 391020 224062 391072 224068
rect 390098 222728 390154 222737
rect 390098 222663 390154 222672
rect 390190 222184 390246 222193
rect 390190 222119 390246 222128
rect 389100 221054 389312 221082
rect 389284 217410 389312 221054
rect 390204 217410 390232 222119
rect 391032 217410 391060 224062
rect 391860 220930 391888 228142
rect 391952 223310 391980 231676
rect 391940 223304 391992 223310
rect 391940 223246 391992 223252
rect 392228 222601 392256 231676
rect 392596 225593 392624 231676
rect 392964 228886 392992 231676
rect 392952 228880 393004 228886
rect 392952 228822 393004 228828
rect 393332 228177 393360 231676
rect 393700 229226 393728 231676
rect 393688 229220 393740 229226
rect 393688 229162 393740 229168
rect 393318 228168 393374 228177
rect 393318 228103 393374 228112
rect 392582 225584 392638 225593
rect 392582 225519 392638 225528
rect 394068 223242 394096 231676
rect 394056 223236 394108 223242
rect 394056 223178 394108 223184
rect 392214 222592 392270 222601
rect 392214 222527 392270 222536
rect 393596 222284 393648 222290
rect 393596 222226 393648 222232
rect 391940 222216 391992 222222
rect 391940 222158 391992 222164
rect 391848 220924 391900 220930
rect 391848 220866 391900 220872
rect 391952 217410 391980 222158
rect 392676 221264 392728 221270
rect 392676 221206 392728 221212
rect 392688 217410 392716 221206
rect 393608 217410 393636 222226
rect 394436 222193 394464 231676
rect 394608 228540 394660 228546
rect 394608 228482 394660 228488
rect 394620 222290 394648 228482
rect 394804 226438 394832 231676
rect 395080 229022 395108 231676
rect 395068 229016 395120 229022
rect 395068 228958 395120 228964
rect 395160 227996 395212 228002
rect 395160 227938 395212 227944
rect 394792 226432 394844 226438
rect 394792 226374 394844 226380
rect 394792 224188 394844 224194
rect 394792 224130 394844 224136
rect 394700 222556 394752 222562
rect 394700 222498 394752 222504
rect 394608 222284 394660 222290
rect 394608 222226 394660 222232
rect 394422 222184 394478 222193
rect 394422 222119 394478 222128
rect 394712 217410 394740 222498
rect 394804 220998 394832 224130
rect 395172 223854 395200 227938
rect 395252 227928 395304 227934
rect 395448 227905 395476 231676
rect 395252 227870 395304 227876
rect 395434 227896 395490 227905
rect 395160 223848 395212 223854
rect 395160 223790 395212 223796
rect 394792 220992 394844 220998
rect 394792 220934 394844 220940
rect 395264 217410 395292 227870
rect 395434 227831 395490 227840
rect 395816 226642 395844 231676
rect 395988 226840 396040 226846
rect 395988 226782 396040 226788
rect 395804 226636 395856 226642
rect 395804 226578 395856 226584
rect 396000 224369 396028 226782
rect 395986 224360 396042 224369
rect 395986 224295 396042 224304
rect 396184 223174 396212 231676
rect 396172 223168 396224 223174
rect 396172 223110 396224 223116
rect 396264 222488 396316 222494
rect 396552 222465 396580 231676
rect 396920 229158 396948 231676
rect 396908 229152 396960 229158
rect 396908 229094 396960 229100
rect 397288 228750 397316 231676
rect 397276 228744 397328 228750
rect 397276 228686 397328 228692
rect 397656 228041 397684 231676
rect 397642 228032 397698 228041
rect 397642 227967 397698 227976
rect 397644 227860 397696 227866
rect 397644 227802 397696 227808
rect 397460 226568 397512 226574
rect 397460 226510 397512 226516
rect 396264 222430 396316 222436
rect 396538 222456 396594 222465
rect 396276 221950 396304 222430
rect 396538 222391 396594 222400
rect 396906 222320 396962 222329
rect 396906 222255 396962 222264
rect 396172 221944 396224 221950
rect 396172 221886 396224 221892
rect 396264 221944 396316 221950
rect 396264 221886 396316 221892
rect 396184 221678 396212 221886
rect 396080 221672 396132 221678
rect 396080 221614 396132 221620
rect 396172 221672 396224 221678
rect 396172 221614 396224 221620
rect 396092 217410 396120 221614
rect 396920 217410 396948 222255
rect 397472 221921 397500 226510
rect 397656 222222 397684 227802
rect 397932 225321 397960 231676
rect 397918 225312 397974 225321
rect 397918 225247 397974 225256
rect 398300 223038 398328 231676
rect 398668 223106 398696 231676
rect 399036 226982 399064 231676
rect 399404 228206 399432 231676
rect 399392 228200 399444 228206
rect 399392 228142 399444 228148
rect 399024 226976 399076 226982
rect 399024 226918 399076 226924
rect 398656 223100 398708 223106
rect 398656 223042 398708 223048
rect 398288 223032 398340 223038
rect 398288 222974 398340 222980
rect 399772 222970 399800 231676
rect 400140 225185 400168 231676
rect 400508 228070 400536 231676
rect 400496 228064 400548 228070
rect 400496 228006 400548 228012
rect 400784 226914 400812 231676
rect 400220 226908 400272 226914
rect 400220 226850 400272 226856
rect 400772 226908 400824 226914
rect 400772 226850 400824 226856
rect 400126 225176 400182 225185
rect 400126 225111 400182 225120
rect 400232 224126 400260 226850
rect 400404 226772 400456 226778
rect 400404 226714 400456 226720
rect 400416 226334 400444 226714
rect 401152 226574 401180 231676
rect 401140 226568 401192 226574
rect 401140 226510 401192 226516
rect 400416 226306 400536 226334
rect 400220 224120 400272 224126
rect 400220 224062 400272 224068
rect 398564 222964 398616 222970
rect 398564 222906 398616 222912
rect 399760 222964 399812 222970
rect 399760 222906 399812 222912
rect 397736 222420 397788 222426
rect 397736 222362 397788 222368
rect 397644 222216 397696 222222
rect 397644 222158 397696 222164
rect 397458 221912 397514 221921
rect 397458 221847 397514 221856
rect 397748 217410 397776 222362
rect 398576 217410 398604 222906
rect 400404 222896 400456 222902
rect 400404 222838 400456 222844
rect 399484 220924 399536 220930
rect 399484 220866 399536 220872
rect 399496 217410 399524 220866
rect 400416 217410 400444 222838
rect 400508 220930 400536 226306
rect 401520 222834 401548 231676
rect 401888 222902 401916 231676
rect 402152 227724 402204 227730
rect 402152 227666 402204 227672
rect 401876 222896 401928 222902
rect 401876 222838 401928 222844
rect 401508 222828 401560 222834
rect 401508 222770 401560 222776
rect 401968 222216 402020 222222
rect 401968 222158 402020 222164
rect 401140 220992 401192 220998
rect 401140 220934 401192 220940
rect 400496 220924 400548 220930
rect 400496 220866 400548 220872
rect 401152 217410 401180 220934
rect 401980 217410 402008 222158
rect 402164 221270 402192 227666
rect 402256 222766 402284 231676
rect 402624 228002 402652 231676
rect 402612 227996 402664 228002
rect 402612 227938 402664 227944
rect 402992 227769 403020 231676
rect 402978 227760 403034 227769
rect 402978 227695 403034 227704
rect 402980 226704 403032 226710
rect 402980 226646 403032 226652
rect 402992 224194 403020 226646
rect 403360 225049 403388 231676
rect 403346 225040 403402 225049
rect 403346 224975 403402 224984
rect 402980 224188 403032 224194
rect 402980 224130 403032 224136
rect 402244 222760 402296 222766
rect 402244 222702 402296 222708
rect 403636 222698 403664 231676
rect 403624 222692 403676 222698
rect 403624 222634 403676 222640
rect 404004 222562 404032 231676
rect 404372 224913 404400 231676
rect 404740 227934 404768 231676
rect 404728 227928 404780 227934
rect 404728 227870 404780 227876
rect 405108 227633 405136 231676
rect 405094 227624 405150 227633
rect 405094 227559 405150 227568
rect 405476 226778 405504 231676
rect 405464 226772 405516 226778
rect 405464 226714 405516 226720
rect 404358 224904 404414 224913
rect 404358 224839 404414 224848
rect 404452 223916 404504 223922
rect 404452 223858 404504 223864
rect 403992 222556 404044 222562
rect 403992 222498 404044 222504
rect 402980 222352 403032 222358
rect 402980 222294 403032 222300
rect 402152 221264 402204 221270
rect 402152 221206 402204 221212
rect 402992 217410 403020 222294
rect 403624 221264 403676 221270
rect 403624 221206 403676 221212
rect 403636 217410 403664 221206
rect 404464 217410 404492 223858
rect 405740 223848 405792 223854
rect 405740 223790 405792 223796
rect 405752 217410 405780 223790
rect 405844 222630 405872 231676
rect 405832 222624 405884 222630
rect 405832 222566 405884 222572
rect 406212 222426 406240 231676
rect 406488 222494 406516 231676
rect 406856 227866 406884 231676
rect 407224 228138 407252 231676
rect 407212 228132 407264 228138
rect 407212 228074 407264 228080
rect 406844 227860 406896 227866
rect 406844 227802 406896 227808
rect 407592 226846 407620 231676
rect 407580 226840 407632 226846
rect 407580 226782 407632 226788
rect 407856 223984 407908 223990
rect 407856 223926 407908 223932
rect 406476 222488 406528 222494
rect 406476 222430 406528 222436
rect 406200 222420 406252 222426
rect 406200 222362 406252 222368
rect 406200 222284 406252 222290
rect 406200 222226 406252 222232
rect 375944 217382 376280 217410
rect 376772 217382 377108 217410
rect 377600 217382 377936 217410
rect 378428 217382 378764 217410
rect 379256 217382 379592 217410
rect 380084 217382 380420 217410
rect 381096 217382 381248 217410
rect 381832 217382 382168 217410
rect 382660 217382 382996 217410
rect 383672 217382 383824 217410
rect 384316 217382 384652 217410
rect 385144 217382 385480 217410
rect 385972 217382 386308 217410
rect 386800 217382 387136 217410
rect 387720 217382 388056 217410
rect 388548 217382 388884 217410
rect 389284 217382 389712 217410
rect 390204 217382 390540 217410
rect 391032 217382 391368 217410
rect 391952 217382 392196 217410
rect 392688 217382 393024 217410
rect 393608 217382 393944 217410
rect 394712 217382 394772 217410
rect 395264 217382 395600 217410
rect 396092 217382 396428 217410
rect 396920 217382 397256 217410
rect 397748 217382 398084 217410
rect 398576 217382 398912 217410
rect 399496 217382 399832 217410
rect 400416 217382 400660 217410
rect 401152 217382 401488 217410
rect 401980 217382 402316 217410
rect 402992 217382 403144 217410
rect 403636 217382 403972 217410
rect 404464 217382 404800 217410
rect 405720 217382 405780 217410
rect 406212 217410 406240 222226
rect 407028 221128 407080 221134
rect 407028 221070 407080 221076
rect 407040 217410 407068 221070
rect 407868 217410 407896 223926
rect 407960 222426 407988 231676
rect 408144 231662 408342 231690
rect 408710 231662 409000 231690
rect 407948 222420 408000 222426
rect 407948 222362 408000 222368
rect 408144 222290 408172 231662
rect 408316 228608 408368 228614
rect 408316 228550 408368 228556
rect 408224 227792 408276 227798
rect 408224 227734 408276 227740
rect 408236 223650 408264 227734
rect 408328 226137 408356 228550
rect 408408 226500 408460 226506
rect 408408 226442 408460 226448
rect 408314 226128 408370 226137
rect 408314 226063 408370 226072
rect 408420 226001 408448 226442
rect 408406 225992 408462 226001
rect 408406 225927 408462 225936
rect 408972 225078 409000 231662
rect 409064 228546 409092 231676
rect 409052 228540 409104 228546
rect 409052 228482 409104 228488
rect 409340 227798 409368 231676
rect 409328 227792 409380 227798
rect 409328 227734 409380 227740
rect 409708 226710 409736 231676
rect 410076 227089 410104 231676
rect 410444 227730 410472 231676
rect 410826 231662 411116 231690
rect 410892 228608 410944 228614
rect 410892 228550 410944 228556
rect 410432 227724 410484 227730
rect 410432 227666 410484 227672
rect 410062 227080 410118 227089
rect 410062 227015 410118 227024
rect 409696 226704 409748 226710
rect 409696 226646 409748 226652
rect 408684 225072 408736 225078
rect 408684 225014 408736 225020
rect 408960 225072 409012 225078
rect 408960 225014 409012 225020
rect 408224 223644 408276 223650
rect 408224 223586 408276 223592
rect 408132 222284 408184 222290
rect 408132 222226 408184 222232
rect 408696 217410 408724 225014
rect 410800 225004 410852 225010
rect 410800 224946 410852 224952
rect 409696 224596 409748 224602
rect 409696 224538 409748 224544
rect 409604 224528 409656 224534
rect 409604 224470 409656 224476
rect 409616 223786 409644 224470
rect 409708 224058 409736 224538
rect 410812 224466 410840 224946
rect 410800 224460 410852 224466
rect 410800 224402 410852 224408
rect 409696 224052 409748 224058
rect 409696 223994 409748 224000
rect 409604 223780 409656 223786
rect 409604 223722 409656 223728
rect 409786 222728 409842 222737
rect 409786 222663 409842 222672
rect 409800 221785 409828 222663
rect 410904 222222 410932 228550
rect 410984 227520 411036 227526
rect 410984 227462 411036 227468
rect 410996 223854 411024 227462
rect 411088 224942 411116 231662
rect 411180 228614 411208 231676
rect 411168 228608 411220 228614
rect 411168 228550 411220 228556
rect 411168 226432 411220 226438
rect 411168 226374 411220 226380
rect 411180 225865 411208 226374
rect 411166 225856 411222 225865
rect 411166 225791 411222 225800
rect 411548 225010 411576 231676
rect 411168 225004 411220 225010
rect 411168 224946 411220 224952
rect 411536 225004 411588 225010
rect 411536 224946 411588 224952
rect 411076 224936 411128 224942
rect 411076 224878 411128 224884
rect 410984 223848 411036 223854
rect 410984 223790 411036 223796
rect 410892 222216 410944 222222
rect 410892 222158 410944 222164
rect 409786 221776 409842 221785
rect 409786 221711 409842 221720
rect 410340 221196 410392 221202
rect 410340 221138 410392 221144
rect 409512 221060 409564 221066
rect 409512 221002 409564 221008
rect 409524 217410 409552 221002
rect 410352 217410 410380 221138
rect 411180 220946 411208 224946
rect 411916 221202 411944 231676
rect 417148 230104 417200 230110
rect 417148 230046 417200 230052
rect 415308 227384 415360 227390
rect 415308 227326 415360 227332
rect 412088 224460 412140 224466
rect 412088 224402 412140 224408
rect 411904 221196 411956 221202
rect 411904 221138 411956 221144
rect 411180 220918 411300 220946
rect 411272 217410 411300 220918
rect 412100 217410 412128 224402
rect 414572 223984 414624 223990
rect 414572 223926 414624 223932
rect 414020 223644 414072 223650
rect 414020 223586 414072 223592
rect 412916 219224 412968 219230
rect 412916 219166 412968 219172
rect 412928 217410 412956 219166
rect 414032 217410 414060 223586
rect 414584 217410 414612 223926
rect 415320 223922 415348 227326
rect 416780 227112 416832 227118
rect 416780 227054 416832 227060
rect 415492 227044 415544 227050
rect 415492 226986 415544 226992
rect 415504 224262 415532 226986
rect 416792 224534 416820 227054
rect 416780 224528 416832 224534
rect 416780 224470 416832 224476
rect 415400 224256 415452 224262
rect 415400 224198 415452 224204
rect 415492 224256 415544 224262
rect 415492 224198 415544 224204
rect 415308 223916 415360 223922
rect 415308 223858 415360 223864
rect 415412 217410 415440 224198
rect 416228 219156 416280 219162
rect 416228 219098 416280 219104
rect 416240 217410 416268 219098
rect 417160 217410 417188 230046
rect 417332 228540 417384 228546
rect 417332 228482 417384 228488
rect 417344 228138 417372 228482
rect 417332 228132 417384 228138
rect 417332 228074 417384 228080
rect 417516 228064 417568 228070
rect 417516 228006 417568 228012
rect 417528 226914 417556 228006
rect 417516 226908 417568 226914
rect 417516 226850 417568 226856
rect 417700 226840 417752 226846
rect 417700 226782 417752 226788
rect 417712 226574 417740 226782
rect 417700 226568 417752 226574
rect 417700 226510 417752 226516
rect 418080 226334 418108 243063
rect 418158 240000 418214 240009
rect 418158 239935 418214 239944
rect 417896 226306 418108 226334
rect 406212 217382 406548 217410
rect 407040 217382 407376 217410
rect 407868 217382 408204 217410
rect 408696 217382 409032 217410
rect 409524 217382 409860 217410
rect 410352 217382 410688 217410
rect 411272 217382 411608 217410
rect 412100 217382 412436 217410
rect 412928 217382 413264 217410
rect 414032 217382 414092 217410
rect 414584 217382 414920 217410
rect 415412 217382 415748 217410
rect 416240 217382 416576 217410
rect 417160 217382 417496 217410
rect 59452 216708 59504 216714
rect 59452 216650 59504 216656
rect 417896 216646 417924 226306
rect 417976 223780 418028 223786
rect 417976 223722 418028 223728
rect 417988 217410 418016 223722
rect 418172 218006 418200 239935
rect 418434 236736 418490 236745
rect 418434 236671 418490 236680
rect 418160 218000 418212 218006
rect 418160 217942 418212 217948
rect 417988 217382 418324 217410
rect 418448 216782 418476 236671
rect 418526 233608 418582 233617
rect 418526 233543 418582 233552
rect 418540 216850 418568 233543
rect 423864 230308 423916 230314
rect 423864 230250 423916 230256
rect 420460 230172 420512 230178
rect 420460 230114 420512 230120
rect 418804 224324 418856 224330
rect 418804 224266 418856 224272
rect 418620 218000 418672 218006
rect 418620 217942 418672 217948
rect 418528 216844 418580 216850
rect 418528 216786 418580 216792
rect 418436 216776 418488 216782
rect 418436 216718 418488 216724
rect 418632 216714 418660 217942
rect 418816 217410 418844 224266
rect 419724 220788 419776 220794
rect 419724 220730 419776 220736
rect 419736 217410 419764 220730
rect 420472 217410 420500 230114
rect 422300 227180 422352 227186
rect 422300 227122 422352 227128
rect 422312 224602 422340 227122
rect 421288 224596 421340 224602
rect 421288 224538 421340 224544
rect 422300 224596 422352 224602
rect 422300 224538 422352 224544
rect 421300 217410 421328 224538
rect 422300 224052 422352 224058
rect 422300 223994 422352 224000
rect 422312 217410 422340 223994
rect 423036 219360 423088 219366
rect 423036 219302 423088 219308
rect 423048 217410 423076 219302
rect 423876 217410 423904 230250
rect 427176 230240 427228 230246
rect 427176 230182 427228 230188
rect 425060 224800 425112 224806
rect 425060 224742 425112 224748
rect 425072 217410 425100 224742
rect 425520 220720 425572 220726
rect 425520 220662 425572 220668
rect 418816 217382 419152 217410
rect 419736 217382 419980 217410
rect 420472 217382 420808 217410
rect 421300 217382 421636 217410
rect 422312 217382 422464 217410
rect 423048 217382 423384 217410
rect 423876 217382 424212 217410
rect 425040 217382 425100 217410
rect 425532 217410 425560 220662
rect 426348 219292 426400 219298
rect 426348 219234 426400 219240
rect 426360 217410 426388 219234
rect 427188 217410 427216 230182
rect 433892 230036 433944 230042
rect 433892 229978 433944 229984
rect 433156 227452 433208 227458
rect 433156 227394 433208 227400
rect 428372 227248 428424 227254
rect 428372 227190 428424 227196
rect 428384 224806 428412 227190
rect 431408 226228 431460 226234
rect 431408 226170 431460 226176
rect 429016 225344 429068 225350
rect 429016 225286 429068 225292
rect 428372 224800 428424 224806
rect 428372 224742 428424 224748
rect 429028 224738 429056 225286
rect 428924 224732 428976 224738
rect 428924 224674 428976 224680
rect 429016 224732 429068 224738
rect 429016 224674 429068 224680
rect 428004 224664 428056 224670
rect 428004 224606 428056 224612
rect 428016 217410 428044 224606
rect 428936 217410 428964 224674
rect 430580 223848 430632 223854
rect 430580 223790 430632 223796
rect 429752 220652 429804 220658
rect 429752 220594 429804 220600
rect 429764 217410 429792 220594
rect 430592 217410 430620 223790
rect 431420 217410 431448 226170
rect 433168 224874 433196 227394
rect 433248 227316 433300 227322
rect 433248 227258 433300 227264
rect 433260 226234 433288 227258
rect 433248 226228 433300 226234
rect 433248 226170 433300 226176
rect 433524 225548 433576 225554
rect 433524 225490 433576 225496
rect 432236 224868 432288 224874
rect 432236 224810 432288 224816
rect 433156 224868 433208 224874
rect 433156 224810 433208 224816
rect 432248 217410 432276 224810
rect 433536 223650 433564 225490
rect 433524 223644 433576 223650
rect 433524 223586 433576 223592
rect 433340 220584 433392 220590
rect 433340 220526 433392 220532
rect 433352 217410 433380 220526
rect 433904 217410 433932 229978
rect 437296 229968 437348 229974
rect 437296 229910 437348 229916
rect 434628 226636 434680 226642
rect 434628 226578 434680 226584
rect 434640 225554 434668 226578
rect 434812 226296 434864 226302
rect 434812 226238 434864 226244
rect 434628 225548 434680 225554
rect 434628 225490 434680 225496
rect 434824 217410 434852 226238
rect 435640 223644 435692 223650
rect 435640 223586 435692 223592
rect 435652 217410 435680 223586
rect 436468 220448 436520 220454
rect 436468 220390 436520 220396
rect 436480 217410 436508 220390
rect 437308 217410 437336 229910
rect 440700 229900 440752 229906
rect 440700 229842 440752 229848
rect 438860 226976 438912 226982
rect 438860 226918 438912 226924
rect 438124 226160 438176 226166
rect 438124 226102 438176 226108
rect 438136 217410 438164 226102
rect 438872 225418 438900 226918
rect 438860 225412 438912 225418
rect 438860 225354 438912 225360
rect 439044 225344 439096 225350
rect 439044 225286 439096 225292
rect 439056 217410 439084 225286
rect 439780 220516 439832 220522
rect 439780 220458 439832 220464
rect 439792 217410 439820 220458
rect 440712 217410 440740 229842
rect 447416 229832 447468 229838
rect 447416 229774 447468 229780
rect 441620 226840 441672 226846
rect 441620 226782 441672 226788
rect 441632 225350 441660 226782
rect 444564 226772 444616 226778
rect 444564 226714 444616 226720
rect 441620 225344 441672 225350
rect 441620 225286 441672 225292
rect 444576 225282 444604 226714
rect 444564 225276 444616 225282
rect 444564 225218 444616 225224
rect 444840 225208 444892 225214
rect 444840 225150 444892 225156
rect 444104 225140 444156 225146
rect 444104 225082 444156 225088
rect 444116 224738 444144 225082
rect 442356 224732 442408 224738
rect 442356 224674 442408 224680
rect 444104 224732 444156 224738
rect 444104 224674 444156 224680
rect 441620 224392 441672 224398
rect 441620 224334 441672 224340
rect 441632 217410 441660 224334
rect 442368 217410 442396 224674
rect 444380 223916 444432 223922
rect 444380 223858 444432 223864
rect 443184 220312 443236 220318
rect 443184 220254 443236 220260
rect 443196 217410 443224 220254
rect 444392 217410 444420 223858
rect 425532 217382 425868 217410
rect 426360 217382 426696 217410
rect 427188 217382 427524 217410
rect 428016 217382 428352 217410
rect 428936 217382 429272 217410
rect 429764 217382 430100 217410
rect 430592 217382 430928 217410
rect 431420 217382 431756 217410
rect 432248 217382 432584 217410
rect 433352 217382 433412 217410
rect 433904 217382 434240 217410
rect 434824 217382 435160 217410
rect 435652 217382 435988 217410
rect 436480 217382 436816 217410
rect 437308 217382 437644 217410
rect 438136 217382 438472 217410
rect 439056 217382 439300 217410
rect 439792 217382 440128 217410
rect 440712 217382 441048 217410
rect 441632 217382 441876 217410
rect 442368 217382 442704 217410
rect 443196 217382 443532 217410
rect 444360 217382 444420 217410
rect 444852 217410 444880 225150
rect 445668 224120 445720 224126
rect 445668 224062 445720 224068
rect 445680 217410 445708 224062
rect 446588 220380 446640 220386
rect 446588 220322 446640 220328
rect 446600 217410 446628 220322
rect 447428 217410 447456 229774
rect 455788 229764 455840 229770
rect 455788 229706 455840 229712
rect 453672 227656 453724 227662
rect 453672 227598 453724 227604
rect 449624 226908 449676 226914
rect 449624 226850 449676 226856
rect 448244 226092 448296 226098
rect 448244 226034 448296 226040
rect 448256 217410 448284 226034
rect 449636 225214 449664 226850
rect 451188 226704 451240 226710
rect 451188 226646 451240 226652
rect 449624 225208 449676 225214
rect 449624 225150 449676 225156
rect 451200 225146 451228 226646
rect 453684 226030 453712 227598
rect 455420 227588 455472 227594
rect 455420 227530 455472 227536
rect 453672 226024 453724 226030
rect 453672 225966 453724 225972
rect 455432 225962 455460 227530
rect 452660 225956 452712 225962
rect 452660 225898 452712 225904
rect 454960 225956 455012 225962
rect 454960 225898 455012 225904
rect 455420 225956 455472 225962
rect 455420 225898 455472 225904
rect 449072 225140 449124 225146
rect 449072 225082 449124 225088
rect 451188 225140 451240 225146
rect 451188 225082 451240 225088
rect 449084 217410 449112 225082
rect 451556 224732 451608 224738
rect 451556 224674 451608 224680
rect 450728 224256 450780 224262
rect 450728 224198 450780 224204
rect 449900 220176 449952 220182
rect 449900 220118 449952 220124
rect 449912 217410 449940 220118
rect 450740 217410 450768 224198
rect 451568 217410 451596 224674
rect 452672 217410 452700 225898
rect 454132 221332 454184 221338
rect 454132 221274 454184 221280
rect 453304 220244 453356 220250
rect 453304 220186 453356 220192
rect 453316 217410 453344 220186
rect 454144 217410 454172 221274
rect 454972 217410 455000 225898
rect 455800 217410 455828 229706
rect 459192 229696 459244 229702
rect 459192 229638 459244 229644
rect 458456 225752 458508 225758
rect 458456 225694 458508 225700
rect 457444 224528 457496 224534
rect 457444 224470 457496 224476
rect 456616 220040 456668 220046
rect 456616 219982 456668 219988
rect 456628 217410 456656 219982
rect 457456 217410 457484 224470
rect 458468 217410 458496 225694
rect 459204 217410 459232 229638
rect 466000 229628 466052 229634
rect 466000 229570 466052 229576
rect 460940 229084 460992 229090
rect 460940 229026 460992 229032
rect 460952 225758 460980 229026
rect 465908 228676 465960 228682
rect 465908 228618 465960 228624
rect 465920 226098 465948 228618
rect 465908 226092 465960 226098
rect 465908 226034 465960 226040
rect 462504 225888 462556 225894
rect 462504 225830 462556 225836
rect 461676 225820 461728 225826
rect 461676 225762 461728 225768
rect 460940 225752 460992 225758
rect 460940 225694 460992 225700
rect 460940 221400 460992 221406
rect 460940 221342 460992 221348
rect 460020 220108 460072 220114
rect 460020 220050 460072 220056
rect 460032 217410 460060 220050
rect 460952 217410 460980 221342
rect 461688 217410 461716 225762
rect 462516 217410 462544 225830
rect 465080 225616 465132 225622
rect 465080 225558 465132 225564
rect 464252 224596 464304 224602
rect 464252 224538 464304 224544
rect 463700 219904 463752 219910
rect 463700 219846 463752 219852
rect 463712 217410 463740 219846
rect 444852 217382 445188 217410
rect 445680 217382 446016 217410
rect 446600 217382 446936 217410
rect 447428 217382 447764 217410
rect 448256 217382 448592 217410
rect 449084 217382 449420 217410
rect 449912 217382 450248 217410
rect 450740 217382 451076 217410
rect 451568 217382 451904 217410
rect 452672 217382 452824 217410
rect 453316 217382 453652 217410
rect 454144 217382 454480 217410
rect 454972 217382 455308 217410
rect 455800 217382 456136 217410
rect 456628 217382 456964 217410
rect 457456 217382 457792 217410
rect 458468 217382 458712 217410
rect 459204 217382 459540 217410
rect 460032 217382 460368 217410
rect 460952 217382 461196 217410
rect 461688 217382 462024 217410
rect 462516 217382 462852 217410
rect 463680 217382 463740 217410
rect 464264 217410 464292 224538
rect 465092 217410 465120 225558
rect 466012 217410 466040 229570
rect 474280 229560 474332 229566
rect 474280 229502 474332 229508
rect 473452 229492 473504 229498
rect 473452 229434 473504 229440
rect 472624 229424 472676 229430
rect 472624 229366 472676 229372
rect 469864 228948 469916 228954
rect 469864 228890 469916 228896
rect 469876 225894 469904 228890
rect 469864 225888 469916 225894
rect 469864 225830 469916 225836
rect 468392 225684 468444 225690
rect 468392 225626 468444 225632
rect 467564 221468 467616 221474
rect 467564 221410 467616 221416
rect 466736 219972 466788 219978
rect 466736 219914 466788 219920
rect 466748 217410 466776 219914
rect 467576 217410 467604 221410
rect 468404 217410 468432 225626
rect 470968 224800 471020 224806
rect 470968 224742 471020 224748
rect 469220 224188 469272 224194
rect 469220 224130 469272 224136
rect 469232 217410 469260 224130
rect 470140 219836 470192 219842
rect 470140 219778 470192 219784
rect 470152 217410 470180 219778
rect 470980 217410 471008 224742
rect 471978 224496 472034 224505
rect 471978 224431 472034 224440
rect 471992 217410 472020 224431
rect 472636 217410 472664 229366
rect 473268 228812 473320 228818
rect 473268 228754 473320 228760
rect 473280 225690 473308 228754
rect 473268 225684 473320 225690
rect 473268 225626 473320 225632
rect 473464 217410 473492 229434
rect 474292 217410 474320 229502
rect 479340 229356 479392 229362
rect 479340 229298 479392 229304
rect 477500 229016 477552 229022
rect 477500 228958 477552 228964
rect 474740 228880 474792 228886
rect 474740 228822 474792 228828
rect 474752 225826 474780 228822
rect 474740 225820 474792 225826
rect 474740 225762 474792 225768
rect 477512 225622 477540 228958
rect 478510 226264 478566 226273
rect 478510 226199 478566 226208
rect 477500 225616 477552 225622
rect 477500 225558 477552 225564
rect 476028 225480 476080 225486
rect 476028 225422 476080 225428
rect 475106 224632 475162 224641
rect 475106 224567 475162 224576
rect 475120 217410 475148 224567
rect 476040 217410 476068 225422
rect 477776 224868 477828 224874
rect 477776 224810 477828 224816
rect 476856 221264 476908 221270
rect 476856 221206 476908 221212
rect 476868 217410 476896 221206
rect 477788 217410 477816 224810
rect 478524 217410 478552 226199
rect 479352 217410 479380 229298
rect 487160 229288 487212 229294
rect 487160 229230 487212 229236
rect 480260 228744 480312 228750
rect 480260 228686 480312 228692
rect 480272 225486 480300 228686
rect 486054 227216 486110 227225
rect 486054 227151 486110 227160
rect 483020 226228 483072 226234
rect 483020 226170 483072 226176
rect 480260 225480 480312 225486
rect 480260 225422 480312 225428
rect 481914 224768 481970 224777
rect 481914 224703 481970 224712
rect 480258 224360 480314 224369
rect 480258 224295 480314 224304
rect 480272 217410 480300 224295
rect 480996 221536 481048 221542
rect 480996 221478 481048 221484
rect 481008 217410 481036 221478
rect 481928 217410 481956 224703
rect 483032 217410 483060 226170
rect 483570 222048 483626 222057
rect 483570 221983 483626 221992
rect 464264 217382 464600 217410
rect 465092 217382 465428 217410
rect 466012 217382 466256 217410
rect 466748 217382 467084 217410
rect 467576 217382 467912 217410
rect 468404 217382 468740 217410
rect 469232 217382 469568 217410
rect 470152 217382 470488 217410
rect 470980 217382 471316 217410
rect 471992 217382 472144 217410
rect 472636 217382 472972 217410
rect 473464 217382 473800 217410
rect 474292 217382 474628 217410
rect 475120 217382 475456 217410
rect 476040 217382 476376 217410
rect 476868 217382 477204 217410
rect 477788 217382 478032 217410
rect 478524 217382 478860 217410
rect 479352 217382 479688 217410
rect 480272 217382 480516 217410
rect 481008 217382 481344 217410
rect 481928 217382 482264 217410
rect 483032 217382 483092 217410
rect 418620 216708 418672 216714
rect 418620 216650 418672 216656
rect 59360 216640 59412 216646
rect 59360 216582 59412 216588
rect 417884 216640 417936 216646
rect 417884 216582 417936 216588
rect 483584 216458 483612 221983
rect 484400 221604 484452 221610
rect 484400 221546 484452 221552
rect 484412 217410 484440 221546
rect 485228 221196 485280 221202
rect 485228 221138 485280 221144
rect 485240 217410 485268 221138
rect 484412 217382 484748 217410
rect 485240 217382 485576 217410
rect 486068 216458 486096 227151
rect 487172 218142 487200 229230
rect 528376 229220 528428 229226
rect 528376 229162 528428 229168
rect 504546 228984 504602 228993
rect 504546 228919 504602 228928
rect 499670 228848 499726 228857
rect 499670 228783 499726 228792
rect 497832 228472 497884 228478
rect 497832 228414 497884 228420
rect 496818 227488 496874 227497
rect 496818 227423 496874 227432
rect 492310 227352 492366 227361
rect 492310 227287 492366 227296
rect 487804 226092 487856 226098
rect 487804 226034 487856 226040
rect 487160 218136 487212 218142
rect 487160 218078 487212 218084
rect 487172 217410 487200 218078
rect 487816 217410 487844 226034
rect 488630 223544 488686 223553
rect 488630 223479 488686 223488
rect 488644 221241 488672 223479
rect 489458 223408 489514 223417
rect 489458 223343 489514 223352
rect 488630 221232 488686 221241
rect 488630 221167 488686 221176
rect 488644 217410 488672 221167
rect 487172 217382 487232 217410
rect 487816 217382 488152 217410
rect 488644 217382 488980 217410
rect 489472 216458 489500 223343
rect 491390 221912 491446 221921
rect 491300 221876 491352 221882
rect 491390 221847 491446 221856
rect 491300 221818 491352 221824
rect 490288 221740 490340 221746
rect 490288 221682 490340 221688
rect 490300 218210 490328 221682
rect 490288 218204 490340 218210
rect 490288 218146 490340 218152
rect 490300 217410 490328 218146
rect 491312 217410 491340 221818
rect 491404 220969 491432 221847
rect 491390 220960 491446 220969
rect 491390 220895 491446 220904
rect 492324 217410 492352 227287
rect 495808 223508 495860 223514
rect 495808 223450 495860 223456
rect 495346 223272 495402 223281
rect 495346 223207 495402 223216
rect 494058 223136 494114 223145
rect 494058 223071 494114 223080
rect 494072 221105 494100 223071
rect 494520 221808 494572 221814
rect 494520 221750 494572 221756
rect 494152 221672 494204 221678
rect 494152 221614 494204 221620
rect 494058 221096 494114 221105
rect 494058 221031 494114 221040
rect 493046 220960 493102 220969
rect 493046 220895 493102 220904
rect 493060 217410 493088 220895
rect 494164 217410 494192 221614
rect 490300 217382 490636 217410
rect 491312 217382 491464 217410
rect 492292 217382 492536 217410
rect 493060 217382 493120 217410
rect 494040 217382 494192 217410
rect 494532 217410 494560 221750
rect 494532 217382 494868 217410
rect 492508 216578 492536 217382
rect 492496 216572 492548 216578
rect 492496 216514 492548 216520
rect 495360 216458 495388 223207
rect 495820 221678 495848 223450
rect 495808 221672 495860 221678
rect 495808 221614 495860 221620
rect 496832 221377 496860 227423
rect 497372 222012 497424 222018
rect 497372 221954 497424 221960
rect 496818 221368 496874 221377
rect 496818 221303 496874 221312
rect 496450 221096 496506 221105
rect 496450 221031 496506 221040
rect 496464 217410 496492 221031
rect 497384 217410 497412 221954
rect 496464 217382 496524 217410
rect 497352 217382 497412 217410
rect 497844 217410 497872 228414
rect 499028 222012 499080 222018
rect 499028 221954 499080 221960
rect 499040 220930 499068 221954
rect 499302 221368 499358 221377
rect 499302 221303 499358 221312
rect 499028 220924 499080 220930
rect 499028 220866 499080 220872
rect 499316 217410 499344 221303
rect 497844 217382 498180 217410
rect 499008 217382 499344 217410
rect 495992 216504 496044 216510
rect 483584 216442 484256 216458
rect 486068 216442 486740 216458
rect 489472 216442 490144 216458
rect 495360 216452 495992 216458
rect 495360 216446 496044 216452
rect 499684 216458 499712 228783
rect 503720 228404 503772 228410
rect 503720 228346 503772 228352
rect 500684 226024 500736 226030
rect 500684 225966 500736 225972
rect 500696 220998 500724 225966
rect 502706 222864 502762 222873
rect 502706 222799 502762 222808
rect 501236 221944 501288 221950
rect 501236 221886 501288 221892
rect 500684 220992 500736 220998
rect 500684 220934 500736 220940
rect 500696 217410 500724 220934
rect 501248 217410 501276 221886
rect 502720 221649 502748 222799
rect 503536 222148 503588 222154
rect 503536 222090 503588 222096
rect 502706 221640 502762 221649
rect 502706 221575 502762 221584
rect 502720 217410 502748 221575
rect 503548 221134 503576 222090
rect 503536 221128 503588 221134
rect 503536 221070 503588 221076
rect 503548 217410 503576 221070
rect 500696 217382 500756 217410
rect 501248 217382 501584 217410
rect 502412 217382 502748 217410
rect 503240 217382 503576 217410
rect 503732 217410 503760 228346
rect 503732 217382 504068 217410
rect 504560 216594 504588 228919
rect 509882 228712 509938 228721
rect 509882 228647 509938 228656
rect 508780 228336 508832 228342
rect 508780 228278 508832 228284
rect 505744 225956 505796 225962
rect 505744 225898 505796 225904
rect 505756 221202 505784 225898
rect 507122 223000 507178 223009
rect 507122 222935 507178 222944
rect 506296 222080 506348 222086
rect 506296 222022 506348 222028
rect 505744 221196 505796 221202
rect 505744 221138 505796 221144
rect 505756 217410 505784 221138
rect 506308 217410 506336 222022
rect 507136 221513 507164 222935
rect 507122 221504 507178 221513
rect 507122 221439 507178 221448
rect 507136 217410 507164 221439
rect 507952 221400 508004 221406
rect 507952 221342 508004 221348
rect 507964 220862 507992 221342
rect 507952 220856 508004 220862
rect 507952 220798 508004 220804
rect 507964 217410 507992 220798
rect 508792 217410 508820 228278
rect 509896 217410 509924 228647
rect 516232 228608 516284 228614
rect 514666 228576 514722 228585
rect 516232 228550 516284 228556
rect 514666 228511 514722 228520
rect 513840 228268 513892 228274
rect 513840 228210 513892 228216
rect 513470 226128 513526 226137
rect 513470 226063 513526 226072
rect 510712 225752 510764 225758
rect 510712 225694 510764 225700
rect 510618 222728 510674 222737
rect 510618 222663 510674 222672
rect 510632 221785 510660 222663
rect 510618 221776 510674 221785
rect 510618 221711 510674 221720
rect 510724 221338 510752 225694
rect 511356 223576 511408 223582
rect 511356 223518 511408 223524
rect 510712 221332 510764 221338
rect 510712 221274 510764 221280
rect 510724 217410 510752 221274
rect 511368 217410 511396 223518
rect 513380 223440 513432 223446
rect 513380 223382 513432 223388
rect 512458 221776 512514 221785
rect 512458 221711 512514 221720
rect 512472 217410 512500 221711
rect 513392 217410 513420 223382
rect 513484 218278 513512 226063
rect 513472 218272 513524 218278
rect 513472 218214 513524 218220
rect 513852 217410 513880 228210
rect 514680 217410 514708 228511
rect 516138 227080 516194 227089
rect 516138 227015 516194 227024
rect 516152 225758 516180 227015
rect 516244 225894 516272 228550
rect 518900 228540 518952 228546
rect 518900 228482 518952 228488
rect 517242 228440 517298 228449
rect 517242 228375 517298 228384
rect 516416 225956 516468 225962
rect 516416 225898 516468 225904
rect 516232 225888 516284 225894
rect 516232 225830 516284 225836
rect 516140 225752 516192 225758
rect 516140 225694 516192 225700
rect 515772 218272 515824 218278
rect 515772 218214 515824 218220
rect 515784 217410 515812 218214
rect 516428 217410 516456 225898
rect 517256 221066 517284 228375
rect 518714 225992 518770 226001
rect 518912 225962 518940 228482
rect 522486 228304 522542 228313
rect 522486 228239 522542 228248
rect 518714 225927 518770 225936
rect 518900 225956 518952 225962
rect 517244 221060 517296 221066
rect 517244 221002 517296 221008
rect 517888 221060 517940 221066
rect 517888 221002 517940 221008
rect 517900 217410 517928 221002
rect 518728 218346 518756 225927
rect 518900 225898 518952 225904
rect 520830 225720 520886 225729
rect 520830 225655 520886 225664
rect 521660 225684 521712 225690
rect 518900 223372 518952 223378
rect 518900 223314 518952 223320
rect 518716 218340 518768 218346
rect 518716 218282 518768 218288
rect 518728 217410 518756 218282
rect 505756 217382 505816 217410
rect 506308 217382 506644 217410
rect 507136 217382 507472 217410
rect 507964 217382 508300 217410
rect 508792 217382 509128 217410
rect 509896 217382 510292 217410
rect 510724 217382 510784 217410
rect 511368 217382 511704 217410
rect 512472 217382 512532 217410
rect 513360 217382 513512 217410
rect 513852 217382 514188 217410
rect 514680 217382 515260 217410
rect 515784 217382 515844 217410
rect 516428 217382 516672 217410
rect 517592 217382 517928 217410
rect 518420 217382 518756 217410
rect 518912 217410 518940 223314
rect 519726 222592 519782 222601
rect 519726 222527 519782 222536
rect 518912 217382 519248 217410
rect 504560 216578 505048 216594
rect 504456 216572 504508 216578
rect 504560 216572 505060 216578
rect 504560 216566 505008 216572
rect 504456 216514 504508 216520
rect 505008 216514 505060 216520
rect 483584 216436 484268 216442
rect 483584 216430 484216 216436
rect 486068 216436 486752 216442
rect 486068 216430 486700 216436
rect 484216 216378 484268 216384
rect 489472 216436 490156 216442
rect 489472 216430 490104 216436
rect 486700 216378 486752 216384
rect 495360 216430 496032 216446
rect 499684 216442 500264 216458
rect 504468 216442 504496 216514
rect 510264 216442 510292 217382
rect 513484 216986 513512 217382
rect 513472 216980 513524 216986
rect 513472 216922 513524 216928
rect 515232 216510 515260 217382
rect 519740 216594 519768 222527
rect 520844 218414 520872 225655
rect 521660 225626 521712 225632
rect 520832 218408 520884 218414
rect 520832 218350 520884 218356
rect 520844 217410 520872 218350
rect 521672 217410 521700 225626
rect 522500 221921 522528 228239
rect 527546 228168 527602 228177
rect 527546 228103 527602 228112
rect 526444 225820 526496 225826
rect 526444 225762 526496 225768
rect 525798 225584 525854 225593
rect 525798 225519 525854 225528
rect 523406 225448 523462 225457
rect 523406 225383 523462 225392
rect 522486 221912 522542 221921
rect 522486 221847 522542 221856
rect 522500 217410 522528 221847
rect 523420 218550 523448 225383
rect 523960 223304 524012 223310
rect 523960 223246 524012 223252
rect 523408 218544 523460 218550
rect 523408 218486 523460 218492
rect 523420 217410 523448 218486
rect 523972 217410 524000 223246
rect 525062 222456 525118 222465
rect 525062 222391 525118 222400
rect 525076 217410 525104 222391
rect 525812 218482 525840 225519
rect 525800 218476 525852 218482
rect 525800 218418 525852 218424
rect 525812 217410 525840 218418
rect 526456 217410 526484 225762
rect 527560 221270 527588 228103
rect 528388 221678 528416 229162
rect 535552 229152 535604 229158
rect 535552 229094 535604 229100
rect 535458 228032 535514 228041
rect 535458 227967 535514 227976
rect 532698 227896 532754 227905
rect 532698 227831 532754 227840
rect 530674 225856 530730 225865
rect 530674 225791 530730 225800
rect 529020 223236 529072 223242
rect 529020 223178 529072 223184
rect 528376 221672 528428 221678
rect 528376 221614 528428 221620
rect 527548 221264 527600 221270
rect 527548 221206 527600 221212
rect 527560 217410 527588 221206
rect 528388 217410 528416 221614
rect 529032 217410 529060 223178
rect 529938 222184 529994 222193
rect 529938 222119 529994 222128
rect 529952 217410 529980 222119
rect 530688 221814 530716 225791
rect 531504 225616 531556 225622
rect 531504 225558 531556 225564
rect 530676 221808 530728 221814
rect 530676 221750 530728 221756
rect 530688 217410 530716 221750
rect 531516 217410 531544 225558
rect 532712 221542 532740 227831
rect 532792 225548 532844 225554
rect 532792 225490 532844 225496
rect 532804 221950 532832 225490
rect 533988 223168 534040 223174
rect 533988 223110 534040 223116
rect 532792 221944 532844 221950
rect 532792 221886 532844 221892
rect 533436 221944 533488 221950
rect 533436 221886 533488 221892
rect 532700 221536 532752 221542
rect 532700 221478 532752 221484
rect 532976 221536 533028 221542
rect 532976 221478 533028 221484
rect 532988 217410 533016 221478
rect 520844 217382 520904 217410
rect 521672 217382 521732 217410
rect 522500 217382 522560 217410
rect 523420 217382 523480 217410
rect 523972 217382 524308 217410
rect 525076 217382 525472 217410
rect 525812 217382 525964 217410
rect 526456 217382 526792 217410
rect 527560 217382 527620 217410
rect 528388 217382 528448 217410
rect 529032 217382 529368 217410
rect 529952 217382 530348 217410
rect 530688 217382 531024 217410
rect 531516 217382 531852 217410
rect 532680 217382 533016 217410
rect 533448 217410 533476 221886
rect 534000 217410 534028 223110
rect 534906 222320 534962 222329
rect 534906 222255 534962 222264
rect 534920 217410 534948 222255
rect 535472 221474 535500 227967
rect 535564 223174 535592 229094
rect 541624 228200 541676 228206
rect 541624 228142 541676 228148
rect 536564 225480 536616 225486
rect 536564 225422 536616 225428
rect 535552 223168 535604 223174
rect 535552 223110 535604 223116
rect 536104 223168 536156 223174
rect 536104 223110 536156 223116
rect 535460 221468 535512 221474
rect 535460 221410 535512 221416
rect 536116 217410 536144 223110
rect 533448 217382 533508 217410
rect 534000 217382 534336 217410
rect 534920 217382 535408 217410
rect 536084 217382 536144 217410
rect 536576 217410 536604 225422
rect 541440 225412 541492 225418
rect 541440 225354 541492 225360
rect 538862 225312 538918 225321
rect 538862 225247 538918 225256
rect 538876 222154 538904 225247
rect 539876 223100 539928 223106
rect 539876 223042 539928 223048
rect 539048 223032 539100 223038
rect 539048 222974 539100 222980
rect 538864 222148 538916 222154
rect 538864 222090 538916 222096
rect 538036 221468 538088 221474
rect 538036 221410 538088 221416
rect 538048 217410 538076 221410
rect 538876 217410 538904 222090
rect 536576 217382 536912 217410
rect 537740 217382 538076 217410
rect 538568 217382 538904 217410
rect 539060 217410 539088 222974
rect 539060 217382 539396 217410
rect 525444 216918 525472 217382
rect 530320 217054 530348 217382
rect 535380 217122 535408 217382
rect 539888 217138 539916 223042
rect 541452 223038 541480 225354
rect 541440 223032 541492 223038
rect 541440 222974 541492 222980
rect 541452 217410 541480 222974
rect 541144 217382 541480 217410
rect 541636 217410 541664 228142
rect 544108 228132 544160 228138
rect 544108 228074 544160 228080
rect 543554 225176 543610 225185
rect 543554 225111 543610 225120
rect 543568 223378 543596 225111
rect 543556 223372 543608 223378
rect 543556 223314 543608 223320
rect 543096 222964 543148 222970
rect 543096 222906 543148 222912
rect 543108 221610 543136 222906
rect 543096 221604 543148 221610
rect 543096 221546 543148 221552
rect 543108 217410 543136 221546
rect 541636 217382 541972 217410
rect 542800 217382 543136 217410
rect 543568 217410 543596 223314
rect 544120 217410 544148 228074
rect 545212 228064 545264 228070
rect 545212 228006 545264 228012
rect 545224 221746 545252 228006
rect 549260 227996 549312 228002
rect 549260 227938 549312 227944
rect 545764 225344 545816 225350
rect 545764 225286 545816 225292
rect 545776 223242 545804 225286
rect 545764 223236 545816 223242
rect 545764 223178 545816 223184
rect 545212 221740 545264 221746
rect 545212 221682 545264 221688
rect 545224 217410 545252 221682
rect 545776 217410 545804 223178
rect 547512 222896 547564 222902
rect 547512 222838 547564 222844
rect 546684 222828 546736 222834
rect 546684 222770 546736 222776
rect 546696 217410 546724 222770
rect 547524 221882 547552 222838
rect 548340 222760 548392 222766
rect 548340 222702 548392 222708
rect 547512 221876 547564 221882
rect 547512 221818 547564 221824
rect 547524 217410 547552 221818
rect 548352 220862 548380 222702
rect 548340 220856 548392 220862
rect 548340 220798 548392 220804
rect 548352 217410 548380 220798
rect 549272 217410 549300 227938
rect 554228 227928 554280 227934
rect 554228 227870 554280 227876
rect 550270 227760 550326 227769
rect 550270 227695 550326 227704
rect 549350 225040 549406 225049
rect 549350 224975 549406 224984
rect 549364 222834 549392 224975
rect 549352 222828 549404 222834
rect 549352 222770 549404 222776
rect 550284 217410 550312 227695
rect 552018 224904 552074 224913
rect 552018 224839 552074 224848
rect 552032 223310 552060 224839
rect 552020 223304 552072 223310
rect 552020 223246 552072 223252
rect 553676 223304 553728 223310
rect 553676 223246 553728 223252
rect 551100 222828 551152 222834
rect 551100 222770 551152 222776
rect 551112 217410 551140 222770
rect 552020 222692 552072 222698
rect 552020 222634 552072 222640
rect 552032 217410 552060 222634
rect 552112 222556 552164 222562
rect 552112 222498 552164 222504
rect 552124 222018 552152 222498
rect 552112 222012 552164 222018
rect 552112 221954 552164 221960
rect 552848 222012 552900 222018
rect 552848 221954 552900 221960
rect 543568 217382 543628 217410
rect 544120 217382 544456 217410
rect 545224 217382 545284 217410
rect 545776 217382 546112 217410
rect 546696 217382 547032 217410
rect 547524 217382 547860 217410
rect 548352 217382 548688 217410
rect 549272 217382 549516 217410
rect 550284 217382 550680 217410
rect 551112 217382 551172 217410
rect 552000 217382 552060 217410
rect 552860 217410 552888 221954
rect 553688 217410 553716 223246
rect 554240 217410 554268 227870
rect 559288 227860 559340 227866
rect 559288 227802 559340 227808
rect 555054 227624 555110 227633
rect 555054 227559 555110 227568
rect 555068 222086 555096 227559
rect 557448 225276 557500 225282
rect 557448 225218 557500 225224
rect 557460 222630 557488 225218
rect 556712 222624 556764 222630
rect 556712 222566 556764 222572
rect 557448 222624 557500 222630
rect 557448 222566 557500 222572
rect 556528 222556 556580 222562
rect 556528 222498 556580 222504
rect 555056 222080 555108 222086
rect 555056 222022 555108 222028
rect 555068 217410 555096 222022
rect 556540 217410 556568 222498
rect 552860 217382 552920 217410
rect 553688 217382 553748 217410
rect 554240 217382 554576 217410
rect 555068 217382 555404 217410
rect 556232 217382 556568 217410
rect 556724 217410 556752 222566
rect 558828 222488 558880 222494
rect 558828 222430 558880 222436
rect 557540 222352 557592 222358
rect 557540 222294 557592 222300
rect 556724 217382 557060 217410
rect 550652 217258 550680 217382
rect 557552 217274 557580 222294
rect 558840 217410 558868 222430
rect 558808 217382 558868 217410
rect 559300 217410 559328 227802
rect 565452 227792 565504 227798
rect 565452 227734 565504 227740
rect 560392 225956 560444 225962
rect 560392 225898 560444 225904
rect 560208 223100 560260 223106
rect 560208 223042 560260 223048
rect 560220 222494 560248 223042
rect 560404 222494 560432 225898
rect 564348 225888 564400 225894
rect 564348 225830 564400 225836
rect 561220 225208 561272 225214
rect 561220 225150 561272 225156
rect 561232 222562 561260 225150
rect 563704 225072 563756 225078
rect 563704 225014 563756 225020
rect 561220 222556 561272 222562
rect 561220 222498 561272 222504
rect 560208 222488 560260 222494
rect 560208 222430 560260 222436
rect 560392 222488 560444 222494
rect 560392 222430 560444 222436
rect 560404 217410 560432 222430
rect 561232 217410 561260 222498
rect 563716 222494 563744 225014
rect 563704 222488 563756 222494
rect 563704 222430 563756 222436
rect 561772 222420 561824 222426
rect 561772 222362 561824 222368
rect 561784 217410 561812 222362
rect 562876 222284 562928 222290
rect 562876 222226 562928 222232
rect 562888 217410 562916 222226
rect 563716 217410 563744 222430
rect 564360 217410 564388 225830
rect 565464 222290 565492 227734
rect 567936 227724 567988 227730
rect 567936 227666 567988 227672
rect 566832 225752 566884 225758
rect 566832 225694 566884 225700
rect 566004 225140 566056 225146
rect 566004 225082 566056 225088
rect 566016 222902 566044 225082
rect 566004 222896 566056 222902
rect 566004 222838 566056 222844
rect 565452 222284 565504 222290
rect 565452 222226 565504 222232
rect 565464 217410 565492 222226
rect 566016 217410 566044 222838
rect 566844 217410 566872 225694
rect 567948 222766 567976 227666
rect 570236 225004 570288 225010
rect 570236 224946 570288 224952
rect 568580 224936 568632 224942
rect 568580 224878 568632 224884
rect 567936 222760 567988 222766
rect 567936 222702 567988 222708
rect 567948 217410 567976 222702
rect 568592 222698 568620 224878
rect 568580 222692 568632 222698
rect 568580 222634 568632 222640
rect 568592 217410 568620 222634
rect 569316 222216 569368 222222
rect 569316 222158 569368 222164
rect 569328 217410 569356 222158
rect 570248 217410 570276 224946
rect 570696 217456 570748 217462
rect 559300 217382 559636 217410
rect 560404 217382 560464 217410
rect 561232 217382 561292 217410
rect 561784 217382 562120 217410
rect 562888 217394 563100 217410
rect 562888 217388 563112 217394
rect 562888 217382 563060 217388
rect 563716 217382 563776 217410
rect 564360 217382 564696 217410
rect 565464 217382 565524 217410
rect 566016 217382 566352 217410
rect 566844 217382 567180 217410
rect 567948 217382 568008 217410
rect 568592 217382 568836 217410
rect 569328 217382 569664 217410
rect 570248 217404 570696 217410
rect 571536 217410 571564 253914
rect 571616 245676 571668 245682
rect 571616 245618 571668 245624
rect 571628 220726 571656 245618
rect 571720 220794 571748 262210
rect 571800 256760 571852 256766
rect 571800 256702 571852 256708
rect 571708 220788 571760 220794
rect 571708 220730 571760 220736
rect 571616 220720 571668 220726
rect 571616 220662 571668 220668
rect 570248 217398 570748 217404
rect 570248 217382 570736 217398
rect 571412 217382 571564 217410
rect 571812 217410 571840 256702
rect 574100 251252 574152 251258
rect 574100 251194 574152 251200
rect 574112 220794 574140 251194
rect 574192 248464 574244 248470
rect 574192 248406 574244 248412
rect 574204 226334 574232 248406
rect 574204 226306 574324 226334
rect 572720 220788 572772 220794
rect 572720 220730 572772 220736
rect 574100 220788 574152 220794
rect 574100 220730 574152 220736
rect 572732 217410 572760 220730
rect 573548 220720 573600 220726
rect 573548 220662 573600 220668
rect 573560 217410 573588 220662
rect 574296 217410 574324 226306
rect 607588 223508 607640 223514
rect 607588 223450 607640 223456
rect 575204 220788 575256 220794
rect 575204 220730 575256 220736
rect 575216 217410 575244 220730
rect 607128 218204 607180 218210
rect 607128 218146 607180 218152
rect 606668 218136 606720 218142
rect 606668 218078 606720 218084
rect 571812 217382 572240 217410
rect 572732 217382 573068 217410
rect 573560 217382 573896 217410
rect 574296 217382 574724 217410
rect 575216 217382 575552 217410
rect 563060 217330 563112 217336
rect 558184 217320 558236 217326
rect 557552 217268 558184 217274
rect 557552 217262 558236 217268
rect 550640 217252 550692 217258
rect 557552 217246 558224 217262
rect 550640 217194 550692 217200
rect 540520 217184 540572 217190
rect 539888 217132 540520 217138
rect 539888 217126 540572 217132
rect 535368 217116 535420 217122
rect 539888 217110 540560 217126
rect 535368 217058 535420 217064
rect 530308 217048 530360 217054
rect 530308 216990 530360 216996
rect 525432 216912 525484 216918
rect 525432 216854 525484 216860
rect 519740 216578 520412 216594
rect 519740 216572 520424 216578
rect 519740 216566 520372 216572
rect 520372 216514 520424 216520
rect 515220 216504 515272 216510
rect 515220 216446 515272 216452
rect 499684 216436 500276 216442
rect 499684 216430 500224 216436
rect 490104 216378 490156 216384
rect 500224 216378 500276 216384
rect 504456 216436 504508 216442
rect 504456 216378 504508 216384
rect 510252 216436 510304 216442
rect 510252 216378 510304 216384
rect 580170 216200 580226 216209
rect 580170 216135 580226 216144
rect 580184 215626 580212 216135
rect 580172 215620 580224 215626
rect 580172 215562 580224 215568
rect 599768 215620 599820 215626
rect 599768 215562 599820 215568
rect 582286 214704 582342 214713
rect 582286 214639 582342 214648
rect 580262 213208 580318 213217
rect 580262 213143 580318 213152
rect 580276 212566 580304 213143
rect 582300 212634 582328 214639
rect 582288 212628 582340 212634
rect 582288 212570 582340 212576
rect 580264 212560 580316 212566
rect 580264 212502 580316 212508
rect 581642 211712 581698 211721
rect 581642 211647 581698 211656
rect 580538 210216 580594 210225
rect 580538 210151 580594 210160
rect 580552 209846 580580 210151
rect 581656 209914 581684 211647
rect 581644 209908 581696 209914
rect 581644 209850 581696 209856
rect 580540 209840 580592 209846
rect 580540 209782 580592 209788
rect 599124 209840 599176 209846
rect 599124 209782 599176 209788
rect 579710 208720 579766 208729
rect 579710 208655 579766 208664
rect 579724 207126 579752 208655
rect 579712 207120 579764 207126
rect 579712 207062 579764 207068
rect 582286 207088 582342 207097
rect 582286 207023 582288 207032
rect 582340 207023 582342 207032
rect 582288 206994 582340 207000
rect 582286 205592 582342 205601
rect 582286 205527 582342 205536
rect 582300 204338 582328 205527
rect 599136 205465 599164 209782
rect 599780 209545 599808 215562
rect 599952 212628 600004 212634
rect 599952 212570 600004 212576
rect 599860 212560 599912 212566
rect 599860 212502 599912 212508
rect 599766 209536 599822 209545
rect 599766 209471 599822 209480
rect 599872 207505 599900 212502
rect 599964 208593 599992 212570
rect 606680 210202 606708 218078
rect 607140 210202 607168 218146
rect 607600 210202 607628 223450
rect 616420 223372 616472 223378
rect 616420 223314 616472 223320
rect 615040 223168 615092 223174
rect 615040 223110 615092 223116
rect 614580 221944 614632 221950
rect 614580 221886 614632 221892
rect 614028 221808 614080 221814
rect 614028 221750 614080 221756
rect 613568 221672 613620 221678
rect 613568 221614 613620 221620
rect 609888 221400 609940 221406
rect 609888 221342 609940 221348
rect 609428 221196 609480 221202
rect 609428 221138 609480 221144
rect 608968 221128 609020 221134
rect 608968 221070 609020 221076
rect 608508 220992 608560 220998
rect 608508 220934 608560 220940
rect 608048 220924 608100 220930
rect 608048 220866 608100 220872
rect 608060 210202 608088 220866
rect 608520 210202 608548 220934
rect 608980 210202 609008 221070
rect 609440 210202 609468 221138
rect 609900 210202 609928 221342
rect 610348 221332 610400 221338
rect 610348 221274 610400 221280
rect 610360 210202 610388 221274
rect 612648 218544 612700 218550
rect 612648 218486 612700 218492
rect 612188 218408 612240 218414
rect 612188 218350 612240 218356
rect 611728 218340 611780 218346
rect 611728 218282 611780 218288
rect 611268 218272 611320 218278
rect 611268 218214 611320 218220
rect 610808 216980 610860 216986
rect 610808 216922 610860 216928
rect 610820 210202 610848 216922
rect 611280 210202 611308 218214
rect 611740 210202 611768 218282
rect 612200 210202 612228 218350
rect 612660 210202 612688 218486
rect 613108 218476 613160 218482
rect 613108 218418 613160 218424
rect 613120 210202 613148 218418
rect 613580 210202 613608 221614
rect 614040 210202 614068 221750
rect 614592 210202 614620 221886
rect 615052 210202 615080 223110
rect 615960 223032 616012 223038
rect 615960 222974 616012 222980
rect 615500 222148 615552 222154
rect 615500 222090 615552 222096
rect 615512 210202 615540 222090
rect 615972 210202 616000 222974
rect 616432 210202 616460 223314
rect 618260 223304 618312 223310
rect 618260 223246 618312 223252
rect 616880 223236 616932 223242
rect 616880 223178 616932 223184
rect 616892 210202 616920 223178
rect 617800 222828 617852 222834
rect 617800 222770 617852 222776
rect 617340 220856 617392 220862
rect 617340 220798 617392 220804
rect 617352 210202 617380 220798
rect 617812 210202 617840 222770
rect 618272 210202 618300 223246
rect 619180 223100 619232 223106
rect 619180 223042 619232 223048
rect 618720 222624 618772 222630
rect 618720 222566 618772 222572
rect 618732 210202 618760 222566
rect 619192 210202 619220 223042
rect 620560 222896 620612 222902
rect 620560 222838 620612 222844
rect 620100 222488 620152 222494
rect 620100 222430 620152 222436
rect 619640 222420 619692 222426
rect 619640 222362 619692 222368
rect 619652 210202 619680 222362
rect 620112 210202 620140 222430
rect 620572 210202 620600 222838
rect 635464 222760 635516 222766
rect 635464 222702 635516 222708
rect 621020 222692 621072 222698
rect 621020 222634 621072 222640
rect 621032 210202 621060 222634
rect 634084 222352 634136 222358
rect 634084 222294 634136 222300
rect 633164 222080 633216 222086
rect 633164 222022 633216 222028
rect 632704 222012 632756 222018
rect 632704 221954 632756 221960
rect 627090 221912 627146 221921
rect 627090 221847 627146 221856
rect 631784 221876 631836 221882
rect 625250 221776 625306 221785
rect 625250 221711 625306 221720
rect 623410 221640 623466 221649
rect 623410 221575 623466 221584
rect 622950 221368 623006 221377
rect 622950 221303 623006 221312
rect 621478 221232 621534 221241
rect 621478 221167 621534 221176
rect 621492 210202 621520 221167
rect 622492 216300 622544 216306
rect 622492 216242 622544 216248
rect 622032 216232 622084 216238
rect 622032 216174 622084 216180
rect 622044 210202 622072 216174
rect 622504 210202 622532 216242
rect 622964 210202 622992 221303
rect 623424 210202 623452 221575
rect 624330 221504 624386 221513
rect 624330 221439 624386 221448
rect 623872 216368 623924 216374
rect 623872 216310 623924 216316
rect 623884 210202 623912 216310
rect 624344 210202 624372 221439
rect 624792 216436 624844 216442
rect 624792 216378 624844 216384
rect 624804 210202 624832 216378
rect 625264 210202 625292 221711
rect 626172 221060 626224 221066
rect 626172 221002 626224 221008
rect 625712 216504 625764 216510
rect 625712 216446 625764 216452
rect 625724 210202 625752 216446
rect 626184 210202 626212 221002
rect 626632 216572 626684 216578
rect 626632 216514 626684 216520
rect 626644 210202 626672 216514
rect 627104 210202 627132 221847
rect 631784 221818 631836 221824
rect 631324 221740 631376 221746
rect 631324 221682 631376 221688
rect 630864 221604 630916 221610
rect 630864 221546 630916 221552
rect 628932 221536 628984 221542
rect 628932 221478 628984 221484
rect 628012 221264 628064 221270
rect 628012 221206 628064 221212
rect 627552 216912 627604 216918
rect 627552 216854 627604 216860
rect 627564 210202 627592 216854
rect 628024 210202 628052 221206
rect 628472 217048 628524 217054
rect 628472 216990 628524 216996
rect 628484 210202 628512 216990
rect 628944 210202 628972 221478
rect 629944 221468 629996 221474
rect 629944 221410 629996 221416
rect 629484 217116 629536 217122
rect 629484 217058 629536 217064
rect 629496 210202 629524 217058
rect 629956 210202 629984 221410
rect 630404 217184 630456 217190
rect 630404 217126 630456 217132
rect 630416 210202 630444 217126
rect 630876 210202 630904 221546
rect 631336 210202 631364 221682
rect 631796 210202 631824 221818
rect 632244 217252 632296 217258
rect 632244 217194 632296 217200
rect 632256 210202 632284 217194
rect 632716 210202 632744 221954
rect 633176 210202 633204 222022
rect 633624 217320 633676 217326
rect 633624 217262 633676 217268
rect 633636 210202 633664 217262
rect 634096 210202 634124 222294
rect 635004 222284 635056 222290
rect 635004 222226 635056 222232
rect 634544 217388 634596 217394
rect 634544 217330 634596 217336
rect 634556 210202 634584 217330
rect 635016 210202 635044 222226
rect 635476 210202 635504 222702
rect 637394 221096 637450 221105
rect 637394 221031 637450 221040
rect 636934 220960 636990 220969
rect 636934 220895 636990 220904
rect 635924 217456 635976 217462
rect 635924 217398 635976 217404
rect 635936 210202 635964 217398
rect 636384 216096 636436 216102
rect 636384 216038 636436 216044
rect 636396 210202 636424 216038
rect 636948 210202 636976 220895
rect 637408 210202 637436 221031
rect 648528 219768 648580 219774
rect 648528 219710 648580 219716
rect 647148 219700 647200 219706
rect 647148 219642 647200 219648
rect 646964 218000 647016 218006
rect 646964 217942 647016 217948
rect 642732 217932 642784 217938
rect 642732 217874 642784 217880
rect 639696 216844 639748 216850
rect 639696 216786 639748 216792
rect 637856 216164 637908 216170
rect 637856 216106 637908 216112
rect 637868 210202 637896 216106
rect 638316 216028 638368 216034
rect 638316 215970 638368 215976
rect 638328 210202 638356 215970
rect 638776 215960 638828 215966
rect 638776 215902 638828 215908
rect 638788 210202 638816 215902
rect 639708 210202 639736 216786
rect 640616 216776 640668 216782
rect 640616 216718 640668 216724
rect 640156 216708 640208 216714
rect 640156 216650 640208 216656
rect 640168 210202 640196 216650
rect 640628 210202 640656 216718
rect 641076 216640 641128 216646
rect 641076 216582 641128 216588
rect 641088 210202 641116 216582
rect 641824 210310 642128 210338
rect 641824 210202 641852 210310
rect 606648 210174 606708 210202
rect 607108 210174 607168 210202
rect 607568 210174 607628 210202
rect 608028 210174 608088 210202
rect 608488 210174 608548 210202
rect 608948 210174 609008 210202
rect 609408 210174 609468 210202
rect 609868 210174 609928 210202
rect 610328 210174 610388 210202
rect 610788 210174 610848 210202
rect 611248 210174 611308 210202
rect 611708 210174 611768 210202
rect 612168 210174 612228 210202
rect 612628 210174 612688 210202
rect 613088 210174 613148 210202
rect 613548 210174 613608 210202
rect 614008 210174 614068 210202
rect 614560 210174 614620 210202
rect 615020 210174 615080 210202
rect 615480 210174 615540 210202
rect 615940 210174 616000 210202
rect 616400 210174 616460 210202
rect 616860 210174 616920 210202
rect 617320 210174 617380 210202
rect 617780 210174 617840 210202
rect 618240 210174 618300 210202
rect 618700 210174 618760 210202
rect 619160 210174 619220 210202
rect 619620 210174 619680 210202
rect 620080 210174 620140 210202
rect 620540 210174 620600 210202
rect 621000 210174 621060 210202
rect 621460 210174 621520 210202
rect 622012 210174 622072 210202
rect 622472 210174 622532 210202
rect 622932 210174 622992 210202
rect 623392 210174 623452 210202
rect 623852 210174 623912 210202
rect 624312 210174 624372 210202
rect 624772 210174 624832 210202
rect 625232 210174 625292 210202
rect 625692 210174 625752 210202
rect 626152 210174 626212 210202
rect 626612 210174 626672 210202
rect 627072 210174 627132 210202
rect 627532 210174 627592 210202
rect 627992 210174 628052 210202
rect 628452 210174 628512 210202
rect 628912 210174 628972 210202
rect 629464 210174 629524 210202
rect 629924 210174 629984 210202
rect 630384 210174 630444 210202
rect 630844 210174 630904 210202
rect 631304 210174 631364 210202
rect 631764 210174 631824 210202
rect 632224 210174 632284 210202
rect 632684 210174 632744 210202
rect 633144 210174 633204 210202
rect 633604 210174 633664 210202
rect 634064 210174 634124 210202
rect 634524 210174 634584 210202
rect 634984 210174 635044 210202
rect 635444 210174 635504 210202
rect 635904 210174 635964 210202
rect 636364 210174 636424 210202
rect 636916 210174 636976 210202
rect 637376 210174 637436 210202
rect 637836 210174 637896 210202
rect 638296 210174 638356 210202
rect 638756 210174 638816 210202
rect 639676 210174 639736 210202
rect 640136 210174 640196 210202
rect 640596 210174 640656 210202
rect 641056 210174 641116 210202
rect 641516 210174 641852 210202
rect 642100 210066 642128 210310
rect 642744 210202 642772 217874
rect 644112 217864 644164 217870
rect 644112 217806 644164 217812
rect 643204 210310 643508 210338
rect 643204 210202 643232 210310
rect 642436 210188 642772 210202
rect 642422 210174 642772 210188
rect 642896 210174 643232 210202
rect 642422 210066 642450 210174
rect 642100 210052 642450 210066
rect 643480 210066 643508 210310
rect 644124 210202 644152 217806
rect 645584 216708 645636 216714
rect 645584 216650 645636 216656
rect 644676 210310 644980 210338
rect 644676 210202 644704 210310
rect 643816 210188 644152 210202
rect 643802 210174 644152 210188
rect 644368 210174 644704 210202
rect 643802 210066 643830 210174
rect 643480 210052 643830 210066
rect 644952 210066 644980 210310
rect 645596 210202 645624 216650
rect 646056 210310 646360 210338
rect 646056 210202 646084 210310
rect 645288 210188 645624 210202
rect 645274 210174 645624 210188
rect 645748 210174 646084 210202
rect 645274 210066 645302 210174
rect 644952 210052 645302 210066
rect 646332 210066 646360 210310
rect 646976 210202 647004 217942
rect 647160 210202 647188 219642
rect 647436 210310 647740 210338
rect 647436 210202 647464 210310
rect 646668 210188 647004 210202
rect 646654 210174 647004 210188
rect 647128 210174 647464 210202
rect 646654 210066 646682 210174
rect 646332 210052 646682 210066
rect 647712 210066 647740 210310
rect 648540 210202 648568 219710
rect 651288 219632 651340 219638
rect 651288 219574 651340 219580
rect 649908 219564 649960 219570
rect 649908 219506 649960 219512
rect 648816 210310 649120 210338
rect 648816 210202 648844 210310
rect 648508 210174 648844 210202
rect 649092 210066 649120 210310
rect 649920 210202 649948 219506
rect 651300 212498 651328 219574
rect 651392 217938 651420 987566
rect 652852 987556 652904 987562
rect 652852 987498 652904 987504
rect 652668 987488 652720 987494
rect 652668 987430 652720 987436
rect 651472 987284 651524 987290
rect 651472 987226 651524 987232
rect 651380 217932 651432 217938
rect 651380 217874 651432 217880
rect 651484 217870 651512 987226
rect 651564 987012 651616 987018
rect 651564 986954 651616 986960
rect 651472 217864 651524 217870
rect 651472 217806 651524 217812
rect 651576 216714 651604 986954
rect 651656 986944 651708 986950
rect 651656 986886 651708 986892
rect 651668 218006 651696 986886
rect 652680 219366 652708 987430
rect 652760 987352 652812 987358
rect 652760 987294 652812 987300
rect 652772 219638 652800 987294
rect 652864 222222 652892 987498
rect 652944 987216 652996 987222
rect 652944 987158 652996 987164
rect 652956 266354 652984 987158
rect 658280 987148 658332 987154
rect 658280 987090 658332 987096
rect 658188 987080 658240 987086
rect 658188 987022 658240 987028
rect 655428 984292 655480 984298
rect 655428 984234 655480 984240
rect 654874 922720 654930 922729
rect 654874 922655 654930 922664
rect 654888 922282 654916 922655
rect 654876 922276 654928 922282
rect 654876 922218 654928 922224
rect 654874 909528 654930 909537
rect 654874 909463 654930 909472
rect 654888 908138 654916 909463
rect 654876 908132 654928 908138
rect 654876 908074 654928 908080
rect 654874 896200 654930 896209
rect 654874 896135 654930 896144
rect 654888 895558 654916 896135
rect 654876 895552 654928 895558
rect 654876 895494 654928 895500
rect 655150 882872 655206 882881
rect 655150 882807 655206 882816
rect 655164 870806 655192 882807
rect 655152 870800 655204 870806
rect 655152 870742 655204 870748
rect 654690 856352 654746 856361
rect 654690 856287 654746 856296
rect 654704 855710 654732 856287
rect 654692 855704 654744 855710
rect 654692 855646 654744 855652
rect 655058 843024 655114 843033
rect 655058 842959 655114 842968
rect 655072 841974 655100 842959
rect 655060 841968 655112 841974
rect 655060 841910 655112 841916
rect 654138 816504 654194 816513
rect 654138 816439 654194 816448
rect 654152 814774 654180 816439
rect 654140 814768 654192 814774
rect 654140 814710 654192 814716
rect 655058 789984 655114 789993
rect 655058 789919 655114 789928
rect 655072 789410 655100 789919
rect 655060 789404 655112 789410
rect 655060 789346 655112 789352
rect 654782 763328 654838 763337
rect 654782 763263 654838 763272
rect 654796 762822 654824 763263
rect 654784 762816 654836 762822
rect 654784 762758 654836 762764
rect 654874 750136 654930 750145
rect 654874 750071 654930 750080
rect 654888 749018 654916 750071
rect 654876 749012 654928 749018
rect 654876 748954 654928 748960
rect 654782 736808 654838 736817
rect 654782 736743 654838 736752
rect 654796 736030 654824 736743
rect 654784 736024 654836 736030
rect 654784 735966 654836 735972
rect 654690 696960 654746 696969
rect 654690 696895 654746 696904
rect 654704 695570 654732 696895
rect 654692 695564 654744 695570
rect 654692 695506 654744 695512
rect 654874 683632 654930 683641
rect 654874 683567 654930 683576
rect 654888 682990 654916 683567
rect 654876 682984 654928 682990
rect 654876 682926 654928 682932
rect 654874 643784 654930 643793
rect 654874 643719 654930 643728
rect 654888 643142 654916 643719
rect 654876 643136 654928 643142
rect 654876 643078 654928 643084
rect 655058 630592 655114 630601
rect 655058 630527 655114 630536
rect 655072 629338 655100 630527
rect 655060 629332 655112 629338
rect 655060 629274 655112 629280
rect 654598 617264 654654 617273
rect 654598 617199 654654 617208
rect 654322 603936 654378 603945
rect 654322 603871 654378 603880
rect 654336 602206 654364 603871
rect 654612 603090 654640 617199
rect 654600 603084 654652 603090
rect 654600 603026 654652 603032
rect 654324 602200 654376 602206
rect 654324 602142 654376 602148
rect 655058 577416 655114 577425
rect 655058 577351 655114 577360
rect 655072 576910 655100 577351
rect 655060 576904 655112 576910
rect 655060 576846 655112 576852
rect 654322 564088 654378 564097
rect 654322 564023 654378 564032
rect 654336 556170 654364 564023
rect 654324 556164 654376 556170
rect 654324 556106 654376 556112
rect 654690 550896 654746 550905
rect 654690 550831 654746 550840
rect 654704 549302 654732 550831
rect 654692 549296 654744 549302
rect 654692 549238 654744 549244
rect 654874 537568 654930 537577
rect 654874 537503 654930 537512
rect 654888 536450 654916 537503
rect 654876 536444 654928 536450
rect 654876 536386 654928 536392
rect 654138 524240 654194 524249
rect 654138 524175 654194 524184
rect 654152 522510 654180 524175
rect 654140 522504 654192 522510
rect 654140 522446 654192 522452
rect 654874 511048 654930 511057
rect 654874 510983 654930 510992
rect 654888 510882 654916 510983
rect 654876 510876 654928 510882
rect 654876 510818 654928 510824
rect 654874 484392 654930 484401
rect 654874 484327 654930 484336
rect 654888 483070 654916 484327
rect 654876 483064 654928 483070
rect 654876 483006 654928 483012
rect 654874 471200 654930 471209
rect 654874 471135 654930 471144
rect 654888 470830 654916 471135
rect 654876 470824 654928 470830
rect 654876 470766 654928 470772
rect 654230 457872 654286 457881
rect 654230 457807 654286 457816
rect 654244 457502 654272 457807
rect 654232 457496 654284 457502
rect 654232 457438 654284 457444
rect 654414 444544 654470 444553
rect 654414 444479 654416 444488
rect 654468 444479 654470 444488
rect 654416 444450 654468 444456
rect 654690 431352 654746 431361
rect 654690 431287 654746 431296
rect 654704 430642 654732 431287
rect 654692 430636 654744 430642
rect 654692 430578 654744 430584
rect 655058 418024 655114 418033
rect 655058 417959 655114 417968
rect 655072 416838 655100 417959
rect 655060 416832 655112 416838
rect 655060 416774 655112 416780
rect 654874 404696 654930 404705
rect 654874 404631 654930 404640
rect 654888 404054 654916 404631
rect 654876 404048 654928 404054
rect 654876 403990 654928 403996
rect 654322 391504 654378 391513
rect 654322 391439 654378 391448
rect 654336 389910 654364 391439
rect 654324 389904 654376 389910
rect 654324 389846 654376 389852
rect 654874 351656 654930 351665
rect 654874 351591 654930 351600
rect 654888 350606 654916 351591
rect 654876 350600 654928 350606
rect 654876 350542 654928 350548
rect 655058 338328 655114 338337
rect 655058 338263 655114 338272
rect 655072 336802 655100 338263
rect 655060 336796 655112 336802
rect 655060 336738 655112 336744
rect 654874 325000 654930 325009
rect 654874 324935 654930 324944
rect 654888 323950 654916 324935
rect 654876 323944 654928 323950
rect 654876 323886 654928 323892
rect 654138 311808 654194 311817
rect 654138 311743 654194 311752
rect 654152 311302 654180 311743
rect 654140 311296 654192 311302
rect 654140 311238 654192 311244
rect 655440 310486 655468 984234
rect 655518 975896 655574 975905
rect 655518 975831 655574 975840
rect 655532 938602 655560 975831
rect 655702 962568 655758 962577
rect 655702 962503 655758 962512
rect 655612 960560 655664 960566
rect 655612 960502 655664 960508
rect 655520 938596 655572 938602
rect 655520 938538 655572 938544
rect 655624 936193 655652 960502
rect 655716 938738 655744 962503
rect 655794 949376 655850 949385
rect 655794 949311 655850 949320
rect 655808 938874 655836 949311
rect 655796 938868 655848 938874
rect 655796 938810 655848 938816
rect 655704 938732 655756 938738
rect 655704 938674 655756 938680
rect 655610 936184 655666 936193
rect 655610 936119 655666 936128
rect 656806 869680 656862 869689
rect 656806 869615 656808 869624
rect 656860 869615 656862 869624
rect 656808 869586 656860 869592
rect 655518 829832 655574 829841
rect 655518 829767 655574 829776
rect 655532 782474 655560 829767
rect 656806 803312 656862 803321
rect 656806 803247 656808 803256
rect 656860 803247 656862 803256
rect 656808 803218 656860 803224
rect 655520 782468 655572 782474
rect 655520 782410 655572 782416
rect 655518 776656 655574 776665
rect 655518 776591 655574 776600
rect 655532 738342 655560 776591
rect 655520 738336 655572 738342
rect 655520 738278 655572 738284
rect 655518 723480 655574 723489
rect 655518 723415 655574 723424
rect 655532 691422 655560 723415
rect 655978 710288 656034 710297
rect 655978 710223 656034 710232
rect 655992 709782 656020 710223
rect 655980 709776 656032 709782
rect 655980 709718 656032 709724
rect 655520 691416 655572 691422
rect 655520 691358 655572 691364
rect 655518 670440 655574 670449
rect 655518 670375 655574 670384
rect 655532 647222 655560 670375
rect 656162 657112 656218 657121
rect 656162 657047 656164 657056
rect 656216 657047 656218 657056
rect 656164 657018 656216 657024
rect 655520 647216 655572 647222
rect 655520 647158 655572 647164
rect 656806 590744 656862 590753
rect 656806 590679 656808 590688
rect 656860 590679 656862 590688
rect 656808 590650 656860 590656
rect 656806 497720 656862 497729
rect 656806 497655 656808 497664
rect 656860 497655 656862 497664
rect 656808 497626 656860 497632
rect 656808 378208 656860 378214
rect 656806 378176 656808 378185
rect 656860 378176 656862 378185
rect 656806 378111 656862 378120
rect 656806 364848 656862 364857
rect 656806 364783 656862 364792
rect 656820 364478 656848 364783
rect 656808 364472 656860 364478
rect 656808 364414 656860 364420
rect 655428 310480 655480 310486
rect 655428 310422 655480 310428
rect 655610 298480 655666 298489
rect 655610 298415 655666 298424
rect 655624 298314 655652 298415
rect 655612 298308 655664 298314
rect 655612 298250 655664 298256
rect 655334 285288 655390 285297
rect 655334 285223 655390 285232
rect 655348 284782 655376 285223
rect 655336 284776 655388 284782
rect 655336 284718 655388 284724
rect 652944 266348 652996 266354
rect 652944 266290 652996 266296
rect 658200 262449 658228 987022
rect 658292 265062 658320 987090
rect 658464 984224 658516 984230
rect 658464 984166 658516 984172
rect 658372 984156 658424 984162
rect 658372 984098 658424 984104
rect 658384 311846 658412 984098
rect 658476 314634 658504 984166
rect 663800 908132 663852 908138
rect 663800 908074 663852 908080
rect 661132 895552 661184 895558
rect 661132 895494 661184 895500
rect 661040 855704 661092 855710
rect 661040 855646 661092 855652
rect 660948 814768 661000 814774
rect 660948 814710 661000 814716
rect 660960 670818 660988 814710
rect 661052 715018 661080 855646
rect 661144 759354 661172 895494
rect 663708 869644 663760 869650
rect 663708 869586 663760 869592
rect 661132 759348 661184 759354
rect 661132 759290 661184 759296
rect 661132 736024 661184 736030
rect 661132 735966 661184 735972
rect 661040 715012 661092 715018
rect 661040 714954 661092 714960
rect 660948 670812 661000 670818
rect 660948 670754 661000 670760
rect 660948 657076 661000 657082
rect 660948 657018 661000 657024
rect 660960 535634 660988 657018
rect 661144 623898 661172 735966
rect 663720 716174 663748 869586
rect 663812 759490 663840 908074
rect 666468 803276 666520 803282
rect 666468 803218 666520 803224
rect 663892 789404 663944 789410
rect 663892 789346 663944 789352
rect 663800 759484 663852 759490
rect 663800 759426 663852 759432
rect 663708 716168 663760 716174
rect 663708 716110 663760 716116
rect 663708 695564 663760 695570
rect 663708 695506 663760 695512
rect 661132 623892 661184 623898
rect 661132 623834 661184 623840
rect 661040 602200 661092 602206
rect 661040 602142 661092 602148
rect 660948 535628 661000 535634
rect 660948 535570 661000 535576
rect 661052 491434 661080 602142
rect 663720 579834 663748 695506
rect 663800 682984 663852 682990
rect 663800 682926 663852 682932
rect 663812 579970 663840 682926
rect 663904 670614 663932 789346
rect 666480 671566 666508 803218
rect 666468 671560 666520 671566
rect 666468 671502 666520 671508
rect 663892 670608 663944 670614
rect 663892 670550 663944 670556
rect 663892 643136 663944 643142
rect 663892 643078 663944 643084
rect 663800 579964 663852 579970
rect 663800 579906 663852 579912
rect 663708 579828 663760 579834
rect 663708 579770 663760 579776
rect 663708 576904 663760 576910
rect 663708 576846 663760 576852
rect 661224 522504 661276 522510
rect 661224 522446 661276 522452
rect 661040 491428 661092 491434
rect 661040 491370 661092 491376
rect 660948 470824 661000 470830
rect 660948 470766 661000 470772
rect 658464 314628 658516 314634
rect 658464 314570 658516 314576
rect 660960 312050 660988 470766
rect 661040 416832 661092 416838
rect 661040 416774 661092 416780
rect 660948 312044 661000 312050
rect 660948 311986 661000 311992
rect 658372 311840 658424 311846
rect 658372 311782 658424 311788
rect 661052 267782 661080 416774
rect 661132 404048 661184 404054
rect 661132 403990 661184 403996
rect 661144 267986 661172 403990
rect 661236 403170 661264 522446
rect 663720 491570 663748 576846
rect 663800 549296 663852 549302
rect 663800 549238 663852 549244
rect 663708 491564 663760 491570
rect 663708 491506 663760 491512
rect 663708 430636 663760 430642
rect 663708 430578 663760 430584
rect 661224 403164 661276 403170
rect 661224 403106 661276 403112
rect 663720 268122 663748 430578
rect 663812 403306 663840 549238
rect 663904 535770 663932 643078
rect 666468 536444 666520 536450
rect 666468 536386 666520 536392
rect 663892 535764 663944 535770
rect 663892 535706 663944 535712
rect 663892 497684 663944 497690
rect 663892 497626 663944 497632
rect 663800 403300 663852 403306
rect 663800 403242 663852 403248
rect 663904 356250 663932 497626
rect 663984 444508 664036 444514
rect 663984 444450 664036 444456
rect 663892 356244 663944 356250
rect 663892 356186 663944 356192
rect 663996 312934 664024 444450
rect 666480 403442 666508 536386
rect 666468 403436 666520 403442
rect 666468 403378 666520 403384
rect 666468 389904 666520 389910
rect 666468 389846 666520 389852
rect 663984 312928 664036 312934
rect 663984 312870 664036 312876
rect 663708 268116 663760 268122
rect 663708 268058 663760 268064
rect 661132 267980 661184 267986
rect 661132 267922 661184 267928
rect 661040 267776 661092 267782
rect 661040 267718 661092 267724
rect 658280 265056 658332 265062
rect 658280 264998 658332 265004
rect 658186 262440 658242 262449
rect 658186 262375 658242 262384
rect 654140 231124 654192 231130
rect 654140 231066 654192 231072
rect 654152 226334 654180 231066
rect 656992 231056 657044 231062
rect 656992 230998 657044 231004
rect 656900 230988 656952 230994
rect 656900 230930 656952 230936
rect 654152 226306 655192 226334
rect 652852 222216 652904 222222
rect 652852 222158 652904 222164
rect 652760 219632 652812 219638
rect 652760 219574 652812 219580
rect 652760 219496 652812 219502
rect 652760 219438 652812 219444
rect 652668 219360 652720 219366
rect 652668 219302 652720 219308
rect 651656 218000 651708 218006
rect 651656 217942 651708 217948
rect 651564 216708 651616 216714
rect 651564 216650 651616 216656
rect 651288 212492 651340 212498
rect 651288 212434 651340 212440
rect 651380 212492 651432 212498
rect 651380 212434 651432 212440
rect 651392 210338 651420 212434
rect 650196 210310 650500 210338
rect 650196 210202 650224 210310
rect 649888 210174 650224 210202
rect 650472 210066 650500 210310
rect 651392 210310 651972 210338
rect 651392 210202 651420 210310
rect 651268 210174 651420 210202
rect 651944 210066 651972 210310
rect 652772 210202 652800 219438
rect 654140 219428 654192 219434
rect 654140 219370 654192 219376
rect 653048 210310 653352 210338
rect 653048 210202 653076 210310
rect 652740 210174 653076 210202
rect 653324 210066 653352 210310
rect 654152 210202 654180 219370
rect 654428 210310 654732 210338
rect 654428 210202 654456 210310
rect 654120 210174 654456 210202
rect 654704 210066 654732 210310
rect 655164 210066 655192 226306
rect 656912 215150 656940 230930
rect 656900 215144 656952 215150
rect 656900 215086 656952 215092
rect 655808 210310 656112 210338
rect 655808 210066 655836 210310
rect 642100 210038 642436 210052
rect 643480 210038 643816 210052
rect 644952 210038 645288 210052
rect 646332 210038 646668 210052
rect 647712 210038 648048 210066
rect 649092 210038 649428 210066
rect 650472 210038 650808 210066
rect 651944 210038 652280 210066
rect 653324 210038 653660 210066
rect 654704 210038 655040 210066
rect 655164 210038 655836 210066
rect 656084 210066 656112 210310
rect 657004 210202 657032 230998
rect 659752 230920 659804 230926
rect 659752 230862 659804 230868
rect 659660 230852 659712 230858
rect 659660 230794 659712 230800
rect 659672 215150 659700 230794
rect 657912 215144 657964 215150
rect 657912 215086 657964 215092
rect 659660 215144 659712 215150
rect 659660 215086 659712 215092
rect 657188 210310 657492 210338
rect 657188 210202 657216 210310
rect 656880 210174 657216 210202
rect 657464 210066 657492 210310
rect 657924 210066 657952 215086
rect 658568 210310 658872 210338
rect 658568 210066 658596 210310
rect 656084 210038 656420 210066
rect 657464 210038 657800 210066
rect 657924 210038 658596 210066
rect 658844 210066 658872 210310
rect 659764 210202 659792 230862
rect 662696 230784 662748 230790
rect 662696 230726 662748 230732
rect 662420 230716 662472 230722
rect 662420 230658 662472 230664
rect 660764 215144 660816 215150
rect 660764 215086 660816 215092
rect 660040 210310 660344 210338
rect 660040 210202 660068 210310
rect 659732 210174 660068 210202
rect 660316 210066 660344 210310
rect 660776 210066 660804 215086
rect 662432 210934 662460 230658
rect 662512 230648 662564 230654
rect 662512 230590 662564 230596
rect 662524 217938 662552 230590
rect 662604 230580 662656 230586
rect 662604 230522 662656 230528
rect 662616 218278 662644 230522
rect 662604 218272 662656 218278
rect 662604 218214 662656 218220
rect 662604 218136 662656 218142
rect 662604 218078 662656 218084
rect 662512 217932 662564 217938
rect 662512 217874 662564 217880
rect 662420 210928 662472 210934
rect 662420 210870 662472 210876
rect 661420 210310 661724 210338
rect 661420 210066 661448 210310
rect 658844 210038 659272 210066
rect 660316 210038 660652 210066
rect 660776 210038 661448 210066
rect 661696 210066 661724 210310
rect 662616 210202 662644 218078
rect 662708 211018 662736 230726
rect 662788 230512 662840 230518
rect 662788 230454 662840 230460
rect 662800 217954 662828 230454
rect 662880 230444 662932 230450
rect 662880 230386 662932 230392
rect 662892 218142 662920 230386
rect 666480 220862 666508 389846
rect 666468 220856 666520 220862
rect 666468 220798 666520 220804
rect 663984 218272 664036 218278
rect 663984 218214 664036 218220
rect 662880 218136 662932 218142
rect 662880 218078 662932 218084
rect 662800 217926 663564 217954
rect 662708 210990 663104 211018
rect 662696 210928 662748 210934
rect 662696 210870 662748 210876
rect 662492 210174 662644 210202
rect 662708 210066 662736 210870
rect 663076 210066 663104 210990
rect 663536 210066 663564 217926
rect 663996 210066 664024 218214
rect 664444 217932 664496 217938
rect 664444 217874 664496 217880
rect 664456 210066 664484 217874
rect 666192 215892 666244 215898
rect 666192 215834 666244 215840
rect 665272 215824 665324 215830
rect 665272 215766 665324 215772
rect 665284 210202 665312 215766
rect 665732 215756 665784 215762
rect 665732 215698 665784 215704
rect 665744 210202 665772 215698
rect 666204 210202 666232 215834
rect 665252 210174 665312 210202
rect 665712 210174 665772 210202
rect 666172 210174 666232 210202
rect 661696 210038 662032 210066
rect 662708 210038 662952 210066
rect 663076 210038 663412 210066
rect 663536 210038 663872 210066
rect 663996 210038 664332 210066
rect 664456 210038 664792 210066
rect 600044 209908 600096 209914
rect 600044 209850 600096 209856
rect 599950 208584 600006 208593
rect 599950 208519 600006 208528
rect 599858 207496 599914 207505
rect 599858 207431 599914 207440
rect 600056 206553 600084 209850
rect 601516 207120 601568 207126
rect 601516 207062 601568 207068
rect 601424 207052 601476 207058
rect 601424 206994 601476 207000
rect 600042 206544 600098 206553
rect 600042 206479 600098 206488
rect 599122 205456 599178 205465
rect 599122 205391 599178 205400
rect 582288 204332 582340 204338
rect 582288 204274 582340 204280
rect 599952 204332 600004 204338
rect 599952 204274 600004 204280
rect 580722 204096 580778 204105
rect 580722 204031 580778 204040
rect 580736 201550 580764 204031
rect 581090 202600 581146 202609
rect 581090 202535 581146 202544
rect 581104 201618 581132 202535
rect 599964 202473 599992 204274
rect 601436 203425 601464 206994
rect 601528 204513 601556 207062
rect 601514 204504 601570 204513
rect 601514 204439 601570 204448
rect 601422 203416 601478 203425
rect 601422 203351 601478 203360
rect 599950 202464 600006 202473
rect 599950 202399 600006 202408
rect 581092 201612 581144 201618
rect 581092 201554 581144 201560
rect 599952 201612 600004 201618
rect 599952 201554 600004 201560
rect 580724 201544 580776 201550
rect 580724 201486 580776 201492
rect 598940 201544 598992 201550
rect 598940 201486 598992 201492
rect 598952 201385 598980 201486
rect 598938 201376 598994 201385
rect 598938 201311 598994 201320
rect 581090 201104 581146 201113
rect 581090 201039 581146 201048
rect 581104 200122 581132 201039
rect 599964 200433 599992 201554
rect 599950 200424 600006 200433
rect 599950 200359 600006 200368
rect 581092 200116 581144 200122
rect 581092 200058 581144 200064
rect 599952 200116 600004 200122
rect 599952 200058 600004 200064
rect 582286 199608 582342 199617
rect 582286 199543 582342 199552
rect 582300 198762 582328 199543
rect 599964 199345 599992 200058
rect 599950 199336 600006 199345
rect 599950 199271 600006 199280
rect 582288 198756 582340 198762
rect 582288 198698 582340 198704
rect 599124 198756 599176 198762
rect 599124 198698 599176 198704
rect 599136 198393 599164 198698
rect 599122 198384 599178 198393
rect 599122 198319 599178 198328
rect 582286 197976 582342 197985
rect 582286 197911 582342 197920
rect 582300 197402 582328 197911
rect 582288 197396 582340 197402
rect 582288 197338 582340 197344
rect 599860 197396 599912 197402
rect 599860 197338 599912 197344
rect 580724 197328 580776 197334
rect 580724 197270 580776 197276
rect 580736 196489 580764 197270
rect 580722 196480 580778 196489
rect 580722 196415 580778 196424
rect 599872 196353 599900 197338
rect 599952 197328 600004 197334
rect 599950 197296 599952 197305
rect 600004 197296 600006 197305
rect 599950 197231 600006 197240
rect 599858 196344 599914 196353
rect 599858 196279 599914 196288
rect 599950 195256 600006 195265
rect 599950 195191 600006 195200
rect 582286 194984 582342 194993
rect 582286 194919 582342 194928
rect 582196 194676 582248 194682
rect 582196 194618 582248 194624
rect 582208 193497 582236 194618
rect 582300 194614 582328 194919
rect 599124 194676 599176 194682
rect 599124 194618 599176 194624
rect 582288 194608 582340 194614
rect 582288 194550 582340 194556
rect 599136 194313 599164 194618
rect 599964 194614 599992 195191
rect 599952 194608 600004 194614
rect 599952 194550 600004 194556
rect 599122 194304 599178 194313
rect 599122 194239 599178 194248
rect 582194 193488 582250 193497
rect 582194 193423 582250 193432
rect 599950 193216 600006 193225
rect 599950 193151 600006 193160
rect 599122 192264 599178 192273
rect 599122 192199 599178 192208
rect 582286 191992 582342 192001
rect 582286 191927 582342 191936
rect 582196 191888 582248 191894
rect 582196 191830 582248 191836
rect 582208 190505 582236 191830
rect 582300 191826 582328 191927
rect 599136 191894 599164 192199
rect 599124 191888 599176 191894
rect 599124 191830 599176 191836
rect 599964 191826 599992 193151
rect 582288 191820 582340 191826
rect 582288 191762 582340 191768
rect 599952 191820 600004 191826
rect 599952 191762 600004 191768
rect 599858 191176 599914 191185
rect 599858 191111 599914 191120
rect 582194 190496 582250 190505
rect 579804 190460 579856 190466
rect 599872 190466 599900 191111
rect 582194 190431 582250 190440
rect 599860 190460 599912 190466
rect 579804 190402 579856 190408
rect 599860 190402 599912 190408
rect 579816 188873 579844 190402
rect 600962 190224 601018 190233
rect 600962 190159 601018 190168
rect 579802 188864 579858 188873
rect 579802 188799 579858 188808
rect 582196 187672 582248 187678
rect 582196 187614 582248 187620
rect 582208 185881 582236 187614
rect 600976 187610 601004 190159
rect 601606 189136 601662 189145
rect 601606 189071 601662 189080
rect 601422 188184 601478 188193
rect 601422 188119 601478 188128
rect 582288 187604 582340 187610
rect 582288 187546 582340 187552
rect 600964 187604 601016 187610
rect 600964 187546 601016 187552
rect 582300 187377 582328 187546
rect 582286 187368 582342 187377
rect 582286 187303 582342 187312
rect 599950 187096 600006 187105
rect 599950 187031 600006 187040
rect 582194 185872 582250 185881
rect 582194 185807 582250 185816
rect 599858 185056 599914 185065
rect 599858 184991 599914 185000
rect 580264 184884 580316 184890
rect 580264 184826 580316 184832
rect 580276 182889 580304 184826
rect 580908 184816 580960 184822
rect 580908 184758 580960 184764
rect 580920 184385 580948 184758
rect 580906 184376 580962 184385
rect 580906 184311 580962 184320
rect 599766 184104 599822 184113
rect 599766 184039 599822 184048
rect 580262 182880 580318 182889
rect 580262 182815 580318 182824
rect 580632 182164 580684 182170
rect 580632 182106 580684 182112
rect 580540 182096 580592 182102
rect 580540 182038 580592 182044
rect 580552 179761 580580 182038
rect 580644 181393 580672 182106
rect 580630 181384 580686 181393
rect 580630 181319 580686 181328
rect 580538 179752 580594 179761
rect 580538 179687 580594 179696
rect 580724 179376 580776 179382
rect 580724 179318 580776 179324
rect 580736 176769 580764 179318
rect 599780 179314 599808 184039
rect 599872 182102 599900 184991
rect 599964 184890 599992 187031
rect 600042 186144 600098 186153
rect 600042 186079 600098 186088
rect 599952 184884 600004 184890
rect 599952 184826 600004 184832
rect 599950 183016 600006 183025
rect 599950 182951 600006 182960
rect 599860 182096 599912 182102
rect 599860 182038 599912 182044
rect 599858 180024 599914 180033
rect 599858 179959 599914 179968
rect 581092 179308 581144 179314
rect 581092 179250 581144 179256
rect 599768 179308 599820 179314
rect 599768 179250 599820 179256
rect 581104 178265 581132 179250
rect 599674 178936 599730 178945
rect 599674 178871 599730 178880
rect 581090 178256 581146 178265
rect 581090 178191 581146 178200
rect 598938 176896 598994 176905
rect 598938 176831 598994 176840
rect 580722 176760 580778 176769
rect 598952 176730 598980 176831
rect 580722 176695 580778 176704
rect 581000 176724 581052 176730
rect 581000 176666 581052 176672
rect 598940 176724 598992 176730
rect 598940 176666 598992 176672
rect 580816 173936 580868 173942
rect 580816 173878 580868 173884
rect 579712 173868 579764 173874
rect 579712 173810 579764 173816
rect 579724 172281 579752 173810
rect 579710 172272 579766 172281
rect 579710 172207 579766 172216
rect 579896 171148 579948 171154
rect 579896 171090 579948 171096
rect 579712 168564 579764 168570
rect 579712 168506 579764 168512
rect 579724 158545 579752 168506
rect 579908 161537 579936 171090
rect 580540 171012 580592 171018
rect 580540 170954 580592 170960
rect 580552 170649 580580 170954
rect 580538 170640 580594 170649
rect 580538 170575 580594 170584
rect 580172 168428 580224 168434
rect 580172 168370 580224 168376
rect 579894 161528 579950 161537
rect 579894 161463 579950 161472
rect 579710 158536 579766 158545
rect 579710 158471 579766 158480
rect 580184 157049 580212 168370
rect 580356 165708 580408 165714
rect 580356 165650 580408 165656
rect 580170 157040 580226 157049
rect 580170 156975 580226 156984
rect 580368 152425 580396 165650
rect 580828 164665 580856 173878
rect 581012 167657 581040 176666
rect 581460 176656 581512 176662
rect 581460 176598 581512 176604
rect 581472 175273 581500 176598
rect 581458 175264 581514 175273
rect 581458 175199 581514 175208
rect 582288 173800 582340 173806
rect 582286 173768 582288 173777
rect 582340 173768 582342 173777
rect 582286 173703 582342 173712
rect 582196 171216 582248 171222
rect 582196 171158 582248 171164
rect 582012 171080 582064 171086
rect 582012 171022 582064 171028
rect 582024 169153 582052 171022
rect 582010 169144 582066 169153
rect 582010 169079 582066 169088
rect 582104 168496 582156 168502
rect 582104 168438 582156 168444
rect 580998 167648 581054 167657
rect 580998 167583 581054 167592
rect 581276 165776 581328 165782
rect 581276 165718 581328 165724
rect 580814 164656 580870 164665
rect 580814 164591 580870 164600
rect 581000 162920 581052 162926
rect 581000 162862 581052 162868
rect 580908 160200 580960 160206
rect 580908 160142 580960 160148
rect 580540 160132 580592 160138
rect 580540 160074 580592 160080
rect 580354 152416 580410 152425
rect 580354 152351 580410 152360
rect 580552 146441 580580 160074
rect 580816 157412 580868 157418
rect 580816 157354 580868 157360
rect 580724 154624 580776 154630
rect 580724 154566 580776 154572
rect 580538 146432 580594 146441
rect 580538 146367 580594 146376
rect 580632 146328 580684 146334
rect 580632 146270 580684 146276
rect 579712 143608 579764 143614
rect 579712 143550 579764 143556
rect 579724 122097 579752 143550
rect 579804 138100 579856 138106
rect 579804 138042 579856 138048
rect 579710 122088 579766 122097
rect 579710 122023 579766 122032
rect 579816 112985 579844 138042
rect 580080 138032 580132 138038
rect 580080 137974 580132 137980
rect 579896 135312 579948 135318
rect 579896 135254 579948 135260
rect 579802 112976 579858 112985
rect 579802 112911 579858 112920
rect 579908 108497 579936 135254
rect 579988 132524 580040 132530
rect 579988 132466 580040 132472
rect 579894 108488 579950 108497
rect 579894 108423 579950 108432
rect 580000 105369 580028 132466
rect 580092 111489 580120 137974
rect 580172 135380 580224 135386
rect 580172 135322 580224 135328
rect 580078 111480 580134 111489
rect 580078 111415 580134 111424
rect 580184 106865 580212 135322
rect 580264 132592 580316 132598
rect 580264 132534 580316 132540
rect 580170 106856 580226 106865
rect 580170 106791 580226 106800
rect 579986 105360 580042 105369
rect 579986 105295 580042 105304
rect 580276 102377 580304 132534
rect 580356 129872 580408 129878
rect 580356 129814 580408 129820
rect 580262 102368 580318 102377
rect 580262 102303 580318 102312
rect 580368 100881 580396 129814
rect 580540 129804 580592 129810
rect 580540 129746 580592 129752
rect 580448 127016 580500 127022
rect 580448 126958 580500 126964
rect 580354 100872 580410 100881
rect 580354 100807 580410 100816
rect 580460 96257 580488 126958
rect 580552 97753 580580 129746
rect 580644 128217 580672 146270
rect 580736 138825 580764 154566
rect 580828 141817 580856 157354
rect 580814 141808 580870 141817
rect 580814 141743 580870 141752
rect 580920 140321 580948 160142
rect 581012 147937 581040 162862
rect 581184 160268 581236 160274
rect 581184 160210 581236 160216
rect 581092 157480 581144 157486
rect 581092 157422 581144 157428
rect 580998 147928 581054 147937
rect 580998 147863 581054 147872
rect 581104 143313 581132 157422
rect 581196 144945 581224 160210
rect 581288 154057 581316 165718
rect 581920 165640 581972 165646
rect 581920 165582 581972 165588
rect 581828 165572 581880 165578
rect 581828 165514 581880 165520
rect 581840 163169 581868 165514
rect 581826 163160 581882 163169
rect 581826 163095 581882 163104
rect 581460 162988 581512 162994
rect 581460 162930 581512 162936
rect 581274 154048 581330 154057
rect 581274 153983 581330 153992
rect 581472 149433 581500 162930
rect 581828 151904 581880 151910
rect 581828 151846 581880 151852
rect 581458 149424 581514 149433
rect 581458 149359 581514 149368
rect 581552 149184 581604 149190
rect 581552 149126 581604 149132
rect 581368 149116 581420 149122
rect 581368 149058 581420 149064
rect 581182 144936 581238 144945
rect 581182 144871 581238 144880
rect 581276 143676 581328 143682
rect 581276 143618 581328 143624
rect 581090 143304 581146 143313
rect 581090 143239 581146 143248
rect 581000 140888 581052 140894
rect 581000 140830 581052 140836
rect 580906 140312 580962 140321
rect 580906 140247 580962 140256
rect 580722 138816 580778 138825
rect 580722 138751 580778 138760
rect 580908 132660 580960 132666
rect 580908 132602 580960 132608
rect 580724 129940 580776 129946
rect 580724 129882 580776 129888
rect 580630 128208 580686 128217
rect 580630 128143 580686 128152
rect 580632 124228 580684 124234
rect 580632 124170 580684 124176
rect 580538 97744 580594 97753
rect 580538 97679 580594 97688
rect 580446 96248 580502 96257
rect 580446 96183 580502 96192
rect 578148 95328 578200 95334
rect 578148 95270 578200 95276
rect 575664 95260 575716 95266
rect 575664 95202 575716 95208
rect 571340 53576 571392 53582
rect 571340 53518 571392 53524
rect 84824 52686 85160 52714
rect 52276 47116 52328 47122
rect 52276 47058 52328 47064
rect 85132 45694 85160 52686
rect 150314 52454 150342 52700
rect 215832 52686 216168 52714
rect 281336 52686 281488 52714
rect 150268 52426 150342 52454
rect 150268 48414 150296 52426
rect 213828 51060 213880 51066
rect 213828 51002 213880 51008
rect 149244 48408 149296 48414
rect 149244 48350 149296 48356
rect 150256 48408 150308 48414
rect 150256 48350 150308 48356
rect 149256 47122 149284 48350
rect 149244 47116 149296 47122
rect 149244 47058 149296 47064
rect 141804 46702 142370 46730
rect 85120 45688 85172 45694
rect 85120 45630 85172 45636
rect 52184 42900 52236 42906
rect 52184 42842 52236 42848
rect 141804 41546 141832 46702
rect 212448 45552 212500 45558
rect 212448 45494 212500 45500
rect 209688 43308 209740 43314
rect 209688 43250 209740 43256
rect 187606 41848 187662 41857
rect 187358 41806 187606 41834
rect 194414 41848 194470 41857
rect 194074 41806 194414 41834
rect 187606 41783 187662 41792
rect 194414 41783 194470 41792
rect 209700 41546 209728 43250
rect 141792 41540 141844 41546
rect 141792 41482 141844 41488
rect 207020 41540 207072 41546
rect 207020 41482 207072 41488
rect 209688 41540 209740 41546
rect 209688 41482 209740 41488
rect 141804 40202 141832 41482
rect 141758 40174 141832 40202
rect 141758 39984 141786 40174
rect 207032 17490 207060 41482
rect 212460 41313 212488 45494
rect 209778 41304 209834 41313
rect 209778 41239 209834 41248
rect 212446 41304 212502 41313
rect 212446 41239 212502 41248
rect 209792 17490 209820 41239
rect 213840 24818 213868 51002
rect 216140 48346 216168 52686
rect 218060 48408 218112 48414
rect 218060 48350 218112 48356
rect 216128 48340 216180 48346
rect 216128 48282 216180 48288
rect 218072 46918 218100 48350
rect 281460 48249 281488 52686
rect 346504 52686 346900 52714
rect 412344 52686 412680 52714
rect 477848 52686 478184 52714
rect 346504 51066 346532 52686
rect 346872 52426 346900 52686
rect 346860 52420 346912 52426
rect 346860 52362 346912 52368
rect 346492 51060 346544 51066
rect 346492 51002 346544 51008
rect 412652 48414 412680 52686
rect 478156 48482 478184 52686
rect 543016 52686 543352 52714
rect 478144 48476 478196 48482
rect 478144 48418 478196 48424
rect 518808 48476 518860 48482
rect 518808 48418 518860 48424
rect 412640 48408 412692 48414
rect 412640 48350 412692 48356
rect 494060 48408 494112 48414
rect 494060 48350 494112 48356
rect 281446 48240 281502 48249
rect 281446 48175 281502 48184
rect 218060 46912 218112 46918
rect 218060 46854 218112 46860
rect 215300 42900 215352 42906
rect 215300 42842 215352 42848
rect 213184 24812 213236 24818
rect 213184 24754 213236 24760
rect 213828 24812 213880 24818
rect 213828 24754 213880 24760
rect 213196 17490 213224 24754
rect 207032 17462 207184 17490
rect 209792 17462 210036 17490
rect 212888 17462 213224 17490
rect 215312 17490 215340 42842
rect 218072 33134 218100 46854
rect 494072 46850 494100 48350
rect 494060 46844 494112 46850
rect 494060 46786 494112 46792
rect 502248 46844 502300 46850
rect 502248 46786 502300 46792
rect 460664 45892 460716 45898
rect 460664 45834 460716 45840
rect 367100 45824 367152 45830
rect 367100 45766 367152 45772
rect 311900 45756 311952 45762
rect 311900 45698 311952 45704
rect 233148 45620 233200 45626
rect 233148 45562 233200 45568
rect 230940 43920 230992 43926
rect 230940 43862 230992 43868
rect 230388 43852 230440 43858
rect 230388 43794 230440 43800
rect 226248 43444 226300 43450
rect 226248 43386 226300 43392
rect 223488 43376 223540 43382
rect 223488 43318 223540 43324
rect 218072 33106 218192 33134
rect 218164 17490 218192 33106
rect 223500 22574 223528 43318
rect 226260 23050 226288 43386
rect 224592 23044 224644 23050
rect 224592 22986 224644 22992
rect 226248 23044 226300 23050
rect 226248 22986 226300 22992
rect 221740 22568 221792 22574
rect 221740 22510 221792 22516
rect 223488 22568 223540 22574
rect 223488 22510 223540 22516
rect 221752 17490 221780 22510
rect 224604 17490 224632 22986
rect 215312 17462 215740 17490
rect 218164 17462 218592 17490
rect 221444 17462 221780 17490
rect 224296 17462 224632 17490
rect 230400 7721 230428 43794
rect 230756 43784 230808 43790
rect 230756 43726 230808 43732
rect 230572 43648 230624 43654
rect 230572 43590 230624 43596
rect 230480 43580 230532 43586
rect 230480 43522 230532 43528
rect 230492 9217 230520 43522
rect 230584 12209 230612 43590
rect 230664 43512 230716 43518
rect 230664 43454 230716 43460
rect 230570 12200 230626 12209
rect 230570 12135 230626 12144
rect 230676 10713 230704 43454
rect 230768 13705 230796 43726
rect 230848 43716 230900 43722
rect 230848 43658 230900 43664
rect 230860 15201 230888 43658
rect 230952 16697 230980 43862
rect 230938 16688 230994 16697
rect 230938 16623 230994 16632
rect 230846 15192 230902 15201
rect 230846 15127 230902 15136
rect 230754 13696 230810 13705
rect 230754 13631 230810 13640
rect 230662 10704 230718 10713
rect 230662 10639 230718 10648
rect 230478 9208 230534 9217
rect 230478 9143 230534 9152
rect 230386 7712 230442 7721
rect 230386 7647 230442 7656
rect 233160 6526 233188 45562
rect 311912 44198 311940 45698
rect 367112 44198 367140 45766
rect 311900 44192 311952 44198
rect 311900 44134 311952 44140
rect 367100 44192 367152 44198
rect 367100 44134 367152 44140
rect 310428 44124 310480 44130
rect 310428 44066 310480 44072
rect 365168 44124 365220 44130
rect 365168 44066 365220 44072
rect 310440 42106 310468 44066
rect 365180 42106 365208 44066
rect 419724 44056 419776 44062
rect 419724 43998 419776 44004
rect 405556 43988 405608 43994
rect 405556 43930 405608 43936
rect 310132 42078 310468 42106
rect 364918 42078 365208 42106
rect 405568 42092 405596 43930
rect 419736 42772 419764 43998
rect 455420 42288 455472 42294
rect 455420 42230 455472 42236
rect 307298 41848 307354 41857
rect 307004 41806 307298 41834
rect 362038 41848 362094 41857
rect 361790 41806 362038 41834
rect 307298 41783 307354 41792
rect 415490 41848 415546 41857
rect 415426 41806 415490 41834
rect 362038 41783 362094 41792
rect 416622 41818 416728 41834
rect 416622 41812 416740 41818
rect 416622 41806 416688 41812
rect 415490 41783 415546 41792
rect 416688 41754 416740 41760
rect 420736 41812 420788 41818
rect 420736 41754 420788 41760
rect 420748 38622 420776 41754
rect 455432 38622 455460 42230
rect 460676 42106 460704 45834
rect 475660 45688 475712 45694
rect 475660 45630 475712 45636
rect 474464 44124 474516 44130
rect 474464 44066 474516 44072
rect 474476 42500 474504 44066
rect 460368 42078 460704 42106
rect 470052 41984 470108 41993
rect 470052 41919 470108 41928
rect 470066 41820 470094 41919
rect 471408 41818 471744 41834
rect 471408 41812 471756 41818
rect 471408 41806 471704 41812
rect 471704 41754 471756 41760
rect 475568 41812 475620 41818
rect 475568 41754 475620 41760
rect 420736 38616 420788 38622
rect 420736 38558 420788 38564
rect 455420 38616 455472 38622
rect 455420 38558 455472 38564
rect 475580 38554 475608 41754
rect 475672 38622 475700 45630
rect 502260 41886 502288 46786
rect 518820 44305 518848 48418
rect 521844 48340 521896 48346
rect 521844 48282 521896 48288
rect 518806 44296 518862 44305
rect 518806 44231 518862 44240
rect 510620 42220 510672 42226
rect 510620 42162 510672 42168
rect 502248 41880 502300 41886
rect 502248 41822 502300 41828
rect 510632 38690 510660 42162
rect 520462 42120 520518 42129
rect 520518 42078 520674 42106
rect 521856 42092 521884 48282
rect 540888 45688 540940 45694
rect 540888 45630 540940 45636
rect 526166 44160 526222 44169
rect 526166 44095 526222 44104
rect 526180 42092 526208 44095
rect 540900 44062 540928 45630
rect 540888 44056 540940 44062
rect 540888 43998 540940 44004
rect 530688 42362 531084 42378
rect 530676 42356 531096 42362
rect 530728 42350 531044 42356
rect 530676 42298 530728 42304
rect 531044 42298 531096 42304
rect 530688 42226 531084 42242
rect 530676 42220 531096 42226
rect 530728 42214 531044 42220
rect 530676 42162 530728 42168
rect 531044 42162 531096 42168
rect 520462 42055 520518 42064
rect 518532 41880 518584 41886
rect 514864 41818 515154 41834
rect 518584 41828 518834 41834
rect 518532 41822 518834 41828
rect 514024 41812 514076 41818
rect 514024 41754 514076 41760
rect 514852 41812 515154 41818
rect 514904 41806 515154 41812
rect 518544 41806 518834 41822
rect 529322 41818 529704 41834
rect 529322 41812 529716 41818
rect 529322 41806 529664 41812
rect 514852 41754 514904 41760
rect 529664 41754 529716 41760
rect 530216 41812 530268 41818
rect 530216 41754 530268 41760
rect 505652 38684 505704 38690
rect 505652 38626 505704 38632
rect 510620 38684 510672 38690
rect 510620 38626 510672 38632
rect 475660 38616 475712 38622
rect 475660 38558 475712 38564
rect 505664 38554 505692 38626
rect 514036 38622 514064 41754
rect 530228 41313 530256 41754
rect 543016 41313 543044 52686
rect 552020 48340 552072 48346
rect 552020 48282 552072 48288
rect 552032 41857 552060 48282
rect 563612 44192 563664 44198
rect 563612 44134 563664 44140
rect 552018 41848 552074 41857
rect 552018 41783 552074 41792
rect 563624 41721 563652 44134
rect 571352 41993 571380 53518
rect 575676 48346 575704 95202
rect 575664 48340 575716 48346
rect 575664 48282 575716 48288
rect 574836 46980 574888 46986
rect 574836 46922 574888 46928
rect 574848 42294 574876 46922
rect 578160 44198 578188 95270
rect 580644 93265 580672 124170
rect 580736 99385 580764 129882
rect 580816 127084 580868 127090
rect 580816 127026 580868 127032
rect 580722 99376 580778 99385
rect 580722 99311 580778 99320
rect 580828 94761 580856 127026
rect 580920 103873 580948 132602
rect 581012 115977 581040 140830
rect 581184 140820 581236 140826
rect 581184 140762 581236 140768
rect 581092 138168 581144 138174
rect 581092 138110 581144 138116
rect 580998 115968 581054 115977
rect 580998 115903 581054 115912
rect 581000 110492 581052 110498
rect 581000 110434 581052 110440
rect 580906 103864 580962 103873
rect 580906 103799 580962 103808
rect 580908 99408 580960 99414
rect 580908 99350 580960 99356
rect 580814 94752 580870 94761
rect 580814 94687 580870 94696
rect 580630 93256 580686 93265
rect 580630 93191 580686 93200
rect 579620 82680 579672 82686
rect 579618 82648 579620 82657
rect 579672 82648 579674 82657
rect 579618 82583 579674 82592
rect 580540 66224 580592 66230
rect 580540 66166 580592 66172
rect 580552 65929 580580 66166
rect 580538 65920 580594 65929
rect 580538 65855 580594 65864
rect 578240 60716 578292 60722
rect 578240 60658 578292 60664
rect 578252 46986 578280 60658
rect 579620 60512 579672 60518
rect 579620 60454 579672 60460
rect 579632 59809 579660 60454
rect 579618 59800 579674 59809
rect 579618 59735 579674 59744
rect 579620 58676 579672 58682
rect 579620 58618 579672 58624
rect 579632 58313 579660 58618
rect 579618 58304 579674 58313
rect 579618 58239 579674 58248
rect 580920 53825 580948 99350
rect 581012 70417 581040 110434
rect 581104 109993 581132 138110
rect 581196 114481 581224 140762
rect 581288 120601 581316 143618
rect 581380 126721 581408 149058
rect 581460 146396 581512 146402
rect 581460 146338 581512 146344
rect 581366 126712 581422 126721
rect 581366 126647 581422 126656
rect 581472 123593 581500 146338
rect 581564 125089 581592 149126
rect 581736 143744 581788 143750
rect 581736 143686 581788 143692
rect 581644 140956 581696 140962
rect 581644 140898 581696 140904
rect 581550 125080 581606 125089
rect 581550 125015 581606 125024
rect 581458 123584 581514 123593
rect 581458 123519 581514 123528
rect 581274 120592 581330 120601
rect 581274 120527 581330 120536
rect 581552 118720 581604 118726
rect 581552 118662 581604 118668
rect 581276 116000 581328 116006
rect 581276 115942 581328 115948
rect 581182 114472 581238 114481
rect 581182 114407 581238 114416
rect 581090 109984 581146 109993
rect 581090 109919 581146 109928
rect 581184 107704 581236 107710
rect 581184 107646 581236 107652
rect 581092 104916 581144 104922
rect 581092 104858 581144 104864
rect 580998 70408 581054 70417
rect 580998 70343 581054 70352
rect 581104 64433 581132 104858
rect 581196 67425 581224 107646
rect 581288 78033 581316 115942
rect 581460 113212 581512 113218
rect 581460 113154 581512 113160
rect 581368 110560 581420 110566
rect 581368 110502 581420 110508
rect 581274 78024 581330 78033
rect 581274 77959 581330 77968
rect 581380 72049 581408 110502
rect 581472 76537 581500 113154
rect 581564 81161 581592 118662
rect 581656 117609 581684 140898
rect 581748 119105 581776 143686
rect 581840 131209 581868 151846
rect 581932 150929 581960 165582
rect 582012 157548 582064 157554
rect 582012 157490 582064 157496
rect 581918 150920 581974 150929
rect 581918 150855 581974 150864
rect 581920 149252 581972 149258
rect 581920 149194 581972 149200
rect 581826 131200 581882 131209
rect 581826 131135 581882 131144
rect 581932 129713 581960 149194
rect 582024 137329 582052 157490
rect 582116 155553 582144 168438
rect 582208 160041 582236 171158
rect 599688 171018 599716 178871
rect 599766 177984 599822 177993
rect 599766 177919 599822 177928
rect 599780 171086 599808 177919
rect 599872 173874 599900 179959
rect 599964 179382 599992 182951
rect 600056 182170 600084 186079
rect 601436 184822 601464 188119
rect 601620 187678 601648 189071
rect 601608 187672 601660 187678
rect 601608 187614 601660 187620
rect 601424 184816 601476 184822
rect 601424 184758 601476 184764
rect 600044 182164 600096 182170
rect 600044 182106 600096 182112
rect 600042 182064 600098 182073
rect 600042 181999 600098 182008
rect 599952 179376 600004 179382
rect 599952 179318 600004 179324
rect 600056 176662 600084 181999
rect 600134 180976 600190 180985
rect 600134 180911 600190 180920
rect 600044 176656 600096 176662
rect 600044 176598 600096 176604
rect 599950 174856 600006 174865
rect 599950 174791 600006 174800
rect 599964 173942 599992 174791
rect 599952 173936 600004 173942
rect 599952 173878 600004 173884
rect 599860 173868 599912 173874
rect 599860 173810 599912 173816
rect 600148 173806 600176 180911
rect 600318 175944 600374 175953
rect 600318 175879 600374 175888
rect 600136 173800 600188 173806
rect 600136 173742 600188 173748
rect 599858 172816 599914 172825
rect 599858 172751 599914 172760
rect 599872 171154 599900 172751
rect 599950 171864 600006 171873
rect 599950 171799 600006 171808
rect 599964 171222 599992 171799
rect 599952 171216 600004 171222
rect 599952 171158 600004 171164
rect 599860 171148 599912 171154
rect 599860 171090 599912 171096
rect 599768 171080 599820 171086
rect 599768 171022 599820 171028
rect 599676 171012 599728 171018
rect 599676 170954 599728 170960
rect 599950 170776 600006 170785
rect 599950 170711 600006 170720
rect 599766 169824 599822 169833
rect 599766 169759 599822 169768
rect 599030 168736 599086 168745
rect 599030 168671 599086 168680
rect 599044 168502 599072 168671
rect 599032 168496 599084 168502
rect 599032 168438 599084 168444
rect 599780 168434 599808 169759
rect 599964 168570 599992 170711
rect 599952 168564 600004 168570
rect 599952 168506 600004 168512
rect 599768 168428 599820 168434
rect 599768 168370 599820 168376
rect 600332 168366 600360 175879
rect 601146 173904 601202 173913
rect 601146 173839 601202 173848
rect 582288 168360 582340 168366
rect 582288 168302 582340 168308
rect 600320 168360 600372 168366
rect 600320 168302 600372 168308
rect 582300 166161 582328 168302
rect 599858 167784 599914 167793
rect 599858 167719 599914 167728
rect 582286 166152 582342 166161
rect 582286 166087 582342 166096
rect 599872 165782 599900 167719
rect 600042 166696 600098 166705
rect 600042 166631 600098 166640
rect 599860 165776 599912 165782
rect 599860 165718 599912 165724
rect 599950 165744 600006 165753
rect 600056 165714 600084 166631
rect 599950 165679 600006 165688
rect 600044 165708 600096 165714
rect 599964 165646 599992 165679
rect 600044 165650 600096 165656
rect 599952 165640 600004 165646
rect 599952 165582 600004 165588
rect 601160 165578 601188 173839
rect 601148 165572 601200 165578
rect 601148 165514 601200 165520
rect 599858 164656 599914 164665
rect 599858 164591 599914 164600
rect 599872 162994 599900 164591
rect 599950 163704 600006 163713
rect 599950 163639 600006 163648
rect 599860 162988 599912 162994
rect 599860 162930 599912 162936
rect 599964 162926 599992 163639
rect 599952 162920 600004 162926
rect 599952 162862 600004 162868
rect 599858 162616 599914 162625
rect 599858 162551 599914 162560
rect 599872 160138 599900 162551
rect 600042 161664 600098 161673
rect 600042 161599 600098 161608
rect 599950 160576 600006 160585
rect 599950 160511 600006 160520
rect 599964 160206 599992 160511
rect 600056 160274 600084 161599
rect 600044 160268 600096 160274
rect 600044 160210 600096 160216
rect 599952 160200 600004 160206
rect 599952 160142 600004 160148
rect 599860 160132 599912 160138
rect 599860 160074 599912 160080
rect 582194 160032 582250 160041
rect 582194 159967 582250 159976
rect 598938 159624 598994 159633
rect 598938 159559 598994 159568
rect 598952 157418 598980 159559
rect 599858 158536 599914 158545
rect 599858 158471 599914 158480
rect 599872 157486 599900 158471
rect 599950 157584 600006 157593
rect 599950 157519 599952 157528
rect 600004 157519 600006 157528
rect 599952 157490 600004 157496
rect 599860 157480 599912 157486
rect 599860 157422 599912 157428
rect 598940 157412 598992 157418
rect 598940 157354 598992 157360
rect 599858 156496 599914 156505
rect 599858 156431 599914 156440
rect 582102 155544 582158 155553
rect 582102 155479 582158 155488
rect 582196 154692 582248 154698
rect 582196 154634 582248 154640
rect 582104 151836 582156 151842
rect 582104 151778 582156 151784
rect 582010 137320 582066 137329
rect 582010 137255 582066 137264
rect 582116 134201 582144 151778
rect 582208 135833 582236 154634
rect 599872 154630 599900 156431
rect 599950 155544 600006 155553
rect 599950 155479 600006 155488
rect 599964 154698 599992 155479
rect 599952 154692 600004 154698
rect 599952 154634 600004 154640
rect 599860 154624 599912 154630
rect 599860 154566 599912 154572
rect 600042 154456 600098 154465
rect 600042 154391 600098 154400
rect 599858 153504 599914 153513
rect 599858 153439 599914 153448
rect 599872 151978 599900 153439
rect 599950 152416 600006 152425
rect 599950 152351 600006 152360
rect 582288 151972 582340 151978
rect 582288 151914 582340 151920
rect 599860 151972 599912 151978
rect 599860 151914 599912 151920
rect 582194 135824 582250 135833
rect 582194 135759 582250 135768
rect 582102 134192 582158 134201
rect 582102 134127 582158 134136
rect 582300 132705 582328 151914
rect 599964 151910 599992 152351
rect 599952 151904 600004 151910
rect 599952 151846 600004 151852
rect 600056 151842 600084 154391
rect 600044 151836 600096 151842
rect 600044 151778 600096 151784
rect 598938 151464 598994 151473
rect 598938 151399 598994 151408
rect 598952 149258 598980 151399
rect 599858 150376 599914 150385
rect 599858 150311 599914 150320
rect 598940 149252 598992 149258
rect 598940 149194 598992 149200
rect 599872 149190 599900 150311
rect 599950 149424 600006 149433
rect 599950 149359 600006 149368
rect 599860 149184 599912 149190
rect 599860 149126 599912 149132
rect 599964 149122 599992 149359
rect 599952 149116 600004 149122
rect 599952 149058 600004 149064
rect 599858 148336 599914 148345
rect 599858 148271 599914 148280
rect 599872 146334 599900 148271
rect 599950 147384 600006 147393
rect 599950 147319 600006 147328
rect 599964 146402 599992 147319
rect 599952 146396 600004 146402
rect 599952 146338 600004 146344
rect 599860 146328 599912 146334
rect 599860 146270 599912 146276
rect 600042 146296 600098 146305
rect 600042 146231 600098 146240
rect 599858 145344 599914 145353
rect 599858 145279 599914 145288
rect 599872 143682 599900 145279
rect 599950 144256 600006 144265
rect 599950 144191 600006 144200
rect 599964 143750 599992 144191
rect 599952 143744 600004 143750
rect 599952 143686 600004 143692
rect 599860 143676 599912 143682
rect 599860 143618 599912 143624
rect 600056 143614 600084 146231
rect 600044 143608 600096 143614
rect 600044 143550 600096 143556
rect 599858 143304 599914 143313
rect 599858 143239 599914 143248
rect 599306 141264 599362 141273
rect 599306 141199 599362 141208
rect 599320 140826 599348 141199
rect 599872 140962 599900 143239
rect 599950 142216 600006 142225
rect 599950 142151 600006 142160
rect 599860 140956 599912 140962
rect 599860 140898 599912 140904
rect 599964 140894 599992 142151
rect 599952 140888 600004 140894
rect 599952 140830 600004 140836
rect 599308 140820 599360 140826
rect 599308 140762 599360 140768
rect 599858 140176 599914 140185
rect 599858 140111 599914 140120
rect 599766 139224 599822 139233
rect 599766 139159 599822 139168
rect 599780 138038 599808 139159
rect 599872 138106 599900 140111
rect 599952 138168 600004 138174
rect 599950 138136 599952 138145
rect 600004 138136 600006 138145
rect 599860 138100 599912 138106
rect 599950 138071 600006 138080
rect 599860 138042 599912 138048
rect 599768 138032 599820 138038
rect 599768 137974 599820 137980
rect 599858 137184 599914 137193
rect 599858 137119 599914 137128
rect 599872 135318 599900 137119
rect 599950 136096 600006 136105
rect 599950 136031 600006 136040
rect 599964 135386 599992 136031
rect 599952 135380 600004 135386
rect 599952 135322 600004 135328
rect 599860 135312 599912 135318
rect 599860 135254 599912 135260
rect 600042 135144 600098 135153
rect 600042 135079 600098 135088
rect 599858 134056 599914 134065
rect 599858 133991 599914 134000
rect 582286 132696 582342 132705
rect 599872 132666 599900 133991
rect 599950 133104 600006 133113
rect 599950 133039 600006 133048
rect 582286 132631 582342 132640
rect 599860 132660 599912 132666
rect 599860 132602 599912 132608
rect 599964 132598 599992 133039
rect 599952 132592 600004 132598
rect 599952 132534 600004 132540
rect 600056 132530 600084 135079
rect 600044 132524 600096 132530
rect 600044 132466 600096 132472
rect 599858 132016 599914 132025
rect 599858 131951 599914 131960
rect 599766 131064 599822 131073
rect 599766 130999 599822 131008
rect 599780 129946 599808 130999
rect 599768 129940 599820 129946
rect 599768 129882 599820 129888
rect 599872 129878 599900 131951
rect 599950 129976 600006 129985
rect 599950 129911 600006 129920
rect 599860 129872 599912 129878
rect 599860 129814 599912 129820
rect 599964 129810 599992 129911
rect 599952 129804 600004 129810
rect 599952 129746 600004 129752
rect 581918 129704 581974 129713
rect 581918 129639 581974 129648
rect 599858 129024 599914 129033
rect 599858 128959 599914 128968
rect 599872 127022 599900 128959
rect 599950 127936 600006 127945
rect 599950 127871 600006 127880
rect 599964 127090 599992 127871
rect 599952 127084 600004 127090
rect 599952 127026 600004 127032
rect 599860 127016 599912 127022
rect 599766 126984 599822 126993
rect 599860 126958 599912 126964
rect 599766 126919 599822 126928
rect 582288 124364 582340 124370
rect 582288 124306 582340 124312
rect 582012 124296 582064 124302
rect 582012 124238 582064 124244
rect 581920 121576 581972 121582
rect 581920 121518 581972 121524
rect 581734 119096 581790 119105
rect 581734 119031 581790 119040
rect 581828 118788 581880 118794
rect 581828 118730 581880 118736
rect 581642 117600 581698 117609
rect 581642 117535 581698 117544
rect 581736 116068 581788 116074
rect 581736 116010 581788 116016
rect 581644 113280 581696 113286
rect 581644 113222 581696 113228
rect 581550 81152 581606 81161
rect 581550 81087 581606 81096
rect 581458 76528 581514 76537
rect 581458 76463 581514 76472
rect 581656 75041 581684 113222
rect 581748 79529 581776 116010
rect 581840 84153 581868 118730
rect 581932 85649 581960 121518
rect 582024 90273 582052 124238
rect 582104 121644 582156 121650
rect 582104 121586 582156 121592
rect 582010 90264 582066 90273
rect 582010 90199 582066 90208
rect 582116 87145 582144 121586
rect 582196 121508 582248 121514
rect 582196 121450 582248 121456
rect 582208 88641 582236 121450
rect 582300 91769 582328 124306
rect 599780 124234 599808 126919
rect 600042 125896 600098 125905
rect 600042 125831 600098 125840
rect 599950 124944 600006 124953
rect 599950 124879 600006 124888
rect 599964 124302 599992 124879
rect 600056 124370 600084 125831
rect 600044 124364 600096 124370
rect 600044 124306 600096 124312
rect 599952 124296 600004 124302
rect 599952 124238 600004 124244
rect 599768 124228 599820 124234
rect 599768 124170 599820 124176
rect 600042 123856 600098 123865
rect 600042 123791 600098 123800
rect 599858 122904 599914 122913
rect 599858 122839 599914 122848
rect 599872 121650 599900 122839
rect 599950 121816 600006 121825
rect 599950 121751 600006 121760
rect 599860 121644 599912 121650
rect 599860 121586 599912 121592
rect 599964 121582 599992 121751
rect 599952 121576 600004 121582
rect 599952 121518 600004 121524
rect 600056 121514 600084 123791
rect 600044 121508 600096 121514
rect 600044 121450 600096 121456
rect 600042 120864 600098 120873
rect 600042 120799 600098 120808
rect 599950 119776 600006 119785
rect 599950 119711 600006 119720
rect 599964 118862 599992 119711
rect 583668 118856 583720 118862
rect 599952 118856 600004 118862
rect 583668 118798 583720 118804
rect 599858 118824 599914 118833
rect 582286 91760 582342 91769
rect 582286 91695 582342 91704
rect 582194 88632 582250 88641
rect 582194 88567 582250 88576
rect 582102 87136 582158 87145
rect 582102 87071 582158 87080
rect 581918 85640 581974 85649
rect 581918 85575 581974 85584
rect 582288 84448 582340 84454
rect 582288 84390 582340 84396
rect 582196 84380 582248 84386
rect 582196 84322 582248 84328
rect 582012 84312 582064 84318
rect 582012 84254 582064 84260
rect 581920 84176 581972 84182
rect 581826 84144 581882 84153
rect 581920 84118 581972 84124
rect 581826 84079 581882 84088
rect 581734 79520 581790 79529
rect 581734 79455 581790 79464
rect 581642 75032 581698 75041
rect 581642 74967 581698 74976
rect 581366 72040 581422 72049
rect 581366 71975 581422 71984
rect 581182 67416 581238 67425
rect 581182 67351 581238 67360
rect 581090 64424 581146 64433
rect 581090 64359 581146 64368
rect 581932 56817 581960 84118
rect 582024 62937 582052 84254
rect 582104 84244 582156 84250
rect 582104 84186 582156 84192
rect 582010 62928 582066 62937
rect 582010 62863 582066 62872
rect 581918 56808 581974 56817
rect 581918 56743 581974 56752
rect 582116 55321 582144 84186
rect 582208 61305 582236 84322
rect 582300 68921 582328 84390
rect 583680 82686 583708 118798
rect 599952 118798 600004 118804
rect 600056 118794 600084 120799
rect 599858 118759 599914 118768
rect 600044 118788 600096 118794
rect 599872 118726 599900 118759
rect 600044 118730 600096 118736
rect 599860 118720 599912 118726
rect 599860 118662 599912 118668
rect 599858 117736 599914 117745
rect 599858 117671 599914 117680
rect 599872 116074 599900 117671
rect 599950 116784 600006 116793
rect 599950 116719 600006 116728
rect 599860 116068 599912 116074
rect 599860 116010 599912 116016
rect 599964 116006 599992 116719
rect 599952 116000 600004 116006
rect 599952 115942 600004 115948
rect 599858 115696 599914 115705
rect 599858 115631 599914 115640
rect 599872 113218 599900 115631
rect 599950 114744 600006 114753
rect 599950 114679 600006 114688
rect 599964 113286 599992 114679
rect 599952 113280 600004 113286
rect 599952 113222 600004 113228
rect 599860 113212 599912 113218
rect 599860 113154 599912 113160
rect 599950 112704 600006 112713
rect 599950 112639 600006 112648
rect 599766 111616 599822 111625
rect 599766 111551 599822 111560
rect 599780 110498 599808 111551
rect 599964 110566 599992 112639
rect 600226 110664 600282 110673
rect 600226 110599 600282 110608
rect 599952 110560 600004 110566
rect 599952 110502 600004 110508
rect 599768 110492 599820 110498
rect 599768 110434 599820 110440
rect 599950 109576 600006 109585
rect 599950 109511 600006 109520
rect 599964 107710 599992 109511
rect 599952 107704 600004 107710
rect 599952 107646 600004 107652
rect 599950 107536 600006 107545
rect 599950 107471 600006 107480
rect 599964 104922 599992 107471
rect 599952 104916 600004 104922
rect 599952 104858 600004 104864
rect 599950 100464 600006 100473
rect 599950 100399 600006 100408
rect 599964 99414 599992 100399
rect 599952 99408 600004 99414
rect 599952 99350 600004 99356
rect 596180 95396 596232 95402
rect 596180 95338 596232 95344
rect 586428 84652 586480 84658
rect 586428 84594 586480 84600
rect 583852 84584 583904 84590
rect 583852 84526 583904 84532
rect 583760 84516 583812 84522
rect 583760 84458 583812 84464
rect 583668 82680 583720 82686
rect 583668 82622 583720 82628
rect 582286 68912 582342 68921
rect 582286 68847 582342 68856
rect 583668 66292 583720 66298
rect 583668 66234 583720 66240
rect 582194 61296 582250 61305
rect 582194 61231 582250 61240
rect 583680 60790 583708 66234
rect 583668 60784 583720 60790
rect 583668 60726 583720 60732
rect 583772 60518 583800 84458
rect 583760 60512 583812 60518
rect 583760 60454 583812 60460
rect 583864 58682 583892 84526
rect 586440 66230 586468 84594
rect 596192 80850 596220 95338
rect 600240 84454 600268 110599
rect 600318 108624 600374 108633
rect 600318 108559 600374 108568
rect 600332 84658 600360 108559
rect 600594 106584 600650 106593
rect 600594 106519 600650 106528
rect 600410 105496 600466 105505
rect 600410 105431 600466 105440
rect 600320 84652 600372 84658
rect 600320 84594 600372 84600
rect 600228 84448 600280 84454
rect 600228 84390 600280 84396
rect 600424 84386 600452 105431
rect 600502 103456 600558 103465
rect 600502 103391 600558 103400
rect 600516 84590 600544 103391
rect 600504 84584 600556 84590
rect 600504 84526 600556 84532
rect 600412 84380 600464 84386
rect 600412 84322 600464 84328
rect 600608 84318 600636 106519
rect 600686 104544 600742 104553
rect 600686 104479 600742 104488
rect 600700 84522 600728 104479
rect 600870 102504 600926 102513
rect 600870 102439 600926 102448
rect 600778 101416 600834 101425
rect 600778 101351 600834 101360
rect 600688 84516 600740 84522
rect 600688 84458 600740 84464
rect 600596 84312 600648 84318
rect 600596 84254 600648 84260
rect 600792 84250 600820 101351
rect 600780 84244 600832 84250
rect 600780 84186 600832 84192
rect 600884 84182 600912 102439
rect 606404 100014 606740 100042
rect 607384 100014 607444 100042
rect 606404 95334 606432 100014
rect 607220 95600 607272 95606
rect 607220 95542 607272 95548
rect 606392 95328 606444 95334
rect 606392 95270 606444 95276
rect 605748 93900 605800 93906
rect 605748 93842 605800 93848
rect 601700 91044 601752 91050
rect 601700 90986 601752 90992
rect 600872 84176 600924 84182
rect 600872 84118 600924 84124
rect 591948 80844 592000 80850
rect 591948 80786 592000 80792
rect 596180 80844 596232 80850
rect 596180 80786 596232 80792
rect 590660 73160 590712 73166
rect 590660 73102 590712 73108
rect 590672 66298 590700 73102
rect 590660 66292 590712 66298
rect 590660 66234 590712 66240
rect 586428 66224 586480 66230
rect 586428 66166 586480 66172
rect 590660 64864 590712 64870
rect 590660 64806 590712 64812
rect 583852 58676 583904 58682
rect 583852 58618 583904 58624
rect 582564 58132 582616 58138
rect 582564 58074 582616 58080
rect 582102 55312 582158 55321
rect 582102 55247 582158 55256
rect 580906 53816 580962 53825
rect 580906 53751 580962 53760
rect 582576 53650 582604 58074
rect 590672 58002 590700 64806
rect 590752 62144 590804 62150
rect 590752 62086 590804 62092
rect 590764 58002 590792 62086
rect 591960 58138 591988 80786
rect 601712 80186 601740 90986
rect 601620 80158 601740 80186
rect 600228 78532 600280 78538
rect 600228 78474 600280 78480
rect 600044 74520 600096 74526
rect 600044 74462 600096 74468
rect 598940 69080 598992 69086
rect 598940 69022 598992 69028
rect 598952 62150 598980 69022
rect 600056 64870 600084 74462
rect 600044 64864 600096 64870
rect 600044 64806 600096 64812
rect 598940 62144 598992 62150
rect 598940 62086 598992 62092
rect 600240 60858 600268 78474
rect 601620 73166 601648 80158
rect 605760 74526 605788 93842
rect 605840 77852 605892 77858
rect 605840 77794 605892 77800
rect 605748 74520 605800 74526
rect 605748 74462 605800 74468
rect 601608 73160 601660 73166
rect 601608 73102 601660 73108
rect 605852 69086 605880 77794
rect 605840 69080 605892 69086
rect 605840 69022 605892 69028
rect 600320 63572 600372 63578
rect 600320 63514 600372 63520
rect 595076 60852 595128 60858
rect 595076 60794 595128 60800
rect 600228 60852 600280 60858
rect 600228 60794 600280 60800
rect 591948 58132 592000 58138
rect 591948 58074 592000 58080
rect 586428 57996 586480 58002
rect 586428 57938 586480 57944
rect 590660 57996 590712 58002
rect 590660 57938 590712 57944
rect 590752 57996 590804 58002
rect 590752 57938 590804 57944
rect 585140 57928 585192 57934
rect 585140 57870 585192 57876
rect 582564 53644 582616 53650
rect 582564 53586 582616 53592
rect 585152 49842 585180 57870
rect 579620 49836 579672 49842
rect 579620 49778 579672 49784
rect 585140 49836 585192 49842
rect 585140 49778 585192 49784
rect 578608 49768 578660 49774
rect 578608 49710 578660 49716
rect 578240 46980 578292 46986
rect 578240 46922 578292 46928
rect 578620 45694 578648 49710
rect 578608 45688 578660 45694
rect 578608 45630 578660 45636
rect 579632 44282 579660 49778
rect 579540 44254 579660 44282
rect 578148 44192 578200 44198
rect 578148 44134 578200 44140
rect 574836 42288 574888 42294
rect 574836 42230 574888 42236
rect 579540 42226 579568 44254
rect 586440 44130 586468 57938
rect 595088 55282 595116 60794
rect 587900 55276 587952 55282
rect 587900 55218 587952 55224
rect 595076 55276 595128 55282
rect 595076 55218 595128 55224
rect 587912 49774 587940 55218
rect 600332 51066 600360 63514
rect 587992 51060 588044 51066
rect 587992 51002 588044 51008
rect 600320 51060 600372 51066
rect 600320 51002 600372 51008
rect 587900 49768 587952 49774
rect 587900 49710 587952 49716
rect 586428 44124 586480 44130
rect 586428 44066 586480 44072
rect 579528 42220 579580 42226
rect 579528 42162 579580 42168
rect 571338 41984 571394 41993
rect 571338 41919 571394 41928
rect 563610 41712 563666 41721
rect 563610 41647 563666 41656
rect 588004 41585 588032 51002
rect 607232 43994 607260 95542
rect 607312 93832 607364 93838
rect 607312 93774 607364 93780
rect 607324 77858 607352 93774
rect 607312 77852 607364 77858
rect 607312 77794 607364 77800
rect 607416 45830 607444 100014
rect 607508 100014 608028 100042
rect 608152 100014 608672 100042
rect 608980 100014 609316 100042
rect 609960 100014 610020 100042
rect 607508 63578 607536 100014
rect 608152 91094 608180 100014
rect 608980 95606 609008 100014
rect 608968 95600 609020 95606
rect 608968 95542 609020 95548
rect 609992 91118 610020 100014
rect 610360 100014 610604 100042
rect 610728 100014 611248 100042
rect 611556 100014 611892 100042
rect 612200 100014 612536 100042
rect 612936 100014 613180 100042
rect 613580 100014 613916 100042
rect 614560 100014 614804 100042
rect 610256 95600 610308 95606
rect 610256 95542 610308 95548
rect 607600 91066 608180 91094
rect 609980 91112 610032 91118
rect 607496 63572 607548 63578
rect 607496 63514 607548 63520
rect 607404 45824 607456 45830
rect 607404 45766 607456 45772
rect 607600 45762 607628 91066
rect 609980 91054 610032 91060
rect 610268 45898 610296 95542
rect 610360 95266 610388 100014
rect 610348 95260 610400 95266
rect 610348 95202 610400 95208
rect 610728 91094 610756 100014
rect 611556 95606 611584 100014
rect 611544 95600 611596 95606
rect 611544 95542 611596 95548
rect 612200 93838 612228 100014
rect 612936 95402 612964 100014
rect 613016 95600 613068 95606
rect 613016 95542 613068 95548
rect 612924 95396 612976 95402
rect 612924 95338 612976 95344
rect 612188 93832 612240 93838
rect 612188 93774 612240 93780
rect 610360 91066 610756 91094
rect 610360 78538 610388 91066
rect 610348 78532 610400 78538
rect 610348 78474 610400 78480
rect 610256 45892 610308 45898
rect 610256 45834 610308 45840
rect 607588 45756 607640 45762
rect 607588 45698 607640 45704
rect 607220 43988 607272 43994
rect 607220 43930 607272 43936
rect 613028 43926 613056 95542
rect 613580 93906 613608 100014
rect 614776 95810 614804 100014
rect 614868 100014 615204 100042
rect 615848 100014 616184 100042
rect 616492 100014 616828 100042
rect 617136 100014 617472 100042
rect 617780 100014 618116 100042
rect 618424 100014 618760 100042
rect 619068 100014 619404 100042
rect 619712 100014 620048 100042
rect 614764 95804 614816 95810
rect 614764 95746 614816 95752
rect 614868 95606 614896 100014
rect 614856 95600 614908 95606
rect 614856 95542 614908 95548
rect 616156 95470 616184 100014
rect 616144 95464 616196 95470
rect 616144 95406 616196 95412
rect 616800 94586 616828 100014
rect 617444 94994 617472 100014
rect 617432 94988 617484 94994
rect 617432 94930 617484 94936
rect 618088 94858 618116 100014
rect 618260 95600 618312 95606
rect 618260 95542 618312 95548
rect 618076 94852 618128 94858
rect 618076 94794 618128 94800
rect 616788 94580 616840 94586
rect 616788 94522 616840 94528
rect 613568 93900 613620 93906
rect 613568 93842 613620 93848
rect 613016 43920 613068 43926
rect 613016 43862 613068 43868
rect 618272 43858 618300 95542
rect 618732 95266 618760 100014
rect 619376 95402 619404 100014
rect 620020 95674 620048 100014
rect 620112 100014 620448 100042
rect 621092 100014 621152 100042
rect 620008 95668 620060 95674
rect 620008 95610 620060 95616
rect 620112 95606 620140 100014
rect 620100 95600 620152 95606
rect 620100 95542 620152 95548
rect 619364 95396 619416 95402
rect 619364 95338 619416 95344
rect 618720 95260 618772 95266
rect 618720 95202 618772 95208
rect 618260 43852 618312 43858
rect 618260 43794 618312 43800
rect 621124 43586 621152 100014
rect 621400 100014 621736 100042
rect 621860 100014 622380 100042
rect 622688 100014 623024 100042
rect 623332 100014 623668 100042
rect 623976 100014 624312 100042
rect 624620 100014 624956 100042
rect 625600 100014 625936 100042
rect 626244 100014 626488 100042
rect 626980 100014 627316 100042
rect 627624 100014 627960 100042
rect 628268 100014 628328 100042
rect 621204 95600 621256 95606
rect 621204 95542 621256 95548
rect 621216 43790 621244 95542
rect 621296 95532 621348 95538
rect 621296 95474 621348 95480
rect 621204 43784 621256 43790
rect 621204 43726 621256 43732
rect 621308 43722 621336 95474
rect 621296 43716 621348 43722
rect 621296 43658 621348 43664
rect 621112 43580 621164 43586
rect 621112 43522 621164 43528
rect 621400 43518 621428 100014
rect 621860 91094 621888 100014
rect 622688 95606 622716 100014
rect 622676 95600 622728 95606
rect 622676 95542 622728 95548
rect 623332 95538 623360 100014
rect 623504 95668 623556 95674
rect 623504 95610 623556 95616
rect 623320 95532 623372 95538
rect 623320 95474 623372 95480
rect 623228 95464 623280 95470
rect 623228 95406 623280 95412
rect 622124 95396 622176 95402
rect 622124 95338 622176 95344
rect 621940 94852 621992 94858
rect 621940 94794 621992 94800
rect 621492 91066 621888 91094
rect 621492 43654 621520 91066
rect 621952 84153 621980 94794
rect 622136 86057 622164 95338
rect 622676 95260 622728 95266
rect 622676 95202 622728 95208
rect 622122 86048 622178 86057
rect 622122 85983 622178 85992
rect 622688 85105 622716 95202
rect 623136 94580 623188 94586
rect 623136 94522 623188 94528
rect 623148 88913 623176 94522
rect 623134 88904 623190 88913
rect 623134 88839 623190 88848
rect 623240 87961 623268 95406
rect 623320 94988 623372 94994
rect 623320 94930 623372 94936
rect 623226 87952 623282 87961
rect 623226 87887 623282 87896
rect 622674 85096 622730 85105
rect 622674 85031 622730 85040
rect 621938 84144 621994 84153
rect 621938 84079 621994 84088
rect 623332 83201 623360 94930
rect 623516 87009 623544 95610
rect 623780 95600 623832 95606
rect 623780 95542 623832 95548
rect 623792 90681 623820 95542
rect 623778 90672 623834 90681
rect 623778 90607 623834 90616
rect 623976 89729 624004 100014
rect 624620 95606 624648 100014
rect 624608 95600 624660 95606
rect 624608 95542 624660 95548
rect 625908 91633 625936 100014
rect 626460 92585 626488 100014
rect 627288 93537 627316 100014
rect 627932 94489 627960 100014
rect 628300 95985 628328 100014
rect 628760 100014 628912 100042
rect 629556 100014 629708 100042
rect 630200 100014 630628 100042
rect 630844 100014 631180 100042
rect 631488 100014 631824 100042
rect 632132 100014 632468 100042
rect 632776 100014 633112 100042
rect 633512 100014 633848 100042
rect 634156 100014 634492 100042
rect 634800 100014 635136 100042
rect 635444 100014 635780 100042
rect 636088 100014 636332 100042
rect 636732 100014 637068 100042
rect 637376 100014 637528 100042
rect 638020 100014 638356 100042
rect 638664 100014 638908 100042
rect 639308 100014 639644 100042
rect 639952 100014 640104 100042
rect 640688 100014 640932 100042
rect 641332 100014 641668 100042
rect 641976 100014 642312 100042
rect 642620 100014 642680 100042
rect 643264 100014 643600 100042
rect 643908 100014 644244 100042
rect 644552 100014 644796 100042
rect 628286 95976 628342 95985
rect 628286 95911 628342 95920
rect 628760 95826 628788 100014
rect 628728 95798 628788 95826
rect 629680 95826 629708 100014
rect 630600 95826 630628 100014
rect 631152 96082 631180 100014
rect 631140 96076 631192 96082
rect 631140 96018 631192 96024
rect 631796 95946 631824 100014
rect 632440 96082 632468 100014
rect 633084 96626 633112 100014
rect 633072 96620 633124 96626
rect 633072 96562 633124 96568
rect 633820 96558 633848 100014
rect 633808 96552 633860 96558
rect 633808 96494 633860 96500
rect 634464 96490 634492 100014
rect 634452 96484 634504 96490
rect 634452 96426 634504 96432
rect 635108 96082 635136 100014
rect 635280 96620 635332 96626
rect 635280 96562 635332 96568
rect 632106 96076 632158 96082
rect 632106 96018 632158 96024
rect 632428 96076 632480 96082
rect 632428 96018 632480 96024
rect 634406 96076 634458 96082
rect 634406 96018 634458 96024
rect 635096 96076 635148 96082
rect 635096 96018 635148 96024
rect 631784 95940 631836 95946
rect 631784 95882 631836 95888
rect 629680 95798 629832 95826
rect 630600 95798 631028 95826
rect 632118 95812 632146 96018
rect 632980 95940 633032 95946
rect 632980 95882 633032 95888
rect 632992 95826 633020 95882
rect 632992 95798 633328 95826
rect 634418 95812 634446 96018
rect 635292 95826 635320 96562
rect 635752 96422 635780 100014
rect 636304 96626 636332 100014
rect 636292 96620 636344 96626
rect 636292 96562 636344 96568
rect 637040 96558 637068 100014
rect 636384 96552 636436 96558
rect 636384 96494 636436 96500
rect 637028 96552 637080 96558
rect 637028 96494 637080 96500
rect 635740 96416 635792 96422
rect 635740 96358 635792 96364
rect 636396 95826 636424 96494
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637500 95742 637528 100014
rect 637580 96484 637632 96490
rect 637580 96426 637632 96432
rect 637592 95826 637620 96426
rect 637592 95798 637928 95826
rect 637488 95736 637540 95742
rect 637488 95678 637540 95684
rect 638328 95606 638356 100014
rect 638880 95878 638908 100014
rect 639006 96076 639058 96082
rect 639006 96018 639058 96024
rect 638868 95872 638920 95878
rect 638868 95814 638920 95820
rect 639018 95812 639046 96018
rect 639616 95810 639644 100014
rect 639880 96416 639932 96422
rect 639880 96358 639932 96364
rect 639892 95826 639920 96358
rect 640076 95946 640104 100014
rect 640064 95940 640116 95946
rect 640064 95882 640116 95888
rect 639604 95804 639656 95810
rect 639892 95798 640228 95826
rect 639604 95746 639656 95752
rect 640904 95742 640932 100014
rect 640984 96620 641036 96626
rect 640984 96562 641036 96568
rect 640996 95826 641024 96562
rect 640996 95798 641332 95826
rect 640524 95736 640576 95742
rect 640522 95704 640524 95713
rect 640892 95736 640944 95742
rect 640576 95704 640578 95713
rect 640892 95678 640944 95684
rect 641640 95674 641668 100014
rect 640522 95639 640578 95648
rect 641628 95668 641680 95674
rect 641628 95610 641680 95616
rect 642284 95606 642312 100014
rect 642364 96552 642416 96558
rect 642364 96494 642416 96500
rect 642376 95826 642404 96494
rect 642376 95798 642528 95826
rect 638316 95600 638368 95606
rect 638316 95542 638368 95548
rect 642272 95600 642324 95606
rect 642272 95542 642324 95548
rect 627918 94480 627974 94489
rect 627918 94415 627974 94424
rect 627274 93528 627330 93537
rect 627274 93463 627330 93472
rect 626446 92576 626502 92585
rect 626446 92511 626502 92520
rect 625894 91624 625950 91633
rect 625894 91559 625950 91568
rect 623962 89720 624018 89729
rect 623962 89655 624018 89664
rect 623502 87000 623558 87009
rect 623502 86935 623558 86944
rect 623318 83192 623374 83201
rect 623318 83127 623374 83136
rect 622306 82240 622362 82249
rect 622306 82175 622362 82184
rect 621480 43648 621532 43654
rect 621480 43590 621532 43596
rect 621388 43512 621440 43518
rect 621388 43454 621440 43460
rect 622320 43382 622348 82175
rect 622490 81424 622546 81433
rect 622490 81359 622546 81368
rect 622504 43450 622532 81359
rect 631856 80974 631916 81002
rect 639308 80974 639368 81002
rect 622492 43444 622544 43450
rect 622492 43386 622544 43392
rect 622308 43376 622360 43382
rect 622308 43318 622360 43324
rect 631888 43314 631916 80974
rect 639340 45558 639368 80974
rect 642652 46918 642680 100014
rect 642824 95668 642876 95674
rect 642824 95610 642876 95616
rect 642732 95532 642784 95538
rect 642732 95474 642784 95480
rect 642744 92721 642772 95474
rect 642730 92712 642786 92721
rect 642730 92647 642786 92656
rect 642640 46912 642692 46918
rect 642640 46854 642692 46860
rect 642836 45626 642864 95610
rect 642916 95600 642968 95606
rect 642916 95542 642968 95548
rect 642928 52426 642956 95542
rect 643100 94988 643152 94994
rect 643100 94930 643152 94936
rect 643112 85270 643140 94930
rect 643572 94246 643600 100014
rect 643560 94240 643612 94246
rect 643560 94182 643612 94188
rect 644216 94110 644244 100014
rect 644204 94104 644256 94110
rect 644204 94046 644256 94052
rect 644768 93906 644796 100014
rect 644860 100014 645196 100042
rect 645840 100014 646176 100042
rect 646484 100014 646820 100042
rect 647220 100014 647556 100042
rect 647864 100014 648108 100042
rect 644860 94994 644888 100014
rect 646044 95940 646096 95946
rect 646044 95882 646096 95888
rect 645952 95804 646004 95810
rect 645952 95746 646004 95752
rect 645860 95736 645912 95742
rect 645860 95678 645912 95684
rect 644848 94988 644900 94994
rect 644848 94930 644900 94936
rect 644756 93900 644808 93906
rect 644756 93842 644808 93848
rect 643100 85264 643152 85270
rect 643100 85206 643152 85212
rect 645872 82249 645900 95678
rect 645964 95010 645992 95746
rect 646056 95146 646084 95882
rect 646148 95334 646176 100014
rect 646792 95946 646820 100014
rect 647528 96082 647556 100014
rect 647516 96076 647568 96082
rect 647516 96018 647568 96024
rect 646780 95940 646832 95946
rect 646780 95882 646832 95888
rect 646228 95872 646280 95878
rect 646228 95814 646280 95820
rect 646136 95328 646188 95334
rect 646136 95270 646188 95276
rect 646056 95118 646176 95146
rect 645964 94982 646084 95010
rect 645952 94920 646004 94926
rect 645952 94862 646004 94868
rect 645964 89729 645992 94862
rect 645950 89720 646006 89729
rect 645950 89655 646006 89664
rect 646056 87145 646084 94982
rect 646042 87136 646098 87145
rect 646042 87071 646098 87080
rect 646148 84697 646176 95118
rect 646240 94926 646268 95814
rect 646412 95600 646464 95606
rect 646412 95542 646464 95548
rect 646228 94920 646280 94926
rect 646228 94862 646280 94868
rect 646424 85202 646452 95542
rect 648080 94518 648108 100014
rect 648172 100014 648508 100042
rect 649152 100014 649396 100042
rect 648172 95606 648200 100014
rect 648160 95600 648212 95606
rect 648160 95542 648212 95548
rect 648620 95396 648672 95402
rect 648620 95338 648672 95344
rect 648068 94512 648120 94518
rect 648068 94454 648120 94460
rect 648632 85338 648660 95338
rect 648712 94716 648764 94722
rect 648712 94658 648764 94664
rect 648724 85406 648752 94658
rect 648896 94580 648948 94586
rect 648896 94522 648948 94528
rect 648908 85542 648936 94522
rect 649368 94042 649396 100014
rect 649460 100014 649796 100042
rect 650104 100014 650440 100042
rect 650748 100014 651084 100042
rect 651728 100014 652064 100042
rect 652372 100014 652708 100042
rect 653016 100014 653352 100042
rect 649460 94722 649488 100014
rect 649448 94716 649500 94722
rect 649448 94658 649500 94664
rect 650104 94586 650132 100014
rect 650748 95402 650776 100014
rect 652036 96490 652064 100014
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 652680 95674 652708 100014
rect 652760 96076 652812 96082
rect 652760 96018 652812 96024
rect 652668 95668 652720 95674
rect 652668 95610 652720 95616
rect 650736 95396 650788 95402
rect 650736 95338 650788 95344
rect 651840 94852 651892 94858
rect 651840 94794 651892 94800
rect 650092 94580 650144 94586
rect 650092 94522 650144 94528
rect 649356 94036 649408 94042
rect 649356 93978 649408 93984
rect 648896 85536 648948 85542
rect 648896 85478 648948 85484
rect 651852 85474 651880 94794
rect 652772 92585 652800 96018
rect 653324 94722 653352 100014
rect 653416 100014 653752 100042
rect 654396 100014 654732 100042
rect 655040 100014 655376 100042
rect 655684 100014 656020 100042
rect 656328 100014 656664 100042
rect 656972 100014 657308 100042
rect 653416 94858 653444 100014
rect 654704 96558 654732 100014
rect 654692 96552 654744 96558
rect 654692 96494 654744 96500
rect 653404 94852 653456 94858
rect 653404 94794 653456 94800
rect 653312 94716 653364 94722
rect 653312 94658 653364 94664
rect 654048 94104 654100 94110
rect 654048 94046 654100 94052
rect 652944 93900 652996 93906
rect 652944 93842 652996 93848
rect 652758 92576 652814 92585
rect 652758 92511 652814 92520
rect 652956 90681 652984 93842
rect 654060 91497 654088 94046
rect 655348 93401 655376 100014
rect 655992 96626 656020 100014
rect 655980 96620 656032 96626
rect 655980 96562 656032 96568
rect 656636 95402 656664 100014
rect 656992 95600 657044 95606
rect 656992 95542 657044 95548
rect 656624 95396 656676 95402
rect 656624 95338 656676 95344
rect 656900 94580 656952 94586
rect 656900 94522 656952 94528
rect 656912 94042 656940 94522
rect 656900 94036 656952 94042
rect 656900 93978 656952 93984
rect 655334 93392 655390 93401
rect 655334 93327 655390 93336
rect 654046 91488 654102 91497
rect 654046 91423 654102 91432
rect 652942 90672 652998 90681
rect 652942 90607 652998 90616
rect 657004 90409 657032 95542
rect 657084 95260 657136 95266
rect 657084 95202 657136 95208
rect 656990 90400 657046 90409
rect 656990 90335 657046 90344
rect 657096 88874 657124 95202
rect 657280 94654 657308 100014
rect 657372 100014 657616 100042
rect 657924 100014 658260 100042
rect 658904 100014 659148 100042
rect 657372 94761 657400 100014
rect 657728 99816 657780 99822
rect 657728 99758 657780 99764
rect 657740 95132 657768 99758
rect 657924 95266 657952 100014
rect 659120 96558 659148 100014
rect 659212 100014 659548 100042
rect 660284 100014 660620 100042
rect 658280 96552 658332 96558
rect 658280 96494 658332 96500
rect 659108 96552 659160 96558
rect 659108 96494 659160 96500
rect 657912 95260 657964 95266
rect 657912 95202 657964 95208
rect 658292 95132 658320 96494
rect 659212 95606 659240 100014
rect 659568 96620 659620 96626
rect 659568 96562 659620 96568
rect 659200 95600 659252 95606
rect 659200 95542 659252 95548
rect 659580 95132 659608 96562
rect 660592 95538 660620 100014
rect 660914 99822 660942 100028
rect 661572 100014 661908 100042
rect 662216 100014 662276 100042
rect 662860 100014 663288 100042
rect 663504 100014 663656 100042
rect 660902 99816 660954 99822
rect 660902 99758 660954 99764
rect 661880 96626 661908 100014
rect 661868 96620 661920 96626
rect 661868 96562 661920 96568
rect 661960 96484 662012 96490
rect 661960 96426 662012 96432
rect 660580 95532 660632 95538
rect 660580 95474 660632 95480
rect 661408 95532 661460 95538
rect 661408 95474 661460 95480
rect 661420 95132 661448 95474
rect 661972 95132 662000 96426
rect 662248 95577 662276 100014
rect 663064 96620 663116 96626
rect 663064 96562 663116 96568
rect 662512 96552 662564 96558
rect 662512 96494 662564 96500
rect 662234 95568 662290 95577
rect 662234 95503 662290 95512
rect 662524 95132 662552 96494
rect 663076 95132 663104 96562
rect 663156 95396 663208 95402
rect 663156 95338 663208 95344
rect 657358 94752 657414 94761
rect 657358 94687 657414 94696
rect 657268 94648 657320 94654
rect 657268 94590 657320 94596
rect 658568 94586 658858 94602
rect 658556 94580 658858 94586
rect 658608 94574 658858 94580
rect 658556 94522 658608 94528
rect 659844 94512 659896 94518
rect 660396 94512 660448 94518
rect 659896 94460 660146 94466
rect 659844 94454 660146 94460
rect 660448 94460 660698 94466
rect 660396 94454 660698 94460
rect 659856 94438 660146 94454
rect 660408 94438 660698 94454
rect 663168 91066 663196 95338
rect 663260 93809 663288 100014
rect 663340 95940 663392 95946
rect 663340 95882 663392 95888
rect 663246 93800 663302 93809
rect 663246 93735 663302 93744
rect 663352 93129 663380 95882
rect 663432 95328 663484 95334
rect 663432 95270 663484 95276
rect 663338 93120 663394 93129
rect 663338 93055 663394 93064
rect 663444 92313 663472 95270
rect 663524 94648 663576 94654
rect 663524 94590 663576 94596
rect 663430 92304 663486 92313
rect 663430 92239 663486 92248
rect 663536 91094 663564 94590
rect 663246 91080 663302 91089
rect 663168 91038 663246 91066
rect 663246 91015 663302 91024
rect 663444 91066 663564 91094
rect 663444 89593 663472 91066
rect 663430 89584 663486 89593
rect 663430 89519 663486 89528
rect 658016 88874 658306 88890
rect 659488 88874 659594 88890
rect 663628 88874 663656 100014
rect 663800 95668 663852 95674
rect 663800 95610 663852 95616
rect 663708 94716 663760 94722
rect 663708 94658 663760 94664
rect 663720 90409 663748 94658
rect 663706 90400 663762 90409
rect 663706 90335 663762 90344
rect 657084 88868 657136 88874
rect 657084 88810 657136 88816
rect 658004 88868 658306 88874
rect 658056 88862 658306 88868
rect 659476 88868 659594 88874
rect 658004 88810 658056 88816
rect 659528 88862 659594 88868
rect 663616 88868 663668 88874
rect 659476 88810 659528 88816
rect 663616 88810 663668 88816
rect 662142 88768 662198 88777
rect 661986 88726 662142 88754
rect 663812 88754 663840 95610
rect 665180 95192 665232 95198
rect 665180 95134 665232 95140
rect 662538 88726 663840 88754
rect 662142 88703 662198 88712
rect 651840 85468 651892 85474
rect 651840 85410 651892 85416
rect 648712 85400 648764 85406
rect 648712 85342 648764 85348
rect 657188 85338 657216 88196
rect 657740 85542 657768 88196
rect 657728 85536 657780 85542
rect 657728 85478 657780 85484
rect 658844 85474 658872 88196
rect 658832 85468 658884 85474
rect 658832 85410 658884 85416
rect 648620 85332 648672 85338
rect 648620 85274 648672 85280
rect 657176 85332 657228 85338
rect 657176 85274 657228 85280
rect 660132 85270 660160 88196
rect 660684 85406 660712 88196
rect 660672 85400 660724 85406
rect 660672 85342 660724 85348
rect 660120 85264 660172 85270
rect 660120 85206 660172 85212
rect 661420 85202 661448 88196
rect 646412 85196 646464 85202
rect 646412 85138 646464 85144
rect 661408 85196 661460 85202
rect 661408 85138 661460 85144
rect 646134 84688 646190 84697
rect 646134 84623 646190 84632
rect 645858 82240 645914 82249
rect 645858 82175 645914 82184
rect 642916 52420 642968 52426
rect 642916 52362 642968 52368
rect 661130 47560 661186 47569
rect 661130 47495 661186 47504
rect 661144 46249 661172 47495
rect 665192 47433 665220 95134
rect 666572 48521 666600 989402
rect 666836 987896 666888 987902
rect 666836 987838 666888 987844
rect 666652 987760 666704 987766
rect 666652 987702 666704 987708
rect 666664 183938 666692 987702
rect 666744 984836 666796 984842
rect 666744 984778 666796 984784
rect 666652 183932 666704 183938
rect 666652 183874 666704 183880
rect 666650 183832 666706 183841
rect 666650 183767 666706 183776
rect 666664 180441 666692 183767
rect 666650 180432 666706 180441
rect 666650 180367 666706 180376
rect 666650 178800 666706 178809
rect 666650 178735 666706 178744
rect 666664 175409 666692 178735
rect 666756 176662 666784 984778
rect 666848 179382 666876 987838
rect 669228 987828 669280 987834
rect 669228 987770 669280 987776
rect 669134 985688 669190 985697
rect 669134 985623 669190 985632
rect 668952 983136 669004 983142
rect 668952 983078 669004 983084
rect 669042 983104 669098 983113
rect 668584 983000 668636 983006
rect 668584 982942 668636 982948
rect 668492 982932 668544 982938
rect 668492 982874 668544 982880
rect 668400 756424 668452 756430
rect 668400 756366 668452 756372
rect 668412 713726 668440 756366
rect 668400 713720 668452 713726
rect 668400 713662 668452 713668
rect 666928 709776 666980 709782
rect 666928 709718 666980 709724
rect 666940 580106 666968 709718
rect 668504 621042 668532 982874
rect 668596 623830 668624 982942
rect 668768 841968 668820 841974
rect 668768 841910 668820 841916
rect 668676 749012 668728 749018
rect 668676 748954 668728 748960
rect 668688 624034 668716 748954
rect 668780 715766 668808 841910
rect 668860 762816 668912 762822
rect 668860 762758 668912 762764
rect 668768 715760 668820 715766
rect 668768 715702 668820 715708
rect 668768 712836 668820 712842
rect 668768 712778 668820 712784
rect 668676 624028 668728 624034
rect 668676 623970 668728 623976
rect 668584 623824 668636 623830
rect 668584 623766 668636 623772
rect 668492 621036 668544 621042
rect 668492 620978 668544 620984
rect 666928 580100 666980 580106
rect 666928 580042 666980 580048
rect 667020 457496 667072 457502
rect 667020 457438 667072 457444
rect 666928 336796 666980 336802
rect 666928 336738 666980 336744
rect 666836 179376 666888 179382
rect 666836 179318 666888 179324
rect 666940 176866 666968 336738
rect 667032 313750 667060 457438
rect 667020 313744 667072 313750
rect 667020 313686 667072 313692
rect 668780 278322 668808 712778
rect 668872 624170 668900 762758
rect 668964 713250 668992 983078
rect 669042 983039 669098 983048
rect 668952 713244 669004 713250
rect 668952 713186 669004 713192
rect 669056 712434 669084 983039
rect 669044 712428 669096 712434
rect 669044 712370 669096 712376
rect 669056 667758 669084 712370
rect 669148 669798 669176 985623
rect 669136 669792 669188 669798
rect 669136 669734 669188 669740
rect 669044 667752 669096 667758
rect 669044 667694 669096 667700
rect 669044 629332 669096 629338
rect 669044 629274 669096 629280
rect 668860 624164 668912 624170
rect 668860 624106 668912 624112
rect 669056 532914 669084 629274
rect 669136 590708 669188 590714
rect 669136 590650 669188 590656
rect 669044 532908 669096 532914
rect 669044 532850 669096 532856
rect 669148 491706 669176 590650
rect 669136 491700 669188 491706
rect 669136 491642 669188 491648
rect 669136 483064 669188 483070
rect 669136 483006 669188 483012
rect 669044 364472 669096 364478
rect 669044 364414 669096 364420
rect 668768 278316 668820 278322
rect 668768 278258 668820 278264
rect 669056 221066 669084 364414
rect 669148 356386 669176 483006
rect 669136 356380 669188 356386
rect 669136 356322 669188 356328
rect 669136 323944 669188 323950
rect 669136 323886 669188 323892
rect 669044 221060 669096 221066
rect 669044 221002 669096 221008
rect 667020 183932 667072 183938
rect 667020 183874 667072 183880
rect 666928 176860 666980 176866
rect 666928 176802 666980 176808
rect 666744 176656 666796 176662
rect 666744 176598 666796 176604
rect 667032 176594 667060 183874
rect 669148 177002 669176 323886
rect 669136 176996 669188 177002
rect 669136 176938 669188 176944
rect 667020 176588 667072 176594
rect 667020 176530 667072 176536
rect 666650 175400 666706 175409
rect 666650 175335 666706 175344
rect 666650 173632 666706 173641
rect 666650 173567 666706 173576
rect 666664 170241 666692 173567
rect 666650 170232 666706 170241
rect 666650 170167 666706 170176
rect 666650 168600 666706 168609
rect 666650 168535 666706 168544
rect 666664 165209 666692 168535
rect 666650 165200 666706 165209
rect 666650 165135 666706 165144
rect 666650 163568 666706 163577
rect 666650 163503 666706 163512
rect 666664 160177 666692 163503
rect 666650 160168 666706 160177
rect 666650 160103 666706 160112
rect 666650 158400 666706 158409
rect 666650 158335 666706 158344
rect 666664 155009 666692 158335
rect 666650 155000 666706 155009
rect 666650 154935 666706 154944
rect 666650 153368 666706 153377
rect 666650 153303 666706 153312
rect 666664 149977 666692 153303
rect 666650 149968 666706 149977
rect 666650 149903 666706 149912
rect 666650 148200 666706 148209
rect 666650 148135 666706 148144
rect 666664 144945 666692 148135
rect 666650 144936 666706 144945
rect 666650 144871 666706 144880
rect 666650 143168 666706 143177
rect 666650 143103 666706 143112
rect 666664 139777 666692 143103
rect 666650 139768 666706 139777
rect 666650 139703 666706 139712
rect 666650 132968 666706 132977
rect 666650 132903 666706 132912
rect 666664 129577 666692 132903
rect 669240 129810 669268 987770
rect 669320 987692 669372 987698
rect 669320 987634 669372 987640
rect 669332 129878 669360 987634
rect 669596 986876 669648 986882
rect 669596 986818 669648 986824
rect 669412 986808 669464 986814
rect 669412 986750 669464 986756
rect 669424 353394 669452 986750
rect 669504 986740 669556 986746
rect 669504 986682 669556 986688
rect 669516 353530 669544 986682
rect 669608 356114 669636 986818
rect 670422 985552 670478 985561
rect 670422 985487 670478 985496
rect 675668 985516 675720 985522
rect 669688 985448 669740 985454
rect 669688 985390 669740 985396
rect 669700 488578 669728 985390
rect 670056 985380 670108 985386
rect 670056 985322 670108 985328
rect 669872 922276 669924 922282
rect 669872 922218 669924 922224
rect 669884 759626 669912 922218
rect 669872 759620 669924 759626
rect 669872 759562 669924 759568
rect 669778 759112 669834 759121
rect 669778 759047 669834 759056
rect 669688 488572 669740 488578
rect 669688 488514 669740 488520
rect 669688 485852 669740 485858
rect 669688 485794 669740 485800
rect 669596 356108 669648 356114
rect 669596 356050 669648 356056
rect 669504 353524 669556 353530
rect 669504 353466 669556 353472
rect 669412 353388 669464 353394
rect 669412 353330 669464 353336
rect 669504 350600 669556 350606
rect 669504 350542 669556 350548
rect 669412 311296 669464 311302
rect 669412 311238 669464 311244
rect 669424 132666 669452 311238
rect 669516 177138 669544 350542
rect 669596 298308 669648 298314
rect 669596 298250 669648 298256
rect 669504 177132 669556 177138
rect 669504 177074 669556 177080
rect 669608 132802 669636 298250
rect 669700 278186 669728 485794
rect 669688 278180 669740 278186
rect 669688 278122 669740 278128
rect 669792 278118 669820 759047
rect 669964 756356 670016 756362
rect 669964 756298 670016 756304
rect 669872 756288 669924 756294
rect 669872 756230 669924 756236
rect 669780 278112 669832 278118
rect 669780 278054 669832 278060
rect 669884 278050 669912 756230
rect 669872 278044 669924 278050
rect 669872 277986 669924 277992
rect 669976 277982 670004 756298
rect 670068 532846 670096 985322
rect 670240 983068 670292 983074
rect 670240 983010 670292 983016
rect 670148 935740 670200 935746
rect 670148 935682 670200 935688
rect 670160 756362 670188 935682
rect 670148 756356 670200 756362
rect 670148 756298 670200 756304
rect 670148 714944 670200 714950
rect 670148 714886 670200 714892
rect 670056 532840 670108 532846
rect 670056 532782 670108 532788
rect 670056 378208 670108 378214
rect 670056 378150 670108 378156
rect 669964 277976 670016 277982
rect 669964 277918 670016 277924
rect 670068 221202 670096 378150
rect 670160 278390 670188 714886
rect 670252 714882 670280 983010
rect 670332 935808 670384 935814
rect 670332 935750 670384 935756
rect 670344 756294 670372 935750
rect 670332 756288 670384 756294
rect 670332 756230 670384 756236
rect 670240 714876 670292 714882
rect 670240 714818 670292 714824
rect 670252 670342 670280 714818
rect 670332 713720 670384 713726
rect 670332 713662 670384 713668
rect 670240 670336 670292 670342
rect 670240 670278 670292 670284
rect 670240 621104 670292 621110
rect 670240 621046 670292 621052
rect 670252 278526 670280 621046
rect 670240 278520 670292 278526
rect 670240 278462 670292 278468
rect 670148 278384 670200 278390
rect 670148 278326 670200 278332
rect 670344 278254 670372 713662
rect 670436 621625 670464 985487
rect 675668 985458 675720 985464
rect 672538 985416 672594 985425
rect 672538 985351 672594 985360
rect 670976 985108 671028 985114
rect 670976 985050 671028 985056
rect 670884 984904 670936 984910
rect 670884 984846 670936 984852
rect 670792 984564 670844 984570
rect 670792 984506 670844 984512
rect 670700 984360 670752 984366
rect 670700 984302 670752 984308
rect 670516 759076 670568 759082
rect 670516 759018 670568 759024
rect 670528 715358 670556 759018
rect 670608 756492 670660 756498
rect 670608 756434 670660 756440
rect 670516 715352 670568 715358
rect 670516 715294 670568 715300
rect 670528 714950 670556 715294
rect 670516 714944 670568 714950
rect 670516 714886 670568 714892
rect 670516 713244 670568 713250
rect 670516 713186 670568 713192
rect 670528 668710 670556 713186
rect 670620 712842 670648 756434
rect 670608 712836 670660 712842
rect 670608 712778 670660 712784
rect 670516 668704 670568 668710
rect 670516 668646 670568 668652
rect 670608 623824 670660 623830
rect 670608 623766 670660 623772
rect 670422 621616 670478 621625
rect 670422 621551 670478 621560
rect 670516 621036 670568 621042
rect 670516 620978 670568 620984
rect 670422 619576 670478 619585
rect 670422 619511 670478 619520
rect 670436 278458 670464 619511
rect 670528 576978 670556 620978
rect 670620 580242 670648 623766
rect 670608 580236 670660 580242
rect 670608 580178 670660 580184
rect 670516 576972 670568 576978
rect 670516 576914 670568 576920
rect 670516 510876 670568 510882
rect 670516 510818 670568 510824
rect 670528 356522 670556 510818
rect 670516 356516 670568 356522
rect 670516 356458 670568 356464
rect 670516 284776 670568 284782
rect 670516 284718 670568 284724
rect 670424 278452 670476 278458
rect 670424 278394 670476 278400
rect 670332 278248 670384 278254
rect 670332 278190 670384 278196
rect 670056 221196 670108 221202
rect 670056 221138 670108 221144
rect 670528 132938 670556 284718
rect 670712 189009 670740 984302
rect 670804 194041 670832 984506
rect 670896 199073 670924 984846
rect 670988 204241 671016 985050
rect 671988 984768 672040 984774
rect 671988 984710 672040 984716
rect 671068 984700 671120 984706
rect 671068 984642 671120 984648
rect 671080 209273 671108 984642
rect 671804 705152 671856 705158
rect 671804 705094 671856 705100
rect 671160 314628 671212 314634
rect 671160 314570 671212 314576
rect 671172 312118 671200 314570
rect 671160 312112 671212 312118
rect 671160 312054 671212 312060
rect 671160 311840 671212 311846
rect 671160 311782 671212 311788
rect 671172 309670 671200 311782
rect 671160 309664 671212 309670
rect 671160 309606 671212 309612
rect 671160 218068 671212 218074
rect 671160 218010 671212 218016
rect 671066 209264 671122 209273
rect 671066 209199 671122 209208
rect 671080 205873 671108 209199
rect 671066 205864 671122 205873
rect 671066 205799 671122 205808
rect 670974 204232 671030 204241
rect 670974 204167 671030 204176
rect 670988 200841 671016 204167
rect 670974 200832 671030 200841
rect 670974 200767 671030 200776
rect 670882 199064 670938 199073
rect 670882 198999 670938 199008
rect 670896 195673 670924 198999
rect 670882 195664 670938 195673
rect 670882 195599 670938 195608
rect 670790 194032 670846 194041
rect 670790 193967 670846 193976
rect 670804 190641 670832 193967
rect 670790 190632 670846 190641
rect 670790 190567 670846 190576
rect 670698 189000 670754 189009
rect 670698 188935 670754 188944
rect 670712 185609 670740 188935
rect 670698 185600 670754 185609
rect 670698 185535 670754 185544
rect 670698 138136 670754 138145
rect 670698 138071 670754 138080
rect 670712 134745 670740 138071
rect 670698 134736 670754 134745
rect 670698 134671 670754 134680
rect 670516 132932 670568 132938
rect 670516 132874 670568 132880
rect 669596 132796 669648 132802
rect 669596 132738 669648 132744
rect 669412 132660 669464 132666
rect 669412 132602 669464 132608
rect 670792 131708 670844 131714
rect 670792 131650 670844 131656
rect 670804 129878 670832 131650
rect 670884 130076 670936 130082
rect 670884 130018 670936 130024
rect 669320 129872 669372 129878
rect 669320 129814 669372 129820
rect 670792 129872 670844 129878
rect 670792 129814 670844 129820
rect 669228 129804 669280 129810
rect 669228 129746 669280 129752
rect 666650 129568 666706 129577
rect 666650 129503 666706 129512
rect 666650 127936 666706 127945
rect 666650 127871 666706 127880
rect 666664 124545 666692 127871
rect 666650 124536 666706 124545
rect 666650 124471 666706 124480
rect 666650 122904 666706 122913
rect 666650 122839 666706 122848
rect 666664 119513 666692 122839
rect 666650 119504 666706 119513
rect 666650 119439 666706 119448
rect 670804 104145 670832 129814
rect 670896 129810 670924 130018
rect 670884 129804 670936 129810
rect 670884 129746 670936 129752
rect 670790 104136 670846 104145
rect 670790 104071 670846 104080
rect 670896 100881 670924 129746
rect 671172 107545 671200 218010
rect 671436 179376 671488 179382
rect 671436 179318 671488 179324
rect 671448 176934 671476 179318
rect 671436 176928 671488 176934
rect 671436 176870 671488 176876
rect 671344 176656 671396 176662
rect 671344 176598 671396 176604
rect 671356 175302 671384 176598
rect 671344 175296 671396 175302
rect 671344 175238 671396 175244
rect 671816 173641 671844 705094
rect 671896 309664 671948 309670
rect 671896 309606 671948 309612
rect 671908 264994 671936 309606
rect 671896 264988 671948 264994
rect 671896 264930 671948 264936
rect 671896 174480 671948 174486
rect 671896 174422 671948 174428
rect 671802 173632 671858 173641
rect 671802 173567 671858 173576
rect 671908 129742 671936 174422
rect 671896 129736 671948 129742
rect 671896 129678 671948 129684
rect 672000 129470 672028 984710
rect 672080 927444 672132 927450
rect 672080 927386 672132 927392
rect 672092 183841 672120 927386
rect 672172 749828 672224 749834
rect 672172 749770 672224 749776
rect 672078 183832 672134 183841
rect 672078 183767 672134 183776
rect 672184 178809 672212 749770
rect 672356 659728 672408 659734
rect 672356 659670 672408 659676
rect 672264 312112 672316 312118
rect 672264 312054 672316 312060
rect 672276 267510 672304 312054
rect 672264 267504 672316 267510
rect 672264 267446 672316 267452
rect 672170 178800 672226 178809
rect 672170 178735 672226 178744
rect 672172 176588 672224 176594
rect 672172 176530 672224 176536
rect 672184 174486 672212 176530
rect 672264 175296 672316 175302
rect 672264 175238 672316 175244
rect 672172 174480 672224 174486
rect 672172 174422 672224 174428
rect 672172 168292 672224 168298
rect 672172 168234 672224 168240
rect 672080 167068 672132 167074
rect 672080 167010 672132 167016
rect 671988 129464 672040 129470
rect 671988 129406 672040 129412
rect 671620 122732 671672 122738
rect 671620 122674 671672 122680
rect 671632 110945 671660 122674
rect 671618 110936 671674 110945
rect 671618 110871 671674 110880
rect 671158 107536 671214 107545
rect 671158 107471 671214 107480
rect 672000 102513 672028 129406
rect 672092 114345 672120 167010
rect 672184 117745 672212 168234
rect 672276 130694 672304 175238
rect 672368 168609 672396 659670
rect 672448 614644 672500 614650
rect 672448 614586 672500 614592
rect 672354 168600 672410 168609
rect 672354 168535 672410 168544
rect 672356 167884 672408 167890
rect 672356 167826 672408 167832
rect 672264 130688 672316 130694
rect 672264 130630 672316 130636
rect 672264 121916 672316 121922
rect 672264 121858 672316 121864
rect 672170 117736 672226 117745
rect 672170 117671 672226 117680
rect 672078 114336 672134 114345
rect 672078 114271 672134 114280
rect 672276 109313 672304 121858
rect 672368 116113 672396 167826
rect 672460 163577 672488 614586
rect 672552 579290 672580 985351
rect 672630 982968 672686 982977
rect 672630 982903 672686 982912
rect 672540 579284 672592 579290
rect 672540 579226 672592 579232
rect 672644 577658 672672 982903
rect 675680 970154 675708 985458
rect 674840 970148 674892 970154
rect 674840 970090 674892 970096
rect 675668 970148 675720 970154
rect 675668 970090 675720 970096
rect 673552 966408 673604 966414
rect 673552 966350 673604 966356
rect 673460 965048 673512 965054
rect 673460 964990 673512 964996
rect 673472 950638 673500 964990
rect 673460 950632 673512 950638
rect 673460 950574 673512 950580
rect 673564 935406 673592 966350
rect 674748 965592 674800 965598
rect 674748 965534 674800 965540
rect 673644 963348 673696 963354
rect 673644 963290 673696 963296
rect 673656 950722 673684 963290
rect 673920 962736 673972 962742
rect 673920 962678 673972 962684
rect 673828 962056 673880 962062
rect 673828 961998 673880 962004
rect 673736 961376 673788 961382
rect 673736 961318 673788 961324
rect 673748 950858 673776 961318
rect 673840 950994 673868 961998
rect 673932 960494 673960 962678
rect 673932 960466 674052 960494
rect 673920 954032 673972 954038
rect 673920 953974 673972 953980
rect 673932 951114 673960 953974
rect 673920 951108 673972 951114
rect 673920 951050 673972 951056
rect 673840 950966 673960 950994
rect 673748 950830 673868 950858
rect 673656 950694 673776 950722
rect 673644 950632 673696 950638
rect 673644 950574 673696 950580
rect 673656 935474 673684 950574
rect 673644 935468 673696 935474
rect 673644 935410 673696 935416
rect 673552 935400 673604 935406
rect 673552 935342 673604 935348
rect 673748 935338 673776 950694
rect 673736 935332 673788 935338
rect 673736 935274 673788 935280
rect 673840 932754 673868 950830
rect 673828 932748 673880 932754
rect 673828 932690 673880 932696
rect 673932 932686 673960 950966
rect 674024 932822 674052 960466
rect 674472 958860 674524 958866
rect 674472 958802 674524 958808
rect 674288 958384 674340 958390
rect 674288 958326 674340 958332
rect 674012 932816 674064 932822
rect 674012 932758 674064 932764
rect 673920 932680 673972 932686
rect 673920 932622 673972 932628
rect 674300 932278 674328 958326
rect 674380 957772 674432 957778
rect 674380 957714 674432 957720
rect 674288 932272 674340 932278
rect 674288 932214 674340 932220
rect 674392 931734 674420 957714
rect 674484 935542 674512 958802
rect 674564 957024 674616 957030
rect 674564 956966 674616 956972
rect 674472 935536 674524 935542
rect 674472 935478 674524 935484
rect 674380 931728 674432 931734
rect 674380 931670 674432 931676
rect 674576 931326 674604 956966
rect 674656 955732 674708 955738
rect 674656 955674 674708 955680
rect 674668 932890 674696 955674
rect 674760 954038 674788 965534
rect 674748 954032 674800 954038
rect 674748 953974 674800 953980
rect 674748 953896 674800 953902
rect 674748 953838 674800 953844
rect 674760 935610 674788 953838
rect 674852 952202 674880 970090
rect 675404 966414 675432 966723
rect 675392 966408 675444 966414
rect 675392 966350 675444 966356
rect 675404 965598 675432 966076
rect 675392 965592 675444 965598
rect 675392 965534 675444 965540
rect 675496 965054 675524 965435
rect 675484 965048 675536 965054
rect 675484 964990 675536 964996
rect 675404 963354 675432 963595
rect 675392 963348 675444 963354
rect 675392 963290 675444 963296
rect 675496 962742 675524 963016
rect 675484 962736 675536 962742
rect 675484 962678 675536 962684
rect 675404 962062 675432 962404
rect 675392 962056 675444 962062
rect 675392 961998 675444 962004
rect 675404 961382 675432 961755
rect 675392 961376 675444 961382
rect 675392 961318 675444 961324
rect 675024 960560 675076 960566
rect 675024 960502 675076 960508
rect 675036 955534 675064 960502
rect 675404 958866 675432 959276
rect 675392 958860 675444 958866
rect 675392 958802 675444 958808
rect 675404 958390 675432 958732
rect 675392 958384 675444 958390
rect 675392 958326 675444 958332
rect 675496 957778 675524 958052
rect 675484 957772 675536 957778
rect 675484 957714 675536 957720
rect 675404 957030 675432 957440
rect 675392 957024 675444 957030
rect 675392 956966 675444 956972
rect 675496 955738 675524 956216
rect 675484 955732 675536 955738
rect 675484 955674 675536 955680
rect 675024 955528 675076 955534
rect 675024 955470 675076 955476
rect 675484 955528 675536 955534
rect 675484 955470 675536 955476
rect 675496 955060 675524 955470
rect 675404 953902 675432 954380
rect 675392 953896 675444 953902
rect 675392 953838 675444 953844
rect 674840 952196 674892 952202
rect 674840 952138 674892 952144
rect 675404 952066 675432 952544
rect 674840 952060 674892 952066
rect 674840 952002 674892 952008
rect 675392 952060 675444 952066
rect 675392 952002 675444 952008
rect 674748 935604 674800 935610
rect 674748 935546 674800 935552
rect 674852 934998 674880 952002
rect 675668 951788 675720 951794
rect 675668 951730 675720 951736
rect 675680 938777 675708 951730
rect 675760 951108 675812 951114
rect 675760 951050 675812 951056
rect 675666 938768 675722 938777
rect 675666 938703 675722 938712
rect 674840 934992 674892 934998
rect 674840 934934 674892 934940
rect 675772 933065 675800 951050
rect 676310 939720 676366 939729
rect 676310 939655 676366 939664
rect 676126 939312 676182 939321
rect 676126 939247 676182 939256
rect 676140 938602 676168 939247
rect 676218 938904 676274 938913
rect 676218 938839 676220 938848
rect 676272 938839 676274 938848
rect 676220 938810 676272 938816
rect 676324 938738 676352 939655
rect 676312 938732 676364 938738
rect 676312 938674 676364 938680
rect 676128 938596 676180 938602
rect 676128 938538 676180 938544
rect 678978 937680 679034 937689
rect 678978 937615 679034 937624
rect 676218 936456 676274 936465
rect 676218 936391 676274 936400
rect 676034 935912 676090 935921
rect 676034 935847 676090 935856
rect 676048 935746 676076 935847
rect 676232 935814 676260 936391
rect 676220 935808 676272 935814
rect 676220 935750 676272 935756
rect 676036 935740 676088 935746
rect 676036 935682 676088 935688
rect 678992 935678 679020 937615
rect 678980 935672 679032 935678
rect 678980 935614 679032 935620
rect 676036 935604 676088 935610
rect 676036 935546 676088 935552
rect 675942 935504 675998 935513
rect 675942 935439 675944 935448
rect 675996 935439 675998 935448
rect 675944 935410 675996 935416
rect 675852 935400 675904 935406
rect 675852 935342 675904 935348
rect 675864 934697 675892 935342
rect 675944 935332 675996 935338
rect 675944 935274 675996 935280
rect 675850 934688 675906 934697
rect 675850 934623 675906 934632
rect 675956 934289 675984 935274
rect 676048 935105 676076 935546
rect 676128 935536 676180 935542
rect 676128 935478 676180 935484
rect 676034 935096 676090 935105
rect 676034 935031 676090 935040
rect 676036 934992 676088 934998
rect 676036 934934 676088 934940
rect 675942 934280 675998 934289
rect 675942 934215 675998 934224
rect 676048 933473 676076 934934
rect 676140 934017 676168 935478
rect 676126 934008 676182 934017
rect 676126 933943 676182 933952
rect 676034 933464 676090 933473
rect 676034 933399 676090 933408
rect 675758 933056 675814 933065
rect 675758 932991 675814 933000
rect 674656 932884 674708 932890
rect 674656 932826 674708 932832
rect 676036 932884 676088 932890
rect 676036 932826 676088 932832
rect 675944 932748 675996 932754
rect 675944 932690 675996 932696
rect 674564 931320 674616 931326
rect 674564 931262 674616 931268
rect 675956 931025 675984 932690
rect 676048 931841 676076 932826
rect 676128 932816 676180 932822
rect 676126 932784 676128 932793
rect 676180 932784 676182 932793
rect 676126 932719 676182 932728
rect 676128 932680 676180 932686
rect 676128 932622 676180 932628
rect 676140 932385 676168 932622
rect 676126 932376 676182 932385
rect 676126 932311 676182 932320
rect 676128 932272 676180 932278
rect 676128 932214 676180 932220
rect 676034 931832 676090 931841
rect 676034 931767 676090 931776
rect 676036 931728 676088 931734
rect 676036 931670 676088 931676
rect 676048 931433 676076 931670
rect 676034 931424 676090 931433
rect 676034 931359 676090 931368
rect 676036 931320 676088 931326
rect 676036 931262 676088 931268
rect 675942 931016 675998 931025
rect 675942 930951 675998 930960
rect 676048 930209 676076 931262
rect 676140 930753 676168 932214
rect 676126 930744 676182 930753
rect 676126 930679 676182 930688
rect 676034 930200 676090 930209
rect 676034 930135 676090 930144
rect 678978 929520 679034 929529
rect 678978 929455 679034 929464
rect 678992 928713 679020 929455
rect 678978 928704 679034 928713
rect 678978 928639 679034 928648
rect 678992 927450 679020 928639
rect 678980 927444 679032 927450
rect 678980 927386 679032 927392
rect 675772 877305 675800 877540
rect 675758 877296 675814 877305
rect 675758 877231 675814 877240
rect 675680 876625 675708 876860
rect 675666 876616 675722 876625
rect 675666 876551 675722 876560
rect 675496 875945 675524 876248
rect 675482 875936 675538 875945
rect 675482 875871 675538 875880
rect 675404 874041 675432 874412
rect 675390 874032 675446 874041
rect 675390 873967 675446 873976
rect 675404 873526 675432 873868
rect 674656 873520 674708 873526
rect 674656 873462 674708 873468
rect 675392 873520 675444 873526
rect 675392 873462 675444 873468
rect 673644 869848 673696 869854
rect 673644 869790 673696 869796
rect 673460 784984 673512 784990
rect 673460 784926 673512 784932
rect 673472 770234 673500 784926
rect 673552 782944 673604 782950
rect 673552 782886 673604 782892
rect 673564 770302 673592 782886
rect 673552 770296 673604 770302
rect 673552 770238 673604 770244
rect 673460 770228 673512 770234
rect 673460 770170 673512 770176
rect 673550 760336 673606 760345
rect 673550 760271 673606 760280
rect 673368 759144 673420 759150
rect 673564 759121 673592 760271
rect 673368 759086 673420 759092
rect 673550 759112 673606 759121
rect 673380 723178 673408 759086
rect 673550 759047 673606 759056
rect 673656 756158 673684 869790
rect 674196 869032 674248 869038
rect 674196 868974 674248 868980
rect 673736 868556 673788 868562
rect 673736 868498 673788 868504
rect 673644 756152 673696 756158
rect 673644 756094 673696 756100
rect 673748 753302 673776 868498
rect 673828 866516 673880 866522
rect 673828 866458 673880 866464
rect 673840 753506 673868 866458
rect 674012 864680 674064 864686
rect 674012 864622 674064 864628
rect 673920 862844 673972 862850
rect 673920 862786 673972 862792
rect 673932 756226 673960 862786
rect 674024 759014 674052 864622
rect 674208 792033 674236 868974
rect 674288 867808 674340 867814
rect 674288 867750 674340 867756
rect 674300 797745 674328 867750
rect 674668 854282 674696 873462
rect 675404 872710 675432 873188
rect 674748 872704 674800 872710
rect 674748 872646 674800 872652
rect 675392 872704 675444 872710
rect 675392 872646 675444 872652
rect 674656 854276 674708 854282
rect 674656 854218 674708 854224
rect 674760 854214 674788 872646
rect 675772 872273 675800 872576
rect 675758 872264 675814 872273
rect 675758 872199 675814 872208
rect 674932 870800 674984 870806
rect 674932 870742 674984 870748
rect 674944 866318 674972 870742
rect 675404 869854 675432 870060
rect 675392 869848 675444 869854
rect 675392 869790 675444 869796
rect 675404 869038 675432 869516
rect 675392 869032 675444 869038
rect 675392 868974 675444 868980
rect 675404 868562 675432 868875
rect 675392 868556 675444 868562
rect 675392 868498 675444 868504
rect 675404 867814 675432 868224
rect 675392 867808 675444 867814
rect 675392 867750 675444 867756
rect 675404 866522 675432 867035
rect 675392 866516 675444 866522
rect 675392 866458 675444 866464
rect 674932 866312 674984 866318
rect 674932 866254 674984 866260
rect 675392 866312 675444 866318
rect 675392 866254 675444 866260
rect 675404 865844 675432 866254
rect 675404 864686 675432 865195
rect 675392 864680 675444 864686
rect 675392 864622 675444 864628
rect 675496 862850 675524 863328
rect 675484 862844 675536 862850
rect 675484 862786 675536 862792
rect 675576 854276 675628 854282
rect 675576 854218 675628 854224
rect 674748 854208 674800 854214
rect 674748 854150 674800 854156
rect 674286 797736 674342 797745
rect 674286 797671 674342 797680
rect 674748 796340 674800 796346
rect 674748 796282 674800 796288
rect 674564 796272 674616 796278
rect 674564 796214 674616 796220
rect 674194 792024 674250 792033
rect 674194 791959 674250 791968
rect 674288 780632 674340 780638
rect 674288 780574 674340 780580
rect 674196 779340 674248 779346
rect 674196 779282 674248 779288
rect 674208 770386 674236 779282
rect 674300 770574 674328 780574
rect 674472 779816 674524 779822
rect 674472 779758 674524 779764
rect 674380 778796 674432 778802
rect 674380 778738 674432 778744
rect 674392 777481 674420 778738
rect 674378 777472 674434 777481
rect 674378 777407 674434 777416
rect 674380 777368 674432 777374
rect 674380 777310 674432 777316
rect 674288 770568 674340 770574
rect 674288 770510 674340 770516
rect 674392 770522 674420 777310
rect 674484 773430 674512 779758
rect 674576 776914 674604 796214
rect 674656 782468 674708 782474
rect 674656 782410 674708 782416
rect 674668 777102 674696 782410
rect 674760 778802 674788 796282
rect 675588 796278 675616 854218
rect 675760 854208 675812 854214
rect 675760 854150 675812 854156
rect 675772 796346 675800 854150
rect 675760 796340 675812 796346
rect 675760 796282 675812 796288
rect 675576 796272 675628 796278
rect 675576 796214 675628 796220
rect 675404 787817 675432 788324
rect 675390 787808 675446 787817
rect 675390 787743 675446 787752
rect 675404 787273 675432 787679
rect 675390 787264 675446 787273
rect 675390 787199 675446 787208
rect 675404 786865 675432 787032
rect 675390 786856 675446 786865
rect 675390 786791 675446 786800
rect 675404 784990 675432 785196
rect 675392 784984 675444 784990
rect 675392 784926 675444 784932
rect 675404 784145 675432 784652
rect 675390 784136 675446 784145
rect 675390 784071 675446 784080
rect 675496 783873 675524 783972
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675496 782950 675524 783360
rect 675484 782944 675536 782950
rect 675484 782886 675536 782892
rect 675496 780638 675524 780844
rect 675484 780632 675536 780638
rect 675484 780574 675536 780580
rect 675496 779822 675524 780300
rect 675484 779816 675536 779822
rect 675484 779758 675536 779764
rect 675404 779346 675432 779688
rect 675392 779340 675444 779346
rect 675392 779282 675444 779288
rect 674748 778796 674800 778802
rect 674748 778738 674800 778744
rect 675496 778666 675524 779008
rect 674748 778660 674800 778666
rect 674748 778602 674800 778608
rect 675484 778660 675536 778666
rect 675484 778602 675536 778608
rect 674656 777096 674708 777102
rect 674656 777038 674708 777044
rect 674576 776886 674696 776914
rect 674564 775532 674616 775538
rect 674564 775474 674616 775480
rect 674472 773424 674524 773430
rect 674472 773366 674524 773372
rect 674576 770658 674604 775474
rect 674668 773906 674696 776886
rect 674656 773900 674708 773906
rect 674656 773842 674708 773848
rect 674656 773628 674708 773634
rect 674656 773570 674708 773576
rect 674668 770794 674696 773570
rect 674760 773158 674788 778602
rect 675404 777374 675432 777852
rect 675392 777368 675444 777374
rect 675392 777310 675444 777316
rect 675392 777096 675444 777102
rect 675392 777038 675444 777044
rect 675404 776628 675432 777038
rect 675404 775538 675432 776016
rect 675392 775532 675444 775538
rect 675392 775474 675444 775480
rect 675208 773900 675260 773906
rect 675208 773842 675260 773848
rect 675220 773362 675248 773842
rect 675496 773634 675524 774180
rect 675484 773628 675536 773634
rect 675484 773570 675536 773576
rect 675668 773424 675720 773430
rect 675668 773366 675720 773372
rect 675758 773392 675814 773401
rect 675208 773356 675260 773362
rect 675208 773298 675260 773304
rect 675576 773356 675628 773362
rect 675576 773298 675628 773304
rect 674748 773152 674800 773158
rect 674748 773094 674800 773100
rect 675484 773152 675536 773158
rect 675484 773094 675536 773100
rect 674668 770766 674788 770794
rect 674576 770630 674696 770658
rect 674564 770568 674616 770574
rect 674392 770494 674512 770522
rect 674564 770510 674616 770516
rect 674208 770358 674420 770386
rect 674196 770296 674248 770302
rect 674196 770238 674248 770244
rect 674012 759008 674064 759014
rect 674012 758950 674064 758956
rect 673920 756220 673972 756226
rect 673920 756162 673972 756168
rect 673828 753500 673880 753506
rect 673828 753442 673880 753448
rect 673736 753296 673788 753302
rect 673736 753238 673788 753244
rect 673920 738472 673972 738478
rect 673920 738414 673972 738420
rect 673644 735004 673696 735010
rect 673644 734946 673696 734952
rect 673552 733644 673604 733650
rect 673552 733586 673604 733592
rect 673368 723172 673420 723178
rect 673368 723114 673420 723120
rect 673092 714060 673144 714066
rect 673092 714002 673144 714008
rect 673000 688628 673052 688634
rect 673000 688570 673052 688576
rect 673012 616758 673040 688570
rect 673104 679046 673132 714002
rect 673564 710734 673592 733586
rect 673656 730674 673684 734946
rect 673828 734392 673880 734398
rect 673828 734334 673880 734340
rect 673736 732352 673788 732358
rect 673736 732294 673788 732300
rect 673748 730810 673776 732294
rect 673840 731762 673868 734334
rect 673932 731882 673960 738414
rect 674012 735480 674064 735486
rect 674012 735422 674064 735428
rect 674024 731950 674052 735422
rect 674012 731944 674064 731950
rect 674012 731886 674064 731892
rect 673920 731876 673972 731882
rect 673920 731818 673972 731824
rect 673840 731734 674052 731762
rect 673920 731604 673972 731610
rect 673920 731546 673972 731552
rect 673748 730782 673868 730810
rect 673656 730646 673776 730674
rect 673644 730516 673696 730522
rect 673644 730458 673696 730464
rect 673656 717670 673684 730458
rect 673644 717664 673696 717670
rect 673644 717606 673696 717612
rect 673552 710728 673604 710734
rect 673552 710670 673604 710676
rect 673748 699553 673776 730646
rect 673840 710870 673868 730782
rect 673932 718010 673960 731546
rect 673920 718004 673972 718010
rect 673920 717946 673972 717952
rect 673920 717664 673972 717670
rect 673920 717606 673972 717612
rect 673828 710864 673880 710870
rect 673828 710806 673880 710812
rect 673828 710728 673880 710734
rect 673828 710670 673880 710676
rect 673840 699825 673868 710670
rect 673826 699816 673882 699825
rect 673826 699751 673882 699760
rect 673734 699544 673790 699553
rect 673734 699479 673790 699488
rect 673736 690464 673788 690470
rect 673736 690406 673788 690412
rect 673184 689172 673236 689178
rect 673184 689114 673236 689120
rect 673092 679040 673144 679046
rect 673092 678982 673144 678988
rect 673092 668092 673144 668098
rect 673092 668034 673144 668040
rect 673104 637906 673132 668034
rect 673092 637900 673144 637906
rect 673092 637842 673144 637848
rect 673196 617982 673224 689114
rect 673276 687336 673328 687342
rect 673276 687278 673328 687284
rect 673288 618254 673316 687278
rect 673552 649596 673604 649602
rect 673552 649538 673604 649544
rect 673460 647352 673512 647358
rect 673460 647294 673512 647300
rect 673472 637566 673500 647294
rect 673460 637560 673512 637566
rect 673460 637502 673512 637508
rect 673368 623960 673420 623966
rect 673368 623902 673420 623908
rect 673276 618248 673328 618254
rect 673276 618190 673328 618196
rect 673184 617976 673236 617982
rect 673184 617918 673236 617924
rect 673000 616752 673052 616758
rect 673000 616694 673052 616700
rect 673380 587926 673408 623902
rect 673460 598460 673512 598466
rect 673460 598402 673512 598408
rect 673368 587920 673420 587926
rect 673368 587862 673420 587868
rect 673368 584316 673420 584322
rect 673368 584258 673420 584264
rect 673380 583658 673408 584258
rect 673472 583778 673500 598402
rect 673564 584322 673592 649538
rect 673644 644156 673696 644162
rect 673644 644098 673696 644104
rect 673552 584316 673604 584322
rect 673552 584258 673604 584264
rect 673552 584180 673604 584186
rect 673552 584122 673604 584128
rect 673460 583772 673512 583778
rect 673460 583714 673512 583720
rect 673380 583630 673500 583658
rect 673276 579284 673328 579290
rect 673276 579226 673328 579232
rect 673092 578468 673144 578474
rect 673092 578410 673144 578416
rect 672632 577652 672684 577658
rect 672632 577594 672684 577600
rect 672540 568608 672592 568614
rect 672540 568550 672592 568556
rect 672446 163568 672502 163577
rect 672446 163503 672502 163512
rect 672552 158409 672580 568550
rect 673104 546310 673132 578410
rect 673184 577652 673236 577658
rect 673184 577594 673236 577600
rect 673092 546304 673144 546310
rect 673092 546246 673144 546252
rect 673196 533322 673224 577594
rect 673288 534954 673316 579226
rect 673368 576904 673420 576910
rect 673368 576846 673420 576852
rect 673276 534948 673328 534954
rect 673276 534890 673328 534896
rect 673184 533316 673236 533322
rect 673184 533258 673236 533264
rect 673380 532642 673408 576846
rect 673472 576706 673500 583630
rect 673460 576700 673512 576706
rect 673460 576642 673512 576648
rect 673564 576094 673592 584122
rect 673552 576088 673604 576094
rect 673552 576030 673604 576036
rect 673656 572830 673684 644098
rect 673748 620906 673776 690406
rect 673828 685500 673880 685506
rect 673828 685442 673880 685448
rect 673840 623762 673868 685442
rect 673932 667894 673960 717606
rect 674024 699689 674052 731734
rect 674208 718146 674236 770238
rect 674288 770228 674340 770234
rect 674288 770170 674340 770176
rect 674196 718140 674248 718146
rect 674196 718082 674248 718088
rect 674196 718004 674248 718010
rect 674196 717946 674248 717952
rect 674208 711890 674236 717946
rect 674300 711958 674328 770170
rect 674288 711952 674340 711958
rect 674288 711894 674340 711900
rect 674196 711884 674248 711890
rect 674196 711826 674248 711832
rect 674392 708286 674420 770358
rect 674484 709306 674512 770494
rect 674576 712026 674604 770510
rect 674668 738478 674696 770630
rect 674656 738472 674708 738478
rect 674656 738414 674708 738420
rect 674656 738336 674708 738342
rect 674656 738278 674708 738284
rect 674668 732086 674696 738278
rect 674656 732080 674708 732086
rect 674656 732022 674708 732028
rect 674656 731944 674708 731950
rect 674656 731886 674708 731892
rect 674564 712020 674616 712026
rect 674564 711962 674616 711968
rect 674668 710734 674696 731886
rect 674760 712094 674788 770766
rect 675496 744161 675524 773094
rect 675588 754225 675616 773298
rect 675574 754216 675630 754225
rect 675574 754151 675630 754160
rect 675482 744152 675538 744161
rect 675482 744087 675538 744096
rect 675680 744025 675708 773366
rect 675758 773327 675814 773336
rect 675772 753817 675800 773327
rect 679070 772712 679126 772721
rect 679070 772647 679126 772656
rect 678978 761288 679034 761297
rect 678978 761223 679034 761232
rect 676218 760880 676274 760889
rect 676218 760815 676274 760824
rect 676126 760472 676182 760481
rect 676126 760407 676182 760416
rect 676140 759354 676168 760407
rect 676232 759626 676260 760815
rect 676310 759656 676366 759665
rect 676220 759620 676272 759626
rect 676310 759591 676366 759600
rect 676220 759562 676272 759568
rect 676128 759348 676180 759354
rect 676128 759290 676180 759296
rect 676036 759144 676088 759150
rect 676034 759112 676036 759121
rect 676088 759112 676090 759121
rect 676324 759082 676352 759591
rect 678992 759490 679020 761223
rect 679084 759665 679112 772647
rect 679070 759656 679126 759665
rect 679070 759591 679126 759600
rect 678980 759484 679032 759490
rect 678980 759426 679032 759432
rect 676034 759047 676090 759056
rect 676312 759076 676364 759082
rect 676312 759018 676364 759024
rect 676036 759008 676088 759014
rect 676036 758950 676088 758956
rect 676048 756673 676076 758950
rect 678978 758432 679034 758441
rect 678978 758367 679034 758376
rect 676310 758024 676366 758033
rect 676310 757959 676366 757968
rect 676126 757616 676182 757625
rect 676126 757551 676182 757560
rect 676034 756664 676090 756673
rect 676034 756599 676090 756608
rect 676140 756362 676168 757551
rect 676218 757208 676274 757217
rect 676218 757143 676274 757152
rect 676232 756498 676260 757143
rect 676220 756492 676272 756498
rect 676220 756434 676272 756440
rect 676324 756430 676352 757959
rect 676312 756424 676364 756430
rect 676312 756366 676364 756372
rect 676128 756356 676180 756362
rect 676128 756298 676180 756304
rect 678992 756294 679020 758367
rect 678980 756288 679032 756294
rect 678980 756230 679032 756236
rect 676036 756220 676088 756226
rect 676036 756162 676088 756168
rect 676048 755041 676076 756162
rect 676128 756152 676180 756158
rect 676128 756094 676180 756100
rect 676140 755585 676168 756094
rect 676126 755576 676182 755585
rect 676126 755511 676182 755520
rect 676034 755032 676090 755041
rect 676034 754967 676090 754976
rect 675758 753808 675814 753817
rect 675758 753743 675814 753752
rect 676036 753500 676088 753506
rect 676036 753442 676088 753448
rect 676048 753409 676076 753442
rect 676034 753400 676090 753409
rect 676034 753335 676090 753344
rect 676036 753296 676088 753302
rect 676036 753238 676088 753244
rect 676048 753001 676076 753238
rect 676034 752992 676090 753001
rect 676034 752927 676090 752936
rect 678978 751088 679034 751097
rect 678978 751023 679034 751032
rect 678992 750281 679020 751023
rect 678978 750272 679034 750281
rect 678978 750207 679034 750216
rect 678992 749834 679020 750207
rect 678980 749828 679032 749834
rect 678980 749770 679032 749776
rect 675666 744016 675722 744025
rect 675666 743951 675722 743960
rect 675772 742937 675800 743308
rect 675758 742928 675814 742937
rect 675758 742863 675814 742872
rect 675772 742529 675800 742696
rect 675758 742520 675814 742529
rect 675758 742455 675814 742464
rect 675496 741713 675524 742016
rect 675482 741704 675538 741713
rect 675482 741639 675538 741648
rect 675404 739809 675432 740180
rect 675390 739800 675446 739809
rect 675390 739735 675446 739744
rect 675404 739129 675432 739636
rect 675390 739120 675446 739129
rect 675390 739055 675446 739064
rect 675680 738585 675708 739024
rect 675666 738576 675722 738585
rect 675666 738511 675722 738520
rect 675772 738041 675800 738344
rect 675758 738032 675814 738041
rect 675758 737967 675814 737976
rect 675404 735486 675432 735896
rect 675392 735480 675444 735486
rect 675392 735422 675444 735428
rect 675404 735010 675432 735319
rect 675392 735004 675444 735010
rect 675392 734946 675444 734952
rect 675404 734398 675432 734672
rect 675392 734392 675444 734398
rect 675392 734334 675444 734340
rect 675404 733650 675432 734031
rect 675392 733644 675444 733650
rect 675392 733586 675444 733592
rect 675404 732358 675432 732836
rect 675392 732352 675444 732358
rect 675392 732294 675444 732300
rect 675392 732080 675444 732086
rect 675392 732022 675444 732028
rect 675404 731612 675432 732022
rect 675404 730522 675432 731000
rect 675392 730516 675444 730522
rect 675392 730458 675444 730464
rect 675680 728686 675708 729164
rect 675668 728680 675720 728686
rect 675668 728622 675720 728628
rect 675668 728408 675720 728414
rect 675668 728350 675720 728356
rect 674840 718140 674892 718146
rect 674840 718082 674892 718088
rect 674748 712088 674800 712094
rect 674748 712030 674800 712036
rect 674656 710728 674708 710734
rect 674656 710670 674708 710676
rect 674472 709300 674524 709306
rect 674472 709242 674524 709248
rect 674380 708280 674432 708286
rect 674380 708222 674432 708228
rect 674852 707878 674880 718082
rect 675484 710864 675536 710870
rect 675484 710806 675536 710812
rect 674840 707872 674892 707878
rect 674840 707814 674892 707820
rect 674564 699780 674616 699786
rect 674564 699722 674616 699728
rect 674010 699680 674066 699689
rect 674010 699615 674066 699624
rect 674472 691416 674524 691422
rect 674472 691358 674524 691364
rect 674484 687070 674512 691358
rect 674472 687064 674524 687070
rect 674472 687006 674524 687012
rect 674288 683664 674340 683670
rect 674288 683606 674340 683612
rect 673920 667888 673972 667894
rect 673920 667830 673972 667836
rect 673920 645448 673972 645454
rect 673920 645390 673972 645396
rect 673828 623756 673880 623762
rect 673828 623698 673880 623704
rect 673736 620900 673788 620906
rect 673736 620842 673788 620848
rect 673736 599004 673788 599010
rect 673736 598946 673788 598952
rect 673644 572824 673696 572830
rect 673644 572766 673696 572772
rect 673552 559564 673604 559570
rect 673552 559506 673604 559512
rect 673460 554600 673512 554606
rect 673460 554542 673512 554548
rect 672816 532636 672868 532642
rect 672816 532578 672868 532584
rect 673368 532636 673420 532642
rect 673368 532578 673420 532584
rect 672632 524476 672684 524482
rect 672632 524418 672684 524424
rect 672538 158400 672594 158409
rect 672538 158335 672594 158344
rect 672644 153377 672672 524418
rect 672724 480752 672776 480758
rect 672724 480694 672776 480700
rect 672630 153368 672686 153377
rect 672630 153303 672686 153312
rect 672736 148209 672764 480694
rect 672828 278594 672856 532578
rect 673472 482934 673500 554542
rect 673564 487966 673592 559506
rect 673644 553240 673696 553246
rect 673644 553182 673696 553188
rect 673552 487960 673604 487966
rect 673552 487902 673604 487908
rect 673656 483002 673684 553182
rect 673748 527882 673776 598946
rect 673828 597168 673880 597174
rect 673828 597110 673880 597116
rect 673840 583930 673868 597110
rect 673932 584186 673960 645390
rect 674012 642116 674064 642122
rect 674012 642058 674064 642064
rect 673920 584180 673972 584186
rect 673920 584122 673972 584128
rect 673840 583902 673960 583930
rect 673828 583772 673880 583778
rect 673828 583714 673880 583720
rect 673736 527876 673788 527882
rect 673736 527818 673788 527824
rect 673840 527134 673868 583714
rect 673932 583710 673960 583902
rect 673920 583704 673972 583710
rect 673920 583646 673972 583652
rect 674024 573646 674052 642058
rect 674196 640280 674248 640286
rect 674196 640222 674248 640228
rect 674208 576842 674236 640222
rect 674300 620974 674328 683606
rect 674472 669792 674524 669798
rect 674472 669734 674524 669740
rect 674380 643408 674432 643414
rect 674380 643350 674432 643356
rect 674288 620968 674340 620974
rect 674288 620910 674340 620916
rect 674392 607753 674420 643350
rect 674484 626550 674512 669734
rect 674576 667826 674604 699722
rect 675496 699718 675524 710806
rect 675576 710728 675628 710734
rect 675576 710670 675628 710676
rect 675588 699786 675616 710670
rect 675576 699780 675628 699786
rect 675576 699722 675628 699728
rect 674748 699712 674800 699718
rect 674748 699654 674800 699660
rect 675484 699712 675536 699718
rect 675484 699654 675536 699660
rect 674656 699644 674708 699650
rect 674656 699586 674708 699592
rect 674564 667820 674616 667826
rect 674564 667762 674616 667768
rect 674668 665174 674696 699586
rect 674760 671294 674788 699654
rect 675680 699650 675708 728350
rect 678980 723172 679032 723178
rect 678980 723114 679032 723120
rect 676034 716544 676090 716553
rect 676034 716479 676090 716488
rect 675944 716168 675996 716174
rect 675942 716136 675944 716145
rect 675996 716136 675998 716145
rect 675942 716071 675998 716080
rect 675944 715760 675996 715766
rect 675942 715728 675944 715737
rect 675996 715728 675998 715737
rect 675942 715663 675998 715672
rect 675944 715352 675996 715358
rect 675942 715320 675944 715329
rect 675996 715320 675998 715329
rect 675942 715255 675998 715264
rect 676048 715018 676076 716479
rect 676036 715012 676088 715018
rect 676036 714954 676088 714960
rect 676034 714912 676090 714921
rect 676034 714847 676036 714856
rect 676088 714847 676090 714856
rect 676036 714818 676088 714824
rect 678992 714513 679020 723114
rect 678978 714504 679034 714513
rect 678978 714439 679034 714448
rect 676034 714096 676090 714105
rect 676034 714031 676036 714040
rect 676088 714031 676090 714040
rect 676036 714002 676088 714008
rect 676036 713720 676088 713726
rect 676034 713688 676036 713697
rect 676088 713688 676090 713697
rect 676034 713623 676090 713632
rect 676034 713280 676090 713289
rect 676034 713215 676036 713224
rect 676088 713215 676090 713224
rect 676036 713186 676088 713192
rect 676034 712872 676090 712881
rect 676034 712807 676036 712816
rect 676088 712807 676090 712816
rect 676036 712778 676088 712784
rect 676034 712464 676090 712473
rect 676034 712399 676036 712408
rect 676088 712399 676090 712408
rect 676036 712370 676088 712376
rect 676036 712088 676088 712094
rect 676036 712030 676088 712036
rect 675944 712020 675996 712026
rect 675944 711962 675996 711968
rect 675852 711952 675904 711958
rect 675852 711894 675904 711900
rect 675760 711884 675812 711890
rect 675760 711826 675812 711832
rect 675772 711657 675800 711826
rect 675758 711648 675814 711657
rect 675758 711583 675814 711592
rect 675864 710841 675892 711894
rect 675850 710832 675906 710841
rect 675850 710767 675906 710776
rect 675956 710433 675984 711962
rect 675942 710424 675998 710433
rect 675942 710359 675998 710368
rect 676048 710025 676076 712030
rect 676310 711886 676366 711895
rect 676310 711821 676366 711830
rect 676954 711886 677010 711895
rect 676954 711821 677010 711830
rect 676034 710016 676090 710025
rect 676034 709951 676090 709960
rect 676036 709300 676088 709306
rect 676036 709242 676088 709248
rect 676048 708393 676076 709242
rect 676034 708384 676090 708393
rect 676034 708319 676090 708328
rect 676036 708280 676088 708286
rect 676036 708222 676088 708228
rect 676048 707985 676076 708222
rect 676034 707976 676090 707985
rect 676034 707911 676090 707920
rect 676036 707872 676088 707878
rect 676036 707814 676088 707820
rect 676048 707577 676076 707814
rect 676034 707568 676090 707577
rect 676034 707503 676090 707512
rect 676036 707464 676088 707470
rect 676036 707406 676088 707412
rect 676048 706761 676076 707406
rect 676324 707169 676352 711821
rect 676968 707470 676996 711821
rect 676956 707464 677008 707470
rect 676956 707406 677008 707412
rect 676310 707160 676366 707169
rect 676310 707095 676366 707104
rect 676034 706752 676090 706761
rect 676034 706687 676090 706696
rect 676034 706344 676090 706353
rect 676034 706279 676090 706288
rect 676048 705158 676076 706279
rect 676036 705152 676088 705158
rect 676034 705120 676036 705129
rect 676088 705120 676090 705129
rect 676034 705055 676090 705064
rect 676048 705029 676076 705055
rect 675668 699644 675720 699650
rect 675668 699586 675720 699592
rect 675496 698193 675524 698323
rect 675482 698184 675538 698193
rect 675482 698119 675538 698128
rect 675404 697241 675432 697680
rect 675390 697232 675446 697241
rect 675390 697167 675446 697176
rect 675404 696697 675432 697035
rect 675390 696688 675446 696697
rect 675390 696623 675446 696632
rect 675404 695065 675432 695195
rect 675390 695056 675446 695065
rect 675390 694991 675446 695000
rect 675496 694249 675524 694620
rect 675482 694240 675538 694249
rect 675482 694175 675538 694184
rect 675404 693705 675432 694008
rect 675390 693696 675446 693705
rect 675390 693631 675446 693640
rect 675772 693025 675800 693328
rect 675758 693016 675814 693025
rect 675758 692951 675814 692960
rect 675404 690470 675432 690880
rect 675392 690464 675444 690470
rect 675392 690406 675444 690412
rect 675772 690169 675800 690336
rect 675758 690160 675814 690169
rect 675758 690095 675814 690104
rect 675496 689178 675524 689656
rect 675484 689172 675536 689178
rect 675484 689114 675536 689120
rect 675404 688634 675432 689044
rect 675392 688628 675444 688634
rect 675392 688570 675444 688576
rect 675404 687342 675432 687820
rect 675392 687336 675444 687342
rect 675392 687278 675444 687284
rect 675484 687064 675536 687070
rect 675484 687006 675536 687012
rect 675496 686664 675524 687006
rect 675404 685506 675432 685984
rect 675392 685500 675444 685506
rect 675392 685442 675444 685448
rect 675496 683670 675524 684148
rect 675484 683664 675536 683670
rect 675484 683606 675536 683612
rect 678980 679040 679032 679046
rect 678980 678982 679032 678988
rect 676220 671560 676272 671566
rect 676218 671528 676220 671537
rect 676272 671528 676274 671537
rect 676218 671463 676274 671472
rect 674748 671288 674800 671294
rect 674748 671230 674800 671236
rect 675208 671288 675260 671294
rect 675208 671230 675260 671236
rect 674748 667956 674800 667962
rect 674748 667898 674800 667904
rect 674656 665168 674708 665174
rect 674656 665110 674708 665116
rect 674656 647760 674708 647766
rect 674656 647702 674708 647708
rect 674564 644836 674616 644842
rect 674564 644778 674616 644784
rect 674576 638602 674604 644778
rect 674668 638858 674696 647702
rect 674760 647358 674788 667898
rect 675220 664766 675248 671230
rect 676034 670984 676090 670993
rect 676034 670919 676090 670928
rect 676048 670818 676076 670919
rect 676036 670812 676088 670818
rect 676036 670754 676088 670760
rect 676036 670608 676088 670614
rect 676034 670576 676036 670585
rect 676088 670576 676090 670585
rect 676034 670511 676090 670520
rect 676220 670336 676272 670342
rect 676218 670304 676220 670313
rect 676272 670304 676274 670313
rect 676218 670239 676274 670248
rect 676036 669792 676088 669798
rect 676034 669760 676036 669769
rect 676088 669760 676090 669769
rect 676034 669695 676090 669704
rect 678992 669497 679020 678982
rect 678978 669488 679034 669497
rect 678978 669423 679034 669432
rect 676034 668944 676090 668953
rect 676034 668879 676090 668888
rect 675942 668128 675998 668137
rect 675942 668063 675944 668072
rect 675996 668063 675998 668072
rect 675944 668034 675996 668040
rect 676048 667962 676076 668879
rect 676220 668704 676272 668710
rect 676218 668672 676220 668681
rect 676272 668672 676274 668681
rect 676218 668607 676274 668616
rect 676036 667956 676088 667962
rect 676036 667898 676088 667904
rect 676128 667888 676180 667894
rect 676128 667830 676180 667836
rect 676036 667820 676088 667826
rect 676036 667762 676088 667768
rect 675944 667752 675996 667758
rect 675942 667720 675944 667729
rect 675996 667720 675998 667729
rect 675942 667655 675998 667664
rect 676048 665281 676076 667762
rect 676140 666641 676168 667830
rect 676126 666632 676182 666641
rect 676126 666567 676182 666576
rect 676034 665272 676090 665281
rect 676034 665207 676090 665216
rect 676036 665168 676088 665174
rect 676036 665110 676088 665116
rect 676048 664873 676076 665110
rect 676034 664864 676090 664873
rect 676034 664799 676090 664808
rect 675208 664760 675260 664766
rect 675208 664702 675260 664708
rect 676036 664760 676088 664766
rect 676036 664702 676088 664708
rect 676048 663241 676076 664702
rect 676034 663232 676090 663241
rect 676034 663167 676090 663176
rect 678978 660920 679034 660929
rect 678978 660855 679034 660864
rect 678992 660113 679020 660855
rect 678978 660104 679034 660113
rect 678978 660039 679034 660048
rect 678992 659734 679020 660039
rect 678980 659728 679032 659734
rect 678980 659670 679032 659676
rect 675404 652633 675432 653140
rect 675390 652624 675446 652633
rect 675390 652559 675446 652568
rect 675496 652225 675524 652460
rect 675482 652216 675538 652225
rect 675482 652151 675538 652160
rect 675404 651681 675432 651848
rect 675390 651672 675446 651681
rect 675390 651607 675446 651616
rect 675404 649602 675432 650012
rect 675392 649596 675444 649602
rect 675392 649538 675444 649544
rect 675772 649233 675800 649468
rect 675758 649224 675814 649233
rect 675758 649159 675814 649168
rect 675680 648689 675708 648788
rect 675666 648680 675722 648689
rect 675666 648615 675722 648624
rect 675496 647766 675524 648176
rect 675484 647760 675536 647766
rect 675484 647702 675536 647708
rect 674748 647352 674800 647358
rect 674748 647294 674800 647300
rect 674748 647216 674800 647222
rect 674748 647158 674800 647164
rect 674760 641918 674788 647158
rect 675404 645454 675432 645660
rect 675392 645448 675444 645454
rect 675392 645390 675444 645396
rect 675404 644842 675432 645116
rect 675392 644836 675444 644842
rect 675392 644778 675444 644784
rect 675404 644162 675432 644475
rect 675392 644156 675444 644162
rect 675392 644098 675444 644104
rect 675404 643414 675432 643824
rect 675392 643408 675444 643414
rect 675392 643350 675444 643356
rect 675404 642122 675432 642635
rect 675392 642116 675444 642122
rect 675392 642058 675444 642064
rect 674748 641912 674800 641918
rect 674748 641854 674800 641860
rect 675392 641912 675444 641918
rect 675392 641854 675444 641860
rect 675404 641444 675432 641854
rect 675404 640286 675432 640795
rect 675392 640280 675444 640286
rect 675392 640222 675444 640228
rect 674656 638852 674708 638858
rect 674656 638794 674708 638800
rect 675208 638716 675260 638722
rect 675208 638658 675260 638664
rect 674576 638574 674788 638602
rect 674564 638444 674616 638450
rect 674564 638386 674616 638392
rect 674472 626544 674524 626550
rect 674472 626486 674524 626492
rect 674472 608796 674524 608802
rect 674472 608738 674524 608744
rect 674378 607744 674434 607753
rect 674378 607679 674434 607688
rect 674288 600432 674340 600438
rect 674288 600374 674340 600380
rect 674196 576836 674248 576842
rect 674196 576778 674248 576784
rect 674012 573640 674064 573646
rect 674012 573582 674064 573588
rect 673920 555280 673972 555286
rect 673920 555222 673972 555228
rect 673828 527128 673880 527134
rect 673828 527070 673880 527076
rect 673932 487150 673960 555222
rect 674012 553784 674064 553790
rect 674012 553726 674064 553732
rect 673920 487144 673972 487150
rect 673920 487086 673972 487092
rect 674024 483585 674052 553726
rect 674196 551948 674248 551954
rect 674196 551890 674248 551896
rect 674208 485518 674236 551890
rect 674300 531146 674328 600374
rect 674484 596630 674512 608738
rect 674472 596624 674524 596630
rect 674472 596566 674524 596572
rect 674472 595332 674524 595338
rect 674472 595274 674524 595280
rect 674380 593700 674432 593706
rect 674380 593642 674432 593648
rect 674392 583794 674420 593642
rect 674484 583914 674512 595274
rect 674472 583908 674524 583914
rect 674472 583850 674524 583856
rect 674392 583766 674512 583794
rect 674380 583704 674432 583710
rect 674380 583646 674432 583652
rect 674288 531140 674340 531146
rect 674288 531082 674340 531088
rect 674392 529514 674420 583646
rect 674484 529922 674512 583766
rect 674576 576774 674604 638386
rect 674760 607481 674788 638574
rect 675220 638246 675248 638658
rect 675496 638450 675524 638928
rect 675484 638444 675536 638450
rect 675484 638386 675536 638392
rect 675208 638240 675260 638246
rect 675208 638182 675260 638188
rect 675668 638240 675720 638246
rect 675668 638182 675720 638188
rect 675680 608802 675708 638182
rect 679164 637900 679216 637906
rect 679164 637842 679216 637848
rect 679072 637560 679124 637566
rect 679072 637502 679124 637508
rect 676036 626544 676088 626550
rect 676036 626486 676088 626492
rect 676048 625161 676076 626486
rect 678978 626104 679034 626113
rect 678978 626039 679034 626048
rect 676218 625696 676274 625705
rect 676218 625631 676274 625640
rect 676034 625152 676090 625161
rect 676034 625087 676090 625096
rect 676126 624472 676182 624481
rect 676126 624407 676182 624416
rect 676036 623960 676088 623966
rect 676034 623928 676036 623937
rect 676088 623928 676090 623937
rect 676034 623863 676090 623872
rect 676140 623830 676168 624407
rect 676232 624170 676260 625631
rect 676310 625288 676366 625297
rect 676310 625223 676366 625232
rect 676220 624164 676272 624170
rect 676220 624106 676272 624112
rect 676324 623898 676352 625223
rect 678992 624034 679020 626039
rect 679084 624481 679112 637502
rect 679070 624472 679126 624481
rect 679070 624407 679126 624416
rect 678980 624028 679032 624034
rect 678980 623970 679032 623976
rect 676312 623892 676364 623898
rect 676312 623834 676364 623840
rect 676128 623824 676180 623830
rect 676128 623766 676180 623772
rect 676036 623756 676088 623762
rect 676036 623698 676088 623704
rect 676048 621489 676076 623698
rect 679176 623665 679204 637842
rect 679162 623656 679218 623665
rect 679162 623591 679218 623600
rect 678978 623248 679034 623257
rect 678978 623183 679034 623192
rect 676218 622024 676274 622033
rect 676218 621959 676274 621968
rect 676034 621480 676090 621489
rect 676034 621415 676090 621424
rect 676232 621042 676260 621959
rect 678992 621110 679020 623183
rect 678980 621104 679032 621110
rect 678980 621046 679032 621052
rect 676220 621036 676272 621042
rect 676220 620978 676272 620984
rect 676036 620968 676088 620974
rect 676036 620910 676088 620916
rect 676048 619857 676076 620910
rect 676128 620900 676180 620906
rect 676128 620842 676180 620848
rect 676140 620401 676168 620842
rect 676126 620392 676182 620401
rect 676126 620327 676182 620336
rect 676034 619848 676090 619857
rect 676034 619783 676090 619792
rect 676036 618248 676088 618254
rect 676034 618216 676036 618225
rect 676088 618216 676090 618225
rect 676034 618151 676090 618160
rect 676220 617976 676272 617982
rect 676218 617944 676220 617953
rect 676272 617944 676274 617953
rect 676218 617879 676274 617888
rect 676220 616752 676272 616758
rect 676218 616720 676220 616729
rect 676272 616720 676274 616729
rect 676218 616655 676274 616664
rect 678978 615904 679034 615913
rect 678978 615839 679034 615848
rect 678992 615097 679020 615839
rect 678978 615088 679034 615097
rect 678978 615023 679034 615032
rect 678992 614650 679020 615023
rect 678980 614644 679032 614650
rect 678980 614586 679032 614592
rect 675668 608796 675720 608802
rect 675668 608738 675720 608744
rect 675496 607617 675524 608124
rect 675482 607608 675538 607617
rect 675482 607543 675538 607552
rect 674746 607472 674802 607481
rect 674746 607407 674802 607416
rect 675772 607345 675800 607479
rect 675758 607336 675814 607345
rect 675758 607271 675814 607280
rect 675404 606529 675432 606832
rect 675390 606520 675446 606529
rect 675390 606455 675446 606464
rect 675404 604761 675432 604996
rect 675390 604752 675446 604761
rect 675390 604687 675446 604696
rect 675404 604353 675432 604452
rect 675390 604344 675446 604353
rect 675390 604279 675446 604288
rect 675496 603537 675524 603772
rect 675482 603528 675538 603537
rect 675482 603463 675538 603472
rect 674656 603084 674708 603090
rect 674656 603026 674708 603032
rect 674668 596902 674696 603026
rect 675772 602993 675800 603160
rect 675758 602984 675814 602993
rect 675758 602919 675814 602928
rect 675496 600438 675524 600644
rect 675484 600432 675536 600438
rect 675484 600374 675536 600380
rect 675496 599622 675524 600100
rect 674748 599616 674800 599622
rect 674748 599558 674800 599564
rect 675484 599616 675536 599622
rect 675484 599558 675536 599564
rect 674656 596896 674708 596902
rect 674656 596838 674708 596844
rect 674760 596714 674788 599558
rect 675404 599010 675432 599488
rect 675392 599004 675444 599010
rect 675392 598946 675444 598952
rect 675496 598466 675524 598808
rect 675484 598460 675536 598466
rect 675484 598402 675536 598408
rect 675404 597174 675432 597652
rect 675392 597168 675444 597174
rect 675392 597110 675444 597116
rect 675392 596896 675444 596902
rect 675392 596838 675444 596844
rect 674668 596686 674788 596714
rect 674564 576768 674616 576774
rect 674564 576710 674616 576716
rect 674668 564505 674696 596686
rect 674748 596624 674800 596630
rect 674748 596566 674800 596572
rect 674760 584050 674788 596566
rect 675404 596428 675432 596838
rect 675404 595338 675432 595816
rect 675392 595332 675444 595338
rect 675392 595274 675444 595280
rect 675496 593706 675524 593980
rect 675484 593700 675536 593706
rect 675484 593642 675536 593648
rect 678980 587920 679032 587926
rect 678980 587862 679032 587868
rect 674748 584044 674800 584050
rect 674748 583986 674800 583992
rect 675668 584044 675720 584050
rect 675668 583986 675720 583992
rect 674748 583908 674800 583914
rect 674748 583850 674800 583856
rect 674654 564496 674710 564505
rect 674654 564431 674710 564440
rect 674564 548344 674616 548350
rect 674564 548286 674616 548292
rect 674472 529916 674524 529922
rect 674472 529858 674524 529864
rect 674380 529508 674432 529514
rect 674380 529450 674432 529456
rect 674576 485790 674604 548286
rect 674656 548276 674708 548282
rect 674656 548218 674708 548224
rect 674668 488238 674696 548218
rect 674760 532710 674788 583850
rect 675680 572121 675708 583986
rect 676310 580952 676366 580961
rect 676310 580887 676366 580896
rect 676126 580544 676182 580553
rect 676126 580479 676182 580488
rect 676036 580236 676088 580242
rect 676036 580178 676088 580184
rect 676048 579873 676076 580178
rect 676140 580106 676168 580479
rect 676218 580136 676274 580145
rect 676128 580100 676180 580106
rect 676218 580071 676274 580080
rect 676128 580042 676180 580048
rect 676232 579970 676260 580071
rect 676220 579964 676272 579970
rect 676220 579906 676272 579912
rect 676034 579864 676090 579873
rect 676324 579834 676352 580887
rect 676034 579799 676090 579808
rect 676312 579828 676364 579834
rect 676312 579770 676364 579776
rect 678992 579329 679020 587862
rect 676218 579320 676274 579329
rect 676218 579255 676220 579264
rect 676272 579255 676274 579264
rect 678978 579320 679034 579329
rect 678978 579255 679034 579264
rect 676220 579226 676272 579232
rect 676218 578504 676274 578513
rect 676218 578439 676220 578448
rect 676272 578439 676274 578448
rect 676220 578410 676272 578416
rect 676218 577688 676274 577697
rect 676218 577623 676220 577632
rect 676272 577623 676274 577632
rect 676220 577594 676272 577600
rect 676218 577280 676274 577289
rect 676218 577215 676274 577224
rect 676034 577008 676090 577017
rect 676232 576978 676260 577215
rect 676034 576943 676090 576952
rect 676220 576972 676272 576978
rect 676048 576910 676076 576943
rect 676220 576914 676272 576920
rect 676036 576904 676088 576910
rect 676036 576846 676088 576852
rect 675944 576836 675996 576842
rect 675944 576778 675996 576784
rect 675956 576201 675984 576778
rect 676036 576768 676088 576774
rect 676036 576710 676088 576716
rect 675942 576192 675998 576201
rect 675942 576127 675998 576136
rect 675944 576088 675996 576094
rect 675944 576030 675996 576036
rect 675956 574977 675984 576030
rect 675942 574968 675998 574977
rect 675942 574903 675998 574912
rect 676048 574569 676076 576710
rect 676128 576700 676180 576706
rect 676128 576642 676180 576648
rect 676140 575657 676168 576642
rect 676126 575648 676182 575657
rect 676126 575583 676182 575592
rect 676034 574560 676090 574569
rect 676034 574495 676090 574504
rect 676036 573640 676088 573646
rect 676036 573582 676088 573588
rect 676048 572937 676076 573582
rect 676034 572928 676090 572937
rect 676034 572863 676090 572872
rect 676036 572824 676088 572830
rect 676036 572766 676088 572772
rect 676048 572529 676076 572766
rect 676034 572520 676090 572529
rect 676034 572455 676090 572464
rect 675666 572112 675722 572121
rect 675666 572047 675722 572056
rect 678978 570752 679034 570761
rect 678978 570687 679034 570696
rect 678992 569945 679020 570687
rect 678978 569936 679034 569945
rect 678978 569871 679034 569880
rect 678992 568614 679020 569871
rect 678980 568608 679032 568614
rect 678980 568550 679032 568556
rect 675772 562465 675800 562904
rect 675758 562456 675814 562465
rect 675758 562391 675814 562400
rect 675772 562057 675800 562292
rect 675758 562048 675814 562057
rect 675758 561983 675814 561992
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675496 559570 675524 559776
rect 675484 559564 675536 559570
rect 675484 559506 675536 559512
rect 675404 558793 675432 559232
rect 675390 558784 675446 558793
rect 675390 558719 675446 558728
rect 675772 558385 675800 558620
rect 675758 558376 675814 558385
rect 675758 558311 675814 558320
rect 675772 557569 675800 557940
rect 675758 557560 675814 557569
rect 675758 557495 675814 557504
rect 675300 556164 675352 556170
rect 675300 556106 675352 556112
rect 675312 551253 675340 556106
rect 675404 555286 675432 555492
rect 675392 555280 675444 555286
rect 675392 555222 675444 555228
rect 675404 554606 675432 554919
rect 675392 554600 675444 554606
rect 675392 554542 675444 554548
rect 675404 553790 675432 554268
rect 675392 553784 675444 553790
rect 675392 553726 675444 553732
rect 675404 553246 675432 553656
rect 675392 553240 675444 553246
rect 675392 553182 675444 553188
rect 675404 551954 675432 552432
rect 675392 551948 675444 551954
rect 675392 551890 675444 551896
rect 675312 551225 675418 551253
rect 675312 550582 675418 550610
rect 675312 548282 675340 550582
rect 675404 548350 675432 548760
rect 675392 548344 675444 548350
rect 675392 548286 675444 548292
rect 675300 548276 675352 548282
rect 675300 548218 675352 548224
rect 679072 546304 679124 546310
rect 679072 546246 679124 546252
rect 676218 535936 676274 535945
rect 676218 535871 676274 535880
rect 676232 535770 676260 535871
rect 676220 535764 676272 535770
rect 676034 535732 676090 535741
rect 676220 535706 676272 535712
rect 676034 535667 676090 535676
rect 676048 535634 676076 535667
rect 676036 535628 676088 535634
rect 676036 535570 676088 535576
rect 678978 535120 679034 535129
rect 678978 535055 679034 535064
rect 676036 534948 676088 534954
rect 676034 534916 676036 534925
rect 676088 534916 676090 534925
rect 676034 534851 676090 534860
rect 676126 534304 676182 534313
rect 676126 534239 676182 534248
rect 676036 533316 676088 533322
rect 676034 533284 676036 533293
rect 676088 533284 676090 533293
rect 676034 533219 676090 533228
rect 675942 532876 675998 532885
rect 675852 532840 675904 532846
rect 676140 532846 676168 534239
rect 678992 532914 679020 535055
rect 679084 534313 679112 546246
rect 679070 534304 679126 534313
rect 679070 534239 679126 534248
rect 679070 533488 679126 533497
rect 679070 533423 679126 533432
rect 678980 532908 679032 532914
rect 678980 532850 679032 532856
rect 675942 532811 675998 532820
rect 676128 532840 676180 532846
rect 675852 532782 675904 532788
rect 674748 532704 674800 532710
rect 674748 532646 674800 532652
rect 675864 524006 675892 532782
rect 675852 524000 675904 524006
rect 675852 523942 675904 523948
rect 675956 496814 675984 532811
rect 676128 532782 676180 532788
rect 676036 532704 676088 532710
rect 676036 532646 676088 532652
rect 676218 532672 676274 532681
rect 676048 531253 676076 532646
rect 676218 532607 676220 532616
rect 676272 532607 676274 532616
rect 676220 532578 676272 532584
rect 676126 531856 676182 531865
rect 676126 531791 676182 531800
rect 676034 531244 676090 531253
rect 676034 531179 676090 531188
rect 676036 531140 676088 531146
rect 676036 531082 676088 531088
rect 676048 530029 676076 531082
rect 676034 530020 676090 530029
rect 676034 529955 676090 529964
rect 676036 529916 676088 529922
rect 676036 529858 676088 529864
rect 676048 529621 676076 529858
rect 676034 529612 676090 529621
rect 676034 529547 676090 529556
rect 676036 529508 676088 529514
rect 676036 529450 676088 529456
rect 676048 527989 676076 529450
rect 676034 527980 676090 527989
rect 676034 527915 676090 527924
rect 676036 527876 676088 527882
rect 676036 527818 676088 527824
rect 676048 527581 676076 527818
rect 676034 527572 676090 527581
rect 676034 527507 676090 527516
rect 676036 527128 676088 527134
rect 676036 527070 676088 527076
rect 676048 526357 676076 527070
rect 676034 526348 676090 526357
rect 676034 526283 676090 526292
rect 676140 524090 676168 531791
rect 678978 525736 679034 525745
rect 678978 525671 679034 525680
rect 678992 524929 679020 525671
rect 678978 524920 679034 524929
rect 678978 524855 679034 524864
rect 678992 524482 679020 524855
rect 678980 524476 679032 524482
rect 678980 524418 679032 524424
rect 679084 524414 679112 533423
rect 677498 524408 677550 524414
rect 677498 524350 677550 524356
rect 679072 524408 679124 524414
rect 679072 524350 679124 524356
rect 675864 496786 675984 496814
rect 676048 524062 676168 524090
rect 675576 492244 675628 492250
rect 675576 492186 675628 492192
rect 675588 488481 675616 492186
rect 675864 489297 675892 496786
rect 676048 492250 676076 524062
rect 676128 524000 676180 524006
rect 676128 523942 676180 523948
rect 676036 492244 676088 492250
rect 676036 492186 676088 492192
rect 676034 492144 676090 492153
rect 676034 492079 676090 492088
rect 675942 491736 675998 491745
rect 676048 491706 676076 492079
rect 675942 491671 675998 491680
rect 676036 491700 676088 491706
rect 675956 491434 675984 491671
rect 676036 491642 676088 491648
rect 676036 491564 676088 491570
rect 676036 491506 676088 491512
rect 675944 491428 675996 491434
rect 675944 491370 675996 491376
rect 676048 491337 676076 491506
rect 676034 491328 676090 491337
rect 676034 491263 676090 491272
rect 676034 490920 676090 490929
rect 676140 490906 676168 523942
rect 677510 504193 677538 524350
rect 677275 504165 677538 504193
rect 677275 503583 677303 504165
rect 677275 503555 677548 503583
rect 677520 491298 677548 503555
rect 676220 491292 676272 491298
rect 676220 491234 676272 491240
rect 677508 491292 677560 491298
rect 677508 491234 677560 491240
rect 676090 490878 676168 490906
rect 676034 490855 676090 490864
rect 675942 490512 675998 490521
rect 675942 490447 675998 490456
rect 675850 489288 675906 489297
rect 675850 489223 675906 489232
rect 675850 488880 675906 488889
rect 675850 488815 675906 488824
rect 675668 488572 675720 488578
rect 675720 488520 675800 488534
rect 675668 488514 675800 488520
rect 675680 488506 675800 488514
rect 675574 488472 675630 488481
rect 675574 488407 675630 488416
rect 674656 488232 674708 488238
rect 674656 488174 674708 488180
rect 675588 485858 675616 488407
rect 675668 487960 675720 487966
rect 675668 487902 675720 487908
rect 675680 486441 675708 487902
rect 675666 486432 675722 486441
rect 675666 486367 675722 486376
rect 675576 485852 675628 485858
rect 675576 485794 675628 485800
rect 674564 485784 674616 485790
rect 674564 485726 674616 485732
rect 674196 485512 674248 485518
rect 674196 485454 674248 485460
rect 674010 483576 674066 483585
rect 674010 483511 674066 483520
rect 673644 482996 673696 483002
rect 673644 482938 673696 482944
rect 673460 482928 673512 482934
rect 673460 482870 673512 482876
rect 675668 482928 675720 482934
rect 675668 482870 675720 482876
rect 675680 482769 675708 482870
rect 675666 482760 675722 482769
rect 675666 482695 675722 482704
rect 675772 411126 675800 488506
rect 675760 411120 675812 411126
rect 675760 411062 675812 411068
rect 675864 410938 675892 488815
rect 675956 488578 675984 490447
rect 676034 490104 676090 490113
rect 676232 490090 676260 491234
rect 676090 490062 676260 490090
rect 676034 490039 676090 490048
rect 676034 489696 676090 489705
rect 676090 489654 676168 489682
rect 676034 489631 676090 489640
rect 675944 488572 675996 488578
rect 675944 488514 675996 488520
rect 676036 488232 676088 488238
rect 676036 488174 676088 488180
rect 675942 488064 675998 488073
rect 675942 487999 675998 488008
rect 675956 478650 675984 487999
rect 676048 487257 676076 488174
rect 676034 487248 676090 487257
rect 676034 487183 676090 487192
rect 676036 487144 676088 487150
rect 676036 487086 676088 487092
rect 676048 486033 676076 487086
rect 676034 486024 676090 486033
rect 676034 485959 676090 485968
rect 676036 485784 676088 485790
rect 676036 485726 676088 485732
rect 676048 485625 676076 485726
rect 676034 485616 676090 485625
rect 676034 485551 676090 485560
rect 676036 485512 676088 485518
rect 676036 485454 676088 485460
rect 676048 483993 676076 485454
rect 676034 483984 676090 483993
rect 676034 483919 676090 483928
rect 676036 482996 676088 483002
rect 676036 482938 676088 482944
rect 676048 482361 676076 482938
rect 676034 482352 676090 482361
rect 676034 482287 676090 482296
rect 676034 481944 676090 481953
rect 676034 481879 676090 481888
rect 676048 480758 676076 481879
rect 676036 480752 676088 480758
rect 676034 480720 676036 480729
rect 676088 480720 676090 480729
rect 676034 480655 676090 480664
rect 676048 480629 676076 480655
rect 675944 478644 675996 478650
rect 675944 478586 675996 478592
rect 676140 478530 676168 489654
rect 675588 410910 675892 410938
rect 675956 478502 676168 478530
rect 675588 401033 675616 410910
rect 675956 410666 675984 478502
rect 676036 478440 676088 478446
rect 676036 478382 676088 478388
rect 675864 410638 675984 410666
rect 675758 402248 675814 402257
rect 675758 402183 675814 402192
rect 675666 401432 675722 401441
rect 675666 401367 675722 401376
rect 675574 401024 675630 401033
rect 675574 400959 675630 400968
rect 675116 400444 675168 400450
rect 675116 400386 675168 400392
rect 674380 399492 674432 399498
rect 674380 399434 674432 399440
rect 673828 397656 673880 397662
rect 673828 397598 673880 397604
rect 673460 396636 673512 396642
rect 673460 396578 673512 396584
rect 672908 392148 672960 392154
rect 672908 392090 672960 392096
rect 672816 278588 672868 278594
rect 672816 278530 672868 278536
rect 672816 256896 672868 256902
rect 672816 256838 672868 256844
rect 672722 148200 672778 148209
rect 672722 148135 672778 148144
rect 672448 130892 672500 130898
rect 672448 130834 672500 130840
rect 672354 116104 672410 116113
rect 672354 116039 672410 116048
rect 672262 109304 672318 109313
rect 672262 109239 672318 109248
rect 672460 105913 672488 130834
rect 672828 127945 672856 256838
rect 672920 143177 672948 392090
rect 673472 372094 673500 396578
rect 673552 395412 673604 395418
rect 673552 395354 673604 395360
rect 673564 376922 673592 395354
rect 673644 394868 673696 394874
rect 673644 394810 673696 394816
rect 673656 378146 673684 394810
rect 673736 392080 673788 392086
rect 673736 392022 673788 392028
rect 673644 378140 673696 378146
rect 673644 378082 673696 378088
rect 673748 376990 673776 392022
rect 673840 379506 673868 397598
rect 674288 397588 674340 397594
rect 674288 397530 674340 397536
rect 674012 392012 674064 392018
rect 674012 391954 674064 391960
rect 673828 379500 673880 379506
rect 673828 379442 673880 379448
rect 674024 378214 674052 391954
rect 674012 378208 674064 378214
rect 674012 378150 674064 378156
rect 673736 376984 673788 376990
rect 673736 376926 673788 376932
rect 673552 376916 673604 376922
rect 673552 376858 673604 376864
rect 674300 373930 674328 397530
rect 674392 383042 674420 399434
rect 674472 398268 674524 398274
rect 674472 398210 674524 398216
rect 674484 385014 674512 398210
rect 674656 397520 674708 397526
rect 674656 397462 674708 397468
rect 674564 390516 674616 390522
rect 674564 390458 674616 390464
rect 674472 385008 674524 385014
rect 674472 384950 674524 384956
rect 674380 383036 674432 383042
rect 674380 382978 674432 382984
rect 674288 373924 674340 373930
rect 674288 373866 674340 373872
rect 673460 372088 673512 372094
rect 673460 372030 673512 372036
rect 674576 370734 674604 390458
rect 674668 383178 674696 397462
rect 675024 395004 675076 395010
rect 675024 394946 675076 394952
rect 674932 394800 674984 394806
rect 674932 394742 674984 394748
rect 674748 390584 674800 390590
rect 674748 390526 674800 390532
rect 674656 383172 674708 383178
rect 674656 383114 674708 383120
rect 674656 383036 674708 383042
rect 674656 382978 674708 382984
rect 674564 370728 674616 370734
rect 674564 370670 674616 370676
rect 674668 361574 674696 382978
rect 674760 370802 674788 390526
rect 674944 381954 674972 394742
rect 675036 382498 675064 394946
rect 675024 382492 675076 382498
rect 675024 382434 675076 382440
rect 674932 381948 674984 381954
rect 674932 381890 674984 381896
rect 675128 374134 675156 400386
rect 675298 396944 675354 396953
rect 675298 396879 675354 396888
rect 675208 394732 675260 394738
rect 675208 394674 675260 394680
rect 675220 384130 675248 394674
rect 675312 385098 675340 396879
rect 675680 390522 675708 401367
rect 675772 390590 675800 402183
rect 675864 401849 675892 410638
rect 675944 403164 675996 403170
rect 675944 403106 675996 403112
rect 675956 403073 675984 403106
rect 675942 403064 675998 403073
rect 675942 402999 675998 403008
rect 675850 401840 675906 401849
rect 675850 401775 675906 401784
rect 676048 400217 676076 478382
rect 676128 411120 676180 411126
rect 676128 411062 676180 411068
rect 676140 402937 676168 411062
rect 676218 403744 676274 403753
rect 676218 403679 676274 403688
rect 676232 403442 676260 403679
rect 676220 403436 676272 403442
rect 676220 403378 676272 403384
rect 676218 403336 676274 403345
rect 676218 403271 676220 403280
rect 676272 403271 676274 403280
rect 676220 403242 676272 403248
rect 676126 402928 676182 402937
rect 676126 402863 676182 402872
rect 676126 400480 676182 400489
rect 676126 400415 676128 400424
rect 676180 400415 676182 400424
rect 676128 400386 676180 400392
rect 676034 400208 676090 400217
rect 676034 400143 676090 400152
rect 676034 399800 676090 399809
rect 676034 399735 676090 399744
rect 676048 399498 676076 399735
rect 676036 399492 676088 399498
rect 676036 399434 676088 399440
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675850 398576 675906 398585
rect 675850 398511 675906 398520
rect 675760 390584 675812 390590
rect 675760 390526 675812 390532
rect 675668 390516 675720 390522
rect 675668 390458 675720 390464
rect 675864 390402 675892 398511
rect 676048 398274 676076 399327
rect 676126 398848 676182 398857
rect 676126 398783 676182 398792
rect 676036 398268 676088 398274
rect 676036 398210 676088 398216
rect 676034 398168 676090 398177
rect 676034 398103 676090 398112
rect 675942 397760 675998 397769
rect 675942 397695 675998 397704
rect 675956 397662 675984 397695
rect 675944 397656 675996 397662
rect 675944 397598 675996 397604
rect 676048 397526 676076 398103
rect 676140 397594 676168 398783
rect 676128 397588 676180 397594
rect 676128 397530 676180 397536
rect 676036 397520 676088 397526
rect 676036 397462 676088 397468
rect 676034 397352 676090 397361
rect 676034 397287 676090 397296
rect 676048 396642 676076 397287
rect 676036 396636 676088 396642
rect 676036 396578 676088 396584
rect 676034 396536 676090 396545
rect 676034 396471 676090 396480
rect 675942 395720 675998 395729
rect 675942 395655 675998 395664
rect 675956 395418 675984 395655
rect 675944 395412 675996 395418
rect 675944 395354 675996 395360
rect 675942 395312 675998 395321
rect 675942 395247 675998 395256
rect 675956 394874 675984 395247
rect 676048 395010 676076 396471
rect 676126 395992 676182 396001
rect 676126 395927 676182 395936
rect 676036 395004 676088 395010
rect 676036 394946 676088 394952
rect 676034 394904 676090 394913
rect 675944 394868 675996 394874
rect 676034 394839 676090 394848
rect 675944 394810 675996 394816
rect 676048 394738 676076 394839
rect 676140 394806 676168 395927
rect 676128 394800 676180 394806
rect 676128 394742 676180 394748
rect 676036 394732 676088 394738
rect 676036 394674 676088 394680
rect 676034 394496 676090 394505
rect 676034 394431 676090 394440
rect 676048 392018 676076 394431
rect 676126 393952 676182 393961
rect 676126 393887 676182 393896
rect 676140 392086 676168 393887
rect 679070 393544 679126 393553
rect 679070 393479 679126 393488
rect 679084 392737 679112 393479
rect 679070 392728 679126 392737
rect 679070 392663 679126 392672
rect 679084 392154 679112 392663
rect 679072 392148 679124 392154
rect 679072 392090 679124 392096
rect 676128 392080 676180 392086
rect 676128 392022 676180 392028
rect 676036 392012 676088 392018
rect 676036 391954 676088 391960
rect 675772 390374 675892 390402
rect 675772 386442 675800 390374
rect 675760 386436 675812 386442
rect 675760 386378 675812 386384
rect 675760 386164 675812 386170
rect 675760 386106 675812 386112
rect 675772 385696 675800 386106
rect 675312 385070 675418 385098
rect 675300 385008 675352 385014
rect 675300 384950 675352 384956
rect 675312 384449 675340 384950
rect 675312 384421 675418 384449
rect 675208 384124 675260 384130
rect 675208 384066 675260 384072
rect 675300 383920 675352 383926
rect 675300 383862 675352 383868
rect 675312 380894 675340 383862
rect 675392 383172 675444 383178
rect 675392 383114 675444 383120
rect 675404 382568 675432 383114
rect 675392 382492 675444 382498
rect 675392 382434 675444 382440
rect 675404 382024 675432 382434
rect 675392 381948 675444 381954
rect 675392 381890 675444 381896
rect 675404 381412 675432 381890
rect 675312 380866 675432 380894
rect 675404 380732 675432 380866
rect 675300 379500 675352 379506
rect 675300 379442 675352 379448
rect 675312 378298 675340 379442
rect 675312 378270 675418 378298
rect 675484 378208 675536 378214
rect 675484 378150 675536 378156
rect 675300 378140 675352 378146
rect 675300 378082 675352 378088
rect 675312 377074 675340 378082
rect 675496 377740 675524 378150
rect 675312 377046 675418 377074
rect 675484 376984 675536 376990
rect 675484 376926 675536 376932
rect 675300 376916 675352 376922
rect 675300 376858 675352 376864
rect 675312 375238 675340 376858
rect 675496 376448 675524 376926
rect 675312 375210 675418 375238
rect 675116 374128 675168 374134
rect 675116 374070 675168 374076
rect 675300 374128 675352 374134
rect 675300 374070 675352 374076
rect 675312 372910 675340 374070
rect 675392 373924 675444 373930
rect 675392 373866 675444 373872
rect 675404 373388 675432 373866
rect 675300 372904 675352 372910
rect 675300 372846 675352 372852
rect 675300 372700 675352 372706
rect 675300 372642 675352 372648
rect 674748 370796 674800 370802
rect 674748 370738 674800 370744
rect 674668 361546 674788 361574
rect 673276 357060 673328 357066
rect 673276 357002 673328 357008
rect 673288 356114 673316 357002
rect 673368 356176 673420 356182
rect 673368 356118 673420 356124
rect 673000 356108 673052 356114
rect 673000 356050 673052 356056
rect 673276 356108 673328 356114
rect 673276 356050 673328 356056
rect 673012 351830 673040 356050
rect 673184 355428 673236 355434
rect 673184 355370 673236 355376
rect 673092 353524 673144 353530
rect 673092 353466 673144 353472
rect 673000 351824 673052 351830
rect 673000 351766 673052 351772
rect 673000 347268 673052 347274
rect 673000 347210 673052 347216
rect 672906 143168 672962 143177
rect 672906 143103 672962 143112
rect 673012 138145 673040 347210
rect 673104 310078 673132 353466
rect 673196 353394 673224 355370
rect 673276 354612 673328 354618
rect 673276 354554 673328 354560
rect 673288 353530 673316 354554
rect 673276 353524 673328 353530
rect 673276 353466 673328 353472
rect 673184 353388 673236 353394
rect 673184 353330 673236 353336
rect 673196 310894 673224 353330
rect 673276 351824 673328 351830
rect 673276 351766 673328 351772
rect 673288 312526 673316 351766
rect 673276 312520 673328 312526
rect 673276 312462 673328 312468
rect 673380 311710 673408 356118
rect 674760 355065 674788 361546
rect 675312 355881 675340 372642
rect 675392 372088 675444 372094
rect 675392 372030 675444 372036
rect 675404 371552 675432 372030
rect 675760 370796 675812 370802
rect 675760 370738 675812 370744
rect 675668 370728 675720 370734
rect 675668 370670 675720 370676
rect 675680 356697 675708 370670
rect 675772 357513 675800 370738
rect 675850 358728 675906 358737
rect 675850 358663 675906 358672
rect 675758 357504 675814 357513
rect 675758 357439 675814 357448
rect 675758 357096 675814 357105
rect 675758 357031 675760 357040
rect 675812 357031 675814 357040
rect 675760 357002 675812 357008
rect 675666 356688 675722 356697
rect 675666 356623 675722 356632
rect 675864 356250 675892 358663
rect 675942 358320 675998 358329
rect 675942 358255 675998 358264
rect 675956 356522 675984 358255
rect 676034 357912 676090 357921
rect 676034 357847 676090 357856
rect 675944 356516 675996 356522
rect 675944 356458 675996 356464
rect 676048 356386 676076 357847
rect 676036 356380 676088 356386
rect 676036 356322 676088 356328
rect 676034 356280 676090 356289
rect 675852 356244 675904 356250
rect 676034 356215 676090 356224
rect 675852 356186 675904 356192
rect 676048 356182 676076 356215
rect 676036 356176 676088 356182
rect 676036 356118 676088 356124
rect 675298 355872 675354 355881
rect 675298 355807 675354 355816
rect 676034 355464 676090 355473
rect 676034 355399 676036 355408
rect 676088 355399 676090 355408
rect 676036 355370 676088 355376
rect 674746 355056 674802 355065
rect 674746 354991 674802 355000
rect 676034 354648 676090 354657
rect 676034 354583 676036 354592
rect 676088 354583 676090 354592
rect 676036 354554 676088 354560
rect 676034 354240 676090 354249
rect 676034 354175 676090 354184
rect 676048 353530 676076 354175
rect 673828 353524 673880 353530
rect 673828 353466 673880 353472
rect 676036 353524 676088 353530
rect 676036 353466 676088 353472
rect 673460 351076 673512 351082
rect 673460 351018 673512 351024
rect 673472 333606 673500 351018
rect 673736 349852 673788 349858
rect 673736 349794 673788 349800
rect 673644 349036 673696 349042
rect 673644 348978 673696 348984
rect 673552 347880 673604 347886
rect 673552 347822 673604 347828
rect 673460 333600 673512 333606
rect 673460 333542 673512 333548
rect 673564 331634 673592 347822
rect 673656 332994 673684 348978
rect 673644 332988 673696 332994
rect 673644 332930 673696 332936
rect 673748 332450 673776 349794
rect 673840 339590 673868 353466
rect 676034 353424 676090 353433
rect 676034 353359 676090 353368
rect 676048 353326 676076 353359
rect 674104 353320 674156 353326
rect 674104 353262 674156 353268
rect 676036 353320 676088 353326
rect 676036 353262 676088 353268
rect 673920 350668 673972 350674
rect 673920 350610 673972 350616
rect 673828 339584 673880 339590
rect 673828 339526 673880 339532
rect 673932 336598 673960 350610
rect 674012 347812 674064 347818
rect 674012 347754 674064 347760
rect 673920 336592 673972 336598
rect 673920 336534 673972 336540
rect 674024 335918 674052 347754
rect 674116 341018 674144 353262
rect 676034 353016 676090 353025
rect 676034 352951 676090 352960
rect 675942 352608 675998 352617
rect 675942 352543 675998 352552
rect 675298 351792 675354 351801
rect 675298 351727 675354 351736
rect 674196 351484 674248 351490
rect 674196 351426 674248 351432
rect 674104 341012 674156 341018
rect 674104 340954 674156 340960
rect 674208 337958 674236 351426
rect 674288 350600 674340 350606
rect 674288 350542 674340 350548
rect 674196 337952 674248 337958
rect 674196 337894 674248 337900
rect 674300 337278 674328 350542
rect 675312 339878 675340 351727
rect 675956 351082 675984 352543
rect 676048 351490 676076 352951
rect 676036 351484 676088 351490
rect 676036 351426 676088 351432
rect 676034 351384 676090 351393
rect 676034 351319 676090 351328
rect 675944 351076 675996 351082
rect 675944 351018 675996 351024
rect 675942 350976 675998 350985
rect 675942 350911 675998 350920
rect 675956 350674 675984 350911
rect 675944 350668 675996 350674
rect 675944 350610 675996 350616
rect 676048 350606 676076 351319
rect 676036 350600 676088 350606
rect 676036 350542 676088 350548
rect 676034 350160 676090 350169
rect 676034 350095 676090 350104
rect 676048 349858 676076 350095
rect 676036 349852 676088 349858
rect 676036 349794 676088 349800
rect 676034 349752 676090 349761
rect 676034 349687 676090 349696
rect 675942 349344 675998 349353
rect 675942 349279 675998 349288
rect 675956 349042 675984 349279
rect 675944 349036 675996 349042
rect 675944 348978 675996 348984
rect 675942 348936 675998 348945
rect 675942 348871 675998 348880
rect 675956 347886 675984 348871
rect 675944 347880 675996 347886
rect 675944 347822 675996 347828
rect 676048 347818 676076 349687
rect 676036 347812 676088 347818
rect 676036 347754 676088 347760
rect 676034 347304 676090 347313
rect 676034 347239 676036 347248
rect 676088 347239 676090 347248
rect 676036 347210 676088 347216
rect 675484 341012 675536 341018
rect 675484 340954 675536 340960
rect 675496 340544 675524 340954
rect 675312 339850 675418 339878
rect 675484 339584 675536 339590
rect 675484 339526 675536 339532
rect 675496 339252 675524 339526
rect 675484 337952 675536 337958
rect 675484 337894 675536 337900
rect 675496 337416 675524 337894
rect 674288 337272 674340 337278
rect 674288 337214 674340 337220
rect 675392 337272 675444 337278
rect 675392 337214 675444 337220
rect 675404 336843 675432 337214
rect 675392 336592 675444 336598
rect 675392 336534 675444 336540
rect 675404 336192 675432 336534
rect 674012 335912 674064 335918
rect 674012 335854 674064 335860
rect 675484 335912 675536 335918
rect 675484 335854 675536 335860
rect 675496 335580 675524 335854
rect 675392 333600 675444 333606
rect 675392 333542 675444 333548
rect 675404 333064 675432 333542
rect 675392 332988 675444 332994
rect 675392 332930 675444 332936
rect 675404 332520 675432 332930
rect 673736 332444 673788 332450
rect 673736 332386 673788 332392
rect 675392 332444 675444 332450
rect 675392 332386 675444 332392
rect 675404 331875 675432 332386
rect 673552 331628 673604 331634
rect 673552 331570 673604 331576
rect 675392 331628 675444 331634
rect 675392 331570 675444 331576
rect 675404 331228 675432 331570
rect 675666 330576 675722 330585
rect 675666 330511 675722 330520
rect 675680 330035 675708 330511
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675758 326904 675814 326913
rect 675758 326839 675814 326848
rect 675772 326332 675800 326839
rect 676036 313744 676088 313750
rect 676034 313712 676036 313721
rect 676088 313712 676090 313721
rect 676034 313647 676090 313656
rect 676218 313168 676274 313177
rect 676218 313103 676274 313112
rect 676036 312928 676088 312934
rect 676034 312896 676036 312905
rect 676088 312896 676090 312905
rect 676034 312831 676090 312840
rect 676036 312520 676088 312526
rect 676034 312488 676036 312497
rect 676088 312488 676090 312497
rect 676034 312423 676090 312432
rect 676036 312112 676088 312118
rect 676034 312080 676036 312089
rect 676088 312080 676090 312089
rect 676232 312050 676260 313103
rect 676034 312015 676090 312024
rect 676220 312044 676272 312050
rect 676220 311986 676272 311992
rect 673368 311704 673420 311710
rect 676036 311704 676088 311710
rect 673368 311646 673420 311652
rect 676034 311672 676036 311681
rect 676088 311672 676090 311681
rect 676034 311607 676090 311616
rect 676034 311264 676090 311273
rect 676034 311199 676090 311208
rect 676048 311030 676076 311199
rect 674748 311024 674800 311030
rect 674748 310966 674800 310972
rect 676036 311024 676088 311030
rect 676036 310966 676088 310972
rect 673184 310888 673236 310894
rect 673184 310830 673236 310836
rect 673276 310480 673328 310486
rect 673276 310422 673328 310428
rect 673092 310072 673144 310078
rect 673092 310014 673144 310020
rect 673092 300892 673144 300898
rect 673092 300834 673144 300840
rect 672998 138136 673054 138145
rect 672998 138071 673054 138080
rect 673104 132977 673132 300834
rect 673288 266150 673316 310422
rect 674196 309188 674248 309194
rect 674196 309130 674248 309136
rect 673552 308100 673604 308106
rect 673552 308042 673604 308048
rect 673460 306536 673512 306542
rect 673460 306478 673512 306484
rect 673472 281926 673500 306478
rect 673564 283762 673592 308042
rect 673920 306400 673972 306406
rect 673920 306342 673972 306348
rect 673644 305108 673696 305114
rect 673644 305050 673696 305056
rect 673656 285598 673684 305050
rect 673736 304700 673788 304706
rect 673736 304642 673788 304648
rect 673748 287230 673776 304642
rect 673828 303884 673880 303890
rect 673828 303826 673880 303832
rect 673736 287224 673788 287230
rect 673736 287166 673788 287172
rect 673840 286618 673868 303826
rect 673932 288590 673960 306342
rect 674012 303816 674064 303822
rect 674012 303758 674064 303764
rect 673920 288584 673972 288590
rect 673920 288526 673972 288532
rect 674024 287978 674052 303758
rect 674208 294574 674236 309130
rect 674472 306468 674524 306474
rect 674472 306410 674524 306416
rect 674196 294568 674248 294574
rect 674196 294510 674248 294516
rect 674484 292942 674512 306410
rect 674656 306060 674708 306066
rect 674656 306002 674708 306008
rect 674564 303748 674616 303754
rect 674564 303690 674616 303696
rect 674472 292936 674524 292942
rect 674472 292878 674524 292884
rect 674576 291106 674604 303690
rect 674668 292330 674696 306002
rect 674656 292324 674708 292330
rect 674656 292266 674708 292272
rect 674564 291100 674616 291106
rect 674564 291042 674616 291048
rect 674012 287972 674064 287978
rect 674012 287914 674064 287920
rect 673828 286612 673880 286618
rect 673828 286554 673880 286560
rect 673644 285592 673696 285598
rect 673644 285534 673696 285540
rect 673552 283756 673604 283762
rect 673552 283698 673604 283704
rect 673460 281920 673512 281926
rect 673460 281862 673512 281868
rect 674760 267714 674788 310966
rect 676036 310888 676088 310894
rect 676034 310856 676036 310865
rect 676088 310856 676090 310865
rect 676034 310791 676090 310800
rect 676036 310480 676088 310486
rect 676034 310448 676036 310457
rect 676088 310448 676090 310457
rect 676034 310383 676090 310392
rect 676036 310072 676088 310078
rect 676034 310040 676036 310049
rect 676088 310040 676090 310049
rect 676034 309975 676090 309984
rect 676036 309664 676088 309670
rect 676034 309632 676036 309641
rect 676088 309632 676090 309641
rect 676034 309567 676090 309576
rect 676034 309224 676090 309233
rect 676034 309159 676036 309168
rect 676088 309159 676090 309168
rect 676036 309130 676088 309136
rect 676034 308816 676090 308825
rect 676034 308751 676090 308760
rect 675758 308408 675814 308417
rect 675758 308343 675814 308352
rect 675482 306776 675538 306785
rect 675482 306711 675538 306720
rect 675496 301034 675524 306711
rect 675208 301028 675260 301034
rect 675208 300970 675260 300976
rect 675484 301028 675536 301034
rect 675484 300970 675536 300976
rect 675220 295118 675248 300970
rect 675772 296206 675800 308343
rect 676048 308106 676076 308751
rect 676036 308100 676088 308106
rect 676036 308042 676088 308048
rect 676034 308000 676090 308009
rect 676034 307935 676090 307944
rect 675942 307184 675998 307193
rect 675942 307119 675998 307128
rect 675956 306542 675984 307119
rect 675944 306536 675996 306542
rect 675944 306478 675996 306484
rect 676048 306474 676076 307935
rect 676126 307456 676182 307465
rect 676126 307391 676182 307400
rect 676036 306468 676088 306474
rect 676036 306410 676088 306416
rect 676140 306406 676168 307391
rect 676128 306400 676180 306406
rect 676034 306368 676090 306377
rect 676128 306342 676180 306348
rect 676034 306303 676090 306312
rect 676048 306066 676076 306303
rect 676036 306060 676088 306066
rect 676036 306002 676088 306008
rect 676126 305416 676182 305425
rect 676126 305351 676182 305360
rect 676140 305114 676168 305351
rect 676128 305108 676180 305114
rect 676128 305050 676180 305056
rect 676126 305008 676182 305017
rect 676126 304943 676182 304952
rect 676140 304706 676168 304943
rect 676128 304700 676180 304706
rect 676128 304642 676180 304648
rect 676126 304600 676182 304609
rect 676126 304535 676182 304544
rect 675942 304328 675998 304337
rect 675942 304263 675998 304272
rect 675850 303920 675906 303929
rect 675850 303855 675852 303864
rect 675904 303855 675906 303864
rect 675852 303826 675904 303832
rect 675956 303822 675984 304263
rect 675944 303816 675996 303822
rect 675944 303758 675996 303764
rect 676140 303754 676168 304535
rect 676128 303748 676180 303754
rect 676128 303690 676180 303696
rect 678978 303376 679034 303385
rect 678978 303311 679034 303320
rect 678992 302569 679020 303311
rect 678978 302560 679034 302569
rect 678978 302495 679034 302504
rect 678992 300898 679020 302495
rect 678980 300892 679032 300898
rect 678980 300834 679032 300840
rect 675760 296200 675812 296206
rect 675760 296142 675812 296148
rect 675760 295996 675812 296002
rect 675760 295938 675812 295944
rect 675772 295528 675800 295938
rect 675208 295112 675260 295118
rect 675208 295054 675260 295060
rect 675392 295112 675444 295118
rect 675392 295054 675444 295060
rect 675404 294879 675432 295054
rect 675392 294568 675444 294574
rect 675392 294510 675444 294516
rect 675404 294236 675432 294510
rect 675392 292936 675444 292942
rect 675392 292878 675444 292884
rect 675404 292400 675432 292878
rect 675392 292324 675444 292330
rect 675392 292266 675444 292272
rect 675404 291856 675432 292266
rect 675758 291680 675814 291689
rect 675758 291615 675814 291624
rect 675772 291176 675800 291615
rect 675392 291100 675444 291106
rect 675392 291042 675444 291048
rect 675404 290564 675432 291042
rect 675392 288584 675444 288590
rect 675392 288526 675444 288532
rect 675404 288048 675432 288526
rect 675392 287972 675444 287978
rect 675392 287914 675444 287920
rect 675404 287504 675432 287914
rect 675484 287224 675536 287230
rect 675484 287166 675536 287172
rect 675496 286892 675524 287166
rect 675392 286612 675444 286618
rect 675392 286554 675444 286560
rect 675404 286212 675432 286554
rect 675484 285592 675536 285598
rect 675484 285534 675536 285540
rect 675496 285056 675524 285534
rect 675484 283756 675536 283762
rect 675484 283698 675536 283704
rect 675496 283220 675524 283698
rect 675392 281920 675444 281926
rect 675392 281862 675444 281868
rect 675404 281355 675432 281862
rect 676126 268560 676182 268569
rect 676126 268495 676182 268504
rect 676036 267980 676088 267986
rect 676036 267922 676088 267928
rect 676048 267889 676076 267922
rect 676034 267880 676090 267889
rect 676034 267815 676090 267824
rect 676140 267782 676168 268495
rect 676218 268152 676274 268161
rect 676218 268087 676220 268096
rect 676272 268087 676274 268096
rect 676220 268058 676272 268064
rect 676128 267776 676180 267782
rect 676128 267718 676180 267724
rect 674748 267708 674800 267714
rect 674748 267650 674800 267656
rect 676036 267708 676088 267714
rect 676036 267650 676088 267656
rect 675944 267504 675996 267510
rect 675942 267472 675944 267481
rect 675996 267472 675998 267481
rect 675942 267407 675998 267416
rect 675758 267064 675814 267073
rect 675758 266999 675814 267008
rect 675668 266348 675720 266354
rect 675668 266290 675720 266296
rect 673276 266144 673328 266150
rect 673276 266086 673328 266092
rect 675680 265441 675708 266290
rect 675666 265432 675722 265441
rect 674748 265396 674800 265402
rect 675666 265367 675722 265376
rect 674748 265338 674800 265344
rect 674760 264974 674788 265338
rect 674576 264946 674788 264974
rect 674196 263084 674248 263090
rect 674196 263026 674248 263032
rect 674012 262540 674064 262546
rect 674012 262482 674064 262488
rect 673736 262336 673788 262342
rect 673736 262278 673788 262284
rect 673460 260228 673512 260234
rect 673460 260170 673512 260176
rect 673472 240582 673500 260170
rect 673552 259752 673604 259758
rect 673552 259694 673604 259700
rect 673564 242214 673592 259694
rect 673644 256828 673696 256834
rect 673644 256770 673696 256776
rect 673552 242208 673604 242214
rect 673552 242150 673604 242156
rect 673656 241602 673684 256770
rect 673748 243642 673776 262278
rect 673828 256760 673880 256766
rect 673828 256702 673880 256708
rect 673736 243636 673788 243642
rect 673736 243578 673788 243584
rect 673840 242962 673868 256702
rect 674024 245654 674052 262482
rect 674104 261860 674156 261866
rect 674104 261802 674156 261808
rect 674116 246378 674144 261802
rect 674208 249626 674236 263026
rect 674288 262268 674340 262274
rect 674288 262210 674340 262216
rect 674196 249620 674248 249626
rect 674196 249562 674248 249568
rect 674300 247926 674328 262210
rect 674472 259684 674524 259690
rect 674472 259626 674524 259632
rect 674380 259616 674432 259622
rect 674380 259558 674432 259564
rect 674288 247920 674340 247926
rect 674288 247862 674340 247868
rect 674392 246566 674420 259558
rect 674484 247314 674512 259626
rect 674472 247308 674524 247314
rect 674472 247250 674524 247256
rect 674380 246560 674432 246566
rect 674380 246502 674432 246508
rect 674116 246350 674512 246378
rect 674024 245626 674420 245654
rect 673828 242956 673880 242962
rect 673828 242898 673880 242904
rect 674392 241942 674420 245626
rect 674380 241936 674432 241942
rect 674380 241878 674432 241884
rect 673644 241596 673696 241602
rect 673644 241538 673696 241544
rect 673460 240576 673512 240582
rect 673460 240518 673512 240524
rect 674484 236910 674512 246350
rect 674472 236904 674524 236910
rect 674472 236846 674524 236852
rect 674576 223582 674604 264946
rect 675574 260536 675630 260545
rect 675574 260471 675630 260480
rect 675588 260234 675616 260471
rect 675576 260228 675628 260234
rect 675576 260170 675628 260176
rect 675574 260128 675630 260137
rect 675574 260063 675630 260072
rect 675588 259758 675616 260063
rect 675576 259752 675628 259758
rect 675576 259694 675628 259700
rect 675024 259548 675076 259554
rect 675024 259490 675076 259496
rect 674748 255332 674800 255338
rect 674748 255274 674800 255280
rect 674656 255264 674708 255270
rect 674656 255206 674708 255212
rect 674668 235550 674696 255206
rect 674760 235618 674788 255274
rect 675036 247602 675064 259490
rect 675208 259480 675260 259486
rect 675208 259422 675260 259428
rect 675220 250442 675248 259422
rect 675680 255338 675708 265367
rect 675772 265062 675800 266999
rect 676048 266665 676076 267650
rect 676034 266656 676090 266665
rect 676034 266591 676090 266600
rect 676034 266248 676090 266257
rect 676034 266183 676090 266192
rect 676048 265402 676076 266183
rect 676220 266144 676272 266150
rect 676218 266112 676220 266121
rect 676272 266112 676274 266121
rect 676218 266047 676274 266056
rect 676036 265396 676088 265402
rect 676036 265338 676088 265344
rect 675760 265056 675812 265062
rect 675760 264998 675812 265004
rect 675668 255332 675720 255338
rect 675668 255274 675720 255280
rect 675772 255270 675800 264998
rect 676220 264988 676272 264994
rect 676220 264930 676272 264936
rect 676232 264897 676260 264930
rect 676218 264888 676274 264897
rect 676218 264823 676274 264832
rect 676034 264208 676090 264217
rect 676034 264143 676090 264152
rect 675850 263392 675906 263401
rect 675850 263327 675906 263336
rect 675760 255264 675812 255270
rect 675760 255206 675812 255212
rect 675864 255082 675892 263327
rect 676048 263090 676076 264143
rect 676126 263664 676182 263673
rect 676126 263599 676182 263608
rect 676036 263084 676088 263090
rect 676036 263026 676088 263032
rect 676034 262984 676090 262993
rect 676034 262919 676090 262928
rect 676048 262274 676076 262919
rect 676140 262546 676168 263599
rect 676128 262540 676180 262546
rect 676128 262482 676180 262488
rect 676126 262440 676182 262449
rect 676126 262375 676182 262384
rect 676140 262342 676168 262375
rect 676128 262336 676180 262342
rect 676128 262278 676180 262284
rect 676036 262268 676088 262274
rect 676036 262210 676088 262216
rect 676034 262168 676090 262177
rect 676034 262103 676090 262112
rect 676048 261866 676076 262103
rect 676036 261860 676088 261866
rect 676036 261802 676088 261808
rect 676034 261760 676090 261769
rect 676034 261695 676090 261704
rect 675942 260944 675998 260953
rect 675942 260879 675998 260888
rect 675956 259622 675984 260879
rect 675944 259616 675996 259622
rect 675944 259558 675996 259564
rect 676048 259486 676076 261695
rect 676126 261216 676182 261225
rect 676126 261151 676182 261160
rect 676140 259690 676168 261151
rect 676128 259684 676180 259690
rect 676128 259626 676180 259632
rect 676126 259584 676182 259593
rect 676126 259519 676128 259528
rect 676180 259519 676182 259528
rect 676128 259490 676180 259496
rect 676036 259480 676088 259486
rect 676036 259422 676088 259428
rect 676034 259312 676090 259321
rect 676034 259247 676090 259256
rect 676048 256766 676076 259247
rect 676126 258768 676182 258777
rect 676126 258703 676182 258712
rect 676140 256834 676168 258703
rect 678978 258360 679034 258369
rect 678978 258295 679034 258304
rect 678992 257553 679020 258295
rect 678978 257544 679034 257553
rect 678978 257479 679034 257488
rect 678992 256902 679020 257479
rect 678980 256896 679032 256902
rect 678980 256838 679032 256844
rect 676128 256828 676180 256834
rect 676128 256770 676180 256776
rect 676036 256760 676088 256766
rect 676036 256702 676088 256708
rect 675772 255054 675892 255082
rect 675772 251258 675800 255054
rect 675760 251252 675812 251258
rect 675760 251194 675812 251200
rect 675760 250980 675812 250986
rect 675760 250922 675812 250928
rect 675772 250512 675800 250922
rect 675208 250436 675260 250442
rect 675208 250378 675260 250384
rect 675484 250436 675536 250442
rect 675484 250378 675536 250384
rect 675496 249900 675524 250378
rect 675392 249620 675444 249626
rect 675392 249562 675444 249568
rect 675404 249220 675432 249562
rect 675484 247920 675536 247926
rect 675484 247862 675536 247868
rect 675036 247574 675156 247602
rect 675128 246090 675156 247574
rect 675496 247384 675524 247862
rect 675392 247308 675444 247314
rect 675392 247250 675444 247256
rect 675404 246840 675432 247250
rect 675392 246560 675444 246566
rect 675392 246502 675444 246508
rect 675404 246199 675432 246502
rect 675116 246084 675168 246090
rect 675116 246026 675168 246032
rect 675392 246084 675444 246090
rect 675392 246026 675444 246032
rect 675404 245548 675432 246026
rect 675300 243636 675352 243642
rect 675300 243578 675352 243584
rect 675312 243085 675340 243578
rect 675312 243057 675418 243085
rect 675300 242956 675352 242962
rect 675300 242898 675352 242904
rect 675312 242533 675340 242898
rect 675312 242505 675418 242533
rect 675392 242208 675444 242214
rect 675392 242150 675444 242156
rect 675300 241936 675352 241942
rect 675300 241878 675352 241884
rect 675312 238218 675340 241878
rect 675404 241876 675432 242150
rect 675392 241596 675444 241602
rect 675392 241538 675444 241544
rect 675404 241231 675432 241538
rect 675392 240576 675444 240582
rect 675392 240518 675444 240524
rect 675404 240040 675432 240518
rect 675312 238190 675418 238218
rect 675392 236904 675444 236910
rect 675392 236846 675444 236852
rect 675404 236368 675432 236846
rect 674748 235612 674800 235618
rect 674748 235554 674800 235560
rect 675668 235612 675720 235618
rect 675668 235554 675720 235560
rect 674656 235544 674708 235550
rect 674656 235486 674708 235492
rect 675680 226334 675708 235554
rect 675760 235544 675812 235550
rect 675760 235486 675812 235492
rect 675588 226306 675708 226334
rect 674564 223576 674616 223582
rect 674564 223518 674616 223524
rect 674656 222216 674708 222222
rect 674656 222158 674708 222164
rect 674104 218340 674156 218346
rect 674104 218282 674156 218288
rect 673460 218136 673512 218142
rect 673460 218078 673512 218084
rect 673184 212084 673236 212090
rect 673184 212026 673236 212032
rect 673090 132968 673146 132977
rect 673090 132903 673146 132912
rect 672814 127936 672870 127945
rect 672814 127871 672870 127880
rect 672908 123140 672960 123146
rect 672908 123082 672960 123088
rect 672920 112713 672948 123082
rect 673196 122913 673224 212026
rect 673472 193526 673500 218078
rect 673644 217116 673696 217122
rect 673644 217058 673696 217064
rect 673552 216300 673604 216306
rect 673552 216242 673604 216248
rect 673460 193520 673512 193526
rect 673460 193462 673512 193468
rect 673564 191690 673592 216242
rect 673656 198422 673684 217058
rect 673920 215484 673972 215490
rect 673920 215426 673972 215432
rect 673828 214668 673880 214674
rect 673828 214610 673880 214616
rect 673736 212628 673788 212634
rect 673736 212570 673788 212576
rect 673644 198416 673696 198422
rect 673644 198358 673696 198364
rect 673748 197606 673776 212570
rect 673736 197600 673788 197606
rect 673736 197542 673788 197548
rect 673840 197062 673868 214610
rect 673932 201550 673960 215426
rect 674012 213852 674064 213858
rect 674012 213794 674064 213800
rect 673920 201544 673972 201550
rect 673920 201486 673972 201492
rect 674024 200734 674052 213794
rect 674116 204610 674144 218282
rect 674380 218068 674432 218074
rect 674380 218010 674432 218016
rect 674196 216708 674248 216714
rect 674196 216650 674248 216656
rect 674104 204604 674156 204610
rect 674104 204546 674156 204552
rect 674208 202774 674236 216650
rect 674288 215416 674340 215422
rect 674288 215358 674340 215364
rect 674196 202768 674248 202774
rect 674196 202710 674248 202716
rect 674300 201890 674328 215358
rect 674392 205562 674420 218010
rect 674472 215348 674524 215354
rect 674472 215290 674524 215296
rect 674380 205556 674432 205562
rect 674380 205498 674432 205504
rect 674380 205420 674432 205426
rect 674380 205362 674432 205368
rect 674288 201884 674340 201890
rect 674288 201826 674340 201832
rect 674012 200728 674064 200734
rect 674012 200670 674064 200676
rect 673828 197056 673880 197062
rect 673828 196998 673880 197004
rect 674392 195226 674420 205362
rect 674484 205222 674512 215290
rect 674564 206168 674616 206174
rect 674564 206110 674616 206116
rect 674472 205216 674524 205222
rect 674472 205158 674524 205164
rect 674470 205048 674526 205057
rect 674470 204983 674526 204992
rect 674484 196450 674512 204983
rect 674472 196444 674524 196450
rect 674472 196386 674524 196392
rect 674380 195220 674432 195226
rect 674380 195162 674432 195168
rect 673552 191684 673604 191690
rect 673552 191626 673604 191632
rect 673276 176928 673328 176934
rect 673276 176870 673328 176876
rect 673288 132326 673316 176870
rect 673368 176044 673420 176050
rect 673368 175986 673420 175992
rect 673276 132320 673328 132326
rect 673276 132262 673328 132268
rect 673380 131510 673408 175986
rect 674576 175574 674604 206110
rect 674668 205850 674696 222158
rect 675588 220697 675616 226306
rect 675666 223136 675722 223145
rect 675666 223071 675722 223080
rect 675680 220862 675708 223071
rect 675772 222329 675800 235486
rect 675852 223576 675904 223582
rect 675852 223518 675904 223524
rect 675942 223544 675998 223553
rect 675758 222320 675814 222329
rect 675758 222255 675814 222264
rect 675760 222216 675812 222222
rect 675760 222158 675812 222164
rect 675772 221921 675800 222158
rect 675758 221912 675814 221921
rect 675758 221847 675814 221856
rect 675864 221513 675892 223518
rect 675942 223479 675998 223488
rect 675850 221504 675906 221513
rect 675850 221439 675906 221448
rect 675956 221202 675984 223479
rect 676034 222728 676090 222737
rect 676034 222663 676090 222672
rect 675944 221196 675996 221202
rect 675944 221138 675996 221144
rect 675758 221096 675814 221105
rect 676048 221066 676076 222663
rect 675758 221031 675814 221040
rect 676036 221060 676088 221066
rect 675668 220856 675720 220862
rect 675668 220798 675720 220804
rect 675574 220688 675630 220697
rect 675574 220623 675630 220632
rect 675576 219564 675628 219570
rect 675576 219506 675628 219512
rect 674840 219360 674892 219366
rect 674840 219302 674892 219308
rect 674852 206174 674880 219302
rect 675390 215384 675446 215393
rect 675390 215319 675446 215328
rect 675208 212560 675260 212566
rect 675208 212502 675260 212508
rect 674840 206168 674892 206174
rect 674840 206110 674892 206116
rect 674840 206032 674892 206038
rect 674840 205974 674892 205980
rect 674668 205822 674788 205850
rect 674656 205760 674708 205766
rect 674656 205702 674708 205708
rect 674668 196586 674696 205702
rect 674656 196580 674708 196586
rect 674656 196522 674708 196528
rect 674656 196444 674708 196450
rect 674656 196386 674708 196392
rect 674668 176390 674696 196386
rect 674760 179382 674788 205822
rect 674852 195362 674880 205974
rect 675220 205766 675248 212502
rect 675404 206038 675432 215319
rect 675392 206032 675444 206038
rect 675588 206009 675616 219506
rect 675772 206038 675800 221031
rect 676036 221002 676088 221008
rect 676034 220280 676090 220289
rect 676034 220215 676090 220224
rect 676048 219570 676076 220215
rect 676036 219564 676088 219570
rect 676036 219506 676088 219512
rect 676034 219464 676090 219473
rect 676034 219399 676090 219408
rect 676048 219366 676076 219399
rect 676036 219360 676088 219366
rect 676036 219302 676088 219308
rect 676034 219056 676090 219065
rect 676034 218991 676090 219000
rect 675942 218648 675998 218657
rect 675942 218583 675998 218592
rect 675956 218142 675984 218583
rect 676048 218346 676076 218991
rect 676036 218340 676088 218346
rect 676036 218282 676088 218288
rect 676034 218240 676090 218249
rect 676034 218175 676090 218184
rect 675944 218136 675996 218142
rect 675944 218078 675996 218084
rect 676048 218074 676076 218175
rect 676036 218068 676088 218074
rect 676036 218010 676088 218016
rect 676034 217832 676090 217841
rect 676034 217767 676090 217776
rect 675942 217424 675998 217433
rect 675942 217359 675998 217368
rect 675956 217122 675984 217359
rect 675944 217116 675996 217122
rect 675944 217058 675996 217064
rect 675942 217016 675998 217025
rect 675942 216951 675998 216960
rect 675956 216306 675984 216951
rect 676048 216714 676076 217767
rect 676036 216708 676088 216714
rect 676036 216650 676088 216656
rect 676034 216608 676090 216617
rect 676034 216543 676090 216552
rect 675944 216300 675996 216306
rect 675944 216242 675996 216248
rect 675942 216200 675998 216209
rect 675942 216135 675998 216144
rect 675850 215792 675906 215801
rect 675850 215727 675906 215736
rect 675864 215490 675892 215727
rect 675852 215484 675904 215490
rect 675852 215426 675904 215432
rect 675956 215422 675984 216135
rect 675944 215416 675996 215422
rect 675944 215358 675996 215364
rect 676048 215354 676076 216543
rect 676036 215348 676088 215354
rect 676036 215290 676088 215296
rect 676034 214976 676090 214985
rect 676034 214911 676090 214920
rect 676048 214674 676076 214911
rect 676036 214668 676088 214674
rect 676036 214610 676088 214616
rect 676034 214568 676090 214577
rect 676034 214503 676090 214512
rect 675942 214160 675998 214169
rect 675942 214095 675998 214104
rect 675956 212634 675984 214095
rect 676048 213858 676076 214503
rect 676036 213852 676088 213858
rect 676036 213794 676088 213800
rect 676034 213752 676090 213761
rect 676034 213687 676090 213696
rect 675944 212628 675996 212634
rect 675944 212570 675996 212576
rect 676048 212566 676076 213687
rect 676036 212560 676088 212566
rect 676036 212502 676088 212508
rect 676034 212120 676090 212129
rect 676034 212055 676036 212064
rect 676088 212055 676090 212064
rect 676036 212026 676088 212032
rect 675760 206032 675812 206038
rect 675392 205974 675444 205980
rect 675574 206000 675630 206009
rect 675760 205974 675812 205980
rect 675574 205935 675630 205944
rect 675208 205760 675260 205766
rect 675208 205702 675260 205708
rect 675300 205556 675352 205562
rect 675300 205498 675352 205504
rect 675312 205337 675340 205498
rect 675312 205309 675418 205337
rect 675300 205216 675352 205222
rect 675300 205158 675352 205164
rect 675312 204694 675340 205158
rect 675312 204666 675418 204694
rect 675300 204604 675352 204610
rect 675300 204546 675352 204552
rect 675312 204049 675340 204546
rect 675312 204021 675418 204049
rect 675484 202768 675536 202774
rect 675484 202710 675536 202716
rect 675496 202195 675524 202710
rect 675392 201884 675444 201890
rect 675392 201826 675444 201832
rect 675404 201620 675432 201826
rect 675392 201544 675444 201550
rect 675392 201486 675444 201492
rect 675404 201008 675432 201486
rect 675392 200728 675444 200734
rect 675392 200670 675444 200676
rect 675404 200328 675432 200670
rect 675392 198416 675444 198422
rect 675392 198358 675444 198364
rect 675404 197880 675432 198358
rect 675484 197600 675536 197606
rect 675484 197542 675536 197548
rect 675496 197336 675524 197542
rect 675392 197056 675444 197062
rect 675392 196998 675444 197004
rect 675404 196656 675432 196998
rect 675392 196580 675444 196586
rect 675392 196522 675444 196528
rect 675404 196044 675432 196522
rect 674840 195356 674892 195362
rect 674840 195298 674892 195304
rect 675392 195356 675444 195362
rect 675392 195298 675444 195304
rect 674840 195220 674892 195226
rect 674840 195162 674892 195168
rect 674748 179376 674800 179382
rect 674748 179318 674800 179324
rect 674852 176662 674880 195162
rect 675404 194820 675432 195298
rect 675392 193520 675444 193526
rect 675392 193462 675444 193468
rect 675404 192984 675432 193462
rect 675392 191684 675444 191690
rect 675392 191626 675444 191632
rect 675404 191148 675432 191626
rect 675852 179376 675904 179382
rect 675852 179318 675904 179324
rect 675758 178528 675814 178537
rect 675758 178463 675814 178472
rect 675772 176866 675800 178463
rect 675864 177313 675892 179318
rect 675942 178120 675998 178129
rect 675942 178055 675998 178064
rect 675850 177304 675906 177313
rect 675850 177239 675906 177248
rect 675956 177138 675984 178055
rect 676034 177712 676090 177721
rect 676034 177647 676090 177656
rect 675944 177132 675996 177138
rect 675944 177074 675996 177080
rect 676048 177002 676076 177647
rect 676036 176996 676088 177002
rect 676036 176938 676088 176944
rect 675944 176928 675996 176934
rect 675942 176896 675944 176905
rect 675996 176896 675998 176905
rect 675760 176860 675812 176866
rect 675942 176831 675998 176840
rect 675760 176802 675812 176808
rect 674840 176656 674892 176662
rect 674840 176598 674892 176604
rect 676036 176656 676088 176662
rect 676036 176598 676088 176604
rect 676048 176497 676076 176598
rect 676034 176488 676090 176497
rect 676034 176423 676090 176432
rect 674656 176384 674708 176390
rect 674656 176326 674708 176332
rect 676036 176384 676088 176390
rect 676036 176326 676088 176332
rect 675942 176080 675998 176089
rect 675942 176015 675944 176024
rect 675996 176015 675998 176024
rect 675944 175986 675996 175992
rect 676048 175681 676076 176326
rect 676034 175672 676090 175681
rect 676034 175607 676090 175616
rect 674564 175568 674616 175574
rect 674564 175510 674616 175516
rect 676036 175568 676088 175574
rect 676036 175510 676088 175516
rect 675944 175296 675996 175302
rect 675942 175264 675944 175273
rect 675996 175264 675998 175273
rect 675942 175199 675998 175208
rect 676048 174865 676076 175510
rect 676034 174856 676090 174865
rect 676034 174791 676090 174800
rect 676036 174480 676088 174486
rect 676034 174448 676036 174457
rect 676088 174448 676090 174457
rect 676034 174383 676090 174392
rect 676034 174040 676090 174049
rect 676034 173975 676090 173984
rect 676048 173942 676076 173975
rect 674104 173936 674156 173942
rect 674104 173878 674156 173884
rect 676036 173936 676088 173942
rect 676036 173878 676088 173884
rect 673736 171352 673788 171358
rect 673736 171294 673788 171300
rect 673460 170060 673512 170066
rect 673460 170002 673512 170008
rect 673472 150414 673500 170002
rect 673644 169244 673696 169250
rect 673644 169186 673696 169192
rect 673552 168564 673604 168570
rect 673552 168506 673604 168512
rect 673564 151434 673592 168506
rect 673656 152046 673684 169186
rect 673748 153406 673776 171294
rect 673828 168768 673880 168774
rect 673828 168710 673880 168716
rect 673736 153400 673788 153406
rect 673736 153342 673788 153348
rect 673840 152590 673868 168710
rect 674116 159390 674144 173878
rect 675758 173224 675814 173233
rect 675758 173159 675814 173168
rect 674656 171692 674708 171698
rect 674656 171634 674708 171640
rect 674564 171216 674616 171222
rect 674564 171158 674616 171164
rect 674104 159384 674156 159390
rect 674104 159326 674156 159332
rect 674576 156942 674604 171158
rect 674668 157758 674696 171634
rect 674840 171148 674892 171154
rect 674840 171090 674892 171096
rect 674748 168700 674800 168706
rect 674748 168642 674800 168648
rect 674656 157752 674708 157758
rect 674656 157694 674708 157700
rect 674564 156936 674616 156942
rect 674564 156878 674616 156884
rect 674760 155718 674788 168642
rect 674852 159934 674880 171090
rect 675772 161022 675800 173159
rect 676034 172816 676090 172825
rect 676034 172751 676090 172760
rect 675942 172408 675998 172417
rect 675942 172343 675998 172352
rect 675956 171358 675984 172343
rect 676048 171698 676076 172751
rect 676036 171692 676088 171698
rect 676036 171634 676088 171640
rect 676034 171592 676090 171601
rect 676034 171527 676090 171536
rect 675944 171352 675996 171358
rect 675944 171294 675996 171300
rect 675944 171216 675996 171222
rect 675942 171184 675944 171193
rect 675996 171184 675998 171193
rect 676048 171154 676076 171527
rect 675942 171119 675998 171128
rect 676036 171148 676088 171154
rect 676036 171090 676088 171096
rect 675942 170368 675998 170377
rect 675942 170303 675998 170312
rect 675956 170066 675984 170303
rect 675944 170060 675996 170066
rect 675944 170002 675996 170008
rect 675942 169960 675998 169969
rect 675942 169895 675998 169904
rect 675956 169250 675984 169895
rect 676034 169552 676090 169561
rect 676034 169487 676090 169496
rect 675944 169244 675996 169250
rect 675944 169186 675996 169192
rect 675942 169144 675998 169153
rect 675942 169079 675998 169088
rect 675956 168774 675984 169079
rect 675944 168768 675996 168774
rect 675850 168736 675906 168745
rect 675944 168710 675996 168716
rect 676048 168706 676076 169487
rect 675850 168671 675906 168680
rect 676036 168700 676088 168706
rect 675864 168570 675892 168671
rect 676036 168642 676088 168648
rect 675852 168564 675904 168570
rect 675852 168506 675904 168512
rect 676034 168328 676090 168337
rect 676034 168263 676036 168272
rect 676088 168263 676090 168272
rect 676036 168234 676088 168240
rect 676034 167920 676090 167929
rect 676034 167855 676036 167864
rect 676088 167855 676090 167864
rect 676036 167826 676088 167832
rect 676034 167104 676090 167113
rect 676034 167039 676036 167048
rect 676088 167039 676090 167048
rect 676036 167010 676088 167016
rect 675760 161016 675812 161022
rect 675760 160958 675812 160964
rect 675760 160812 675812 160818
rect 675760 160754 675812 160760
rect 675772 160344 675800 160754
rect 674840 159928 674892 159934
rect 674840 159870 674892 159876
rect 675392 159928 675444 159934
rect 675392 159870 675444 159876
rect 675404 159664 675432 159870
rect 675484 159384 675536 159390
rect 675484 159326 675536 159332
rect 675496 159052 675524 159326
rect 675484 157752 675536 157758
rect 675484 157694 675536 157700
rect 675496 157216 675524 157694
rect 675392 156936 675444 156942
rect 675392 156878 675444 156884
rect 675404 156643 675432 156878
rect 675758 156496 675814 156505
rect 675758 156431 675814 156440
rect 675772 155992 675800 156431
rect 674748 155712 674800 155718
rect 674748 155654 674800 155660
rect 675484 155712 675536 155718
rect 675484 155654 675536 155660
rect 675496 155380 675524 155654
rect 675392 153400 675444 153406
rect 675392 153342 675444 153348
rect 675404 152864 675432 153342
rect 673828 152584 673880 152590
rect 673828 152526 673880 152532
rect 675392 152584 675444 152590
rect 675392 152526 675444 152532
rect 675404 152320 675432 152526
rect 673644 152040 673696 152046
rect 673644 151982 673696 151988
rect 675392 152040 675444 152046
rect 675392 151982 675444 151988
rect 675404 151675 675432 151982
rect 673552 151428 673604 151434
rect 673552 151370 673604 151376
rect 675392 151428 675444 151434
rect 675392 151370 675444 151376
rect 675404 151028 675432 151370
rect 673460 150408 673512 150414
rect 673460 150350 673512 150356
rect 675392 150408 675444 150414
rect 675392 150350 675444 150356
rect 675404 149835 675432 150350
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675758 146296 675814 146305
rect 675758 146231 675814 146240
rect 675772 146132 675800 146231
rect 676126 133104 676182 133113
rect 676126 133039 676182 133048
rect 676034 132968 676090 132977
rect 676034 132903 676090 132912
rect 676048 132666 676076 132903
rect 676140 132802 676168 133039
rect 676220 132932 676272 132938
rect 676220 132874 676272 132880
rect 676128 132796 676180 132802
rect 676128 132738 676180 132744
rect 676232 132705 676260 132874
rect 676218 132696 676274 132705
rect 676036 132660 676088 132666
rect 676218 132631 676274 132640
rect 676036 132602 676088 132608
rect 676220 132320 676272 132326
rect 676218 132288 676220 132297
rect 676272 132288 676274 132297
rect 676218 132223 676274 132232
rect 676034 131744 676090 131753
rect 676034 131679 676036 131688
rect 676088 131679 676090 131688
rect 676036 131650 676088 131656
rect 673368 131504 673420 131510
rect 676220 131504 676272 131510
rect 673368 131446 673420 131452
rect 676218 131472 676220 131481
rect 676272 131472 676274 131481
rect 676218 131407 676274 131416
rect 676034 130928 676090 130937
rect 676034 130863 676036 130872
rect 676088 130863 676090 130872
rect 676036 130834 676088 130840
rect 676220 130688 676272 130694
rect 676218 130656 676220 130665
rect 676272 130656 676274 130665
rect 676218 130591 676274 130600
rect 676034 130112 676090 130121
rect 676034 130047 676036 130056
rect 676088 130047 676090 130056
rect 676036 130018 676088 130024
rect 676036 129736 676088 129742
rect 676034 129704 676036 129713
rect 676088 129704 676090 129713
rect 676034 129639 676090 129648
rect 676220 129464 676272 129470
rect 676218 129432 676220 129441
rect 676272 129432 676274 129441
rect 676218 129367 676274 129376
rect 676034 128888 676090 128897
rect 676034 128823 676090 128832
rect 675758 128072 675814 128081
rect 675758 128007 675814 128016
rect 674380 127764 674432 127770
rect 674380 127706 674432 127712
rect 673644 127084 673696 127090
rect 673644 127026 673696 127032
rect 673552 124568 673604 124574
rect 673552 124510 673604 124516
rect 673182 122904 673238 122913
rect 673182 122839 673238 122848
rect 672906 112704 672962 112713
rect 672906 112639 672962 112648
rect 673564 107030 673592 124510
rect 673656 108254 673684 127026
rect 673828 123276 673880 123282
rect 673828 123218 673880 123224
rect 673736 121508 673788 121514
rect 673736 121450 673788 121456
rect 673644 108248 673696 108254
rect 673644 108190 673696 108196
rect 673552 107024 673604 107030
rect 673552 106966 673604 106972
rect 673748 106418 673776 121450
rect 673840 107574 673868 123218
rect 674392 114238 674420 127706
rect 674564 127016 674616 127022
rect 674564 126958 674616 126964
rect 674472 124432 674524 124438
rect 674472 124374 674524 124380
rect 674380 114232 674432 114238
rect 674380 114174 674432 114180
rect 673828 107568 673880 107574
rect 673828 107510 673880 107516
rect 673736 106412 673788 106418
rect 673736 106354 673788 106360
rect 672446 105904 672502 105913
rect 672446 105839 672502 105848
rect 674484 105194 674512 124374
rect 674576 112402 674604 126958
rect 675666 124808 675722 124817
rect 675666 124743 675722 124752
rect 675680 124574 675708 124743
rect 675668 124568 675720 124574
rect 675668 124510 675720 124516
rect 674748 124500 674800 124506
rect 674748 124442 674800 124448
rect 674656 124364 674708 124370
rect 674656 124306 674708 124312
rect 674564 112396 674616 112402
rect 674564 112338 674616 112344
rect 674668 111178 674696 124306
rect 674760 111926 674788 124442
rect 675116 124296 675168 124302
rect 675116 124238 675168 124244
rect 674748 111920 674800 111926
rect 674748 111862 674800 111868
rect 674656 111172 674708 111178
rect 674656 111114 674708 111120
rect 675128 110702 675156 124238
rect 675208 124228 675260 124234
rect 675208 124170 675260 124176
rect 675220 115054 675248 124170
rect 675772 115802 675800 128007
rect 676048 127770 676076 128823
rect 676036 127764 676088 127770
rect 676036 127706 676088 127712
rect 676034 127664 676090 127673
rect 676034 127599 676090 127608
rect 675942 127256 675998 127265
rect 675942 127191 675998 127200
rect 675956 127090 675984 127191
rect 675944 127084 675996 127090
rect 675944 127026 675996 127032
rect 676048 127022 676076 127599
rect 676036 127016 676088 127022
rect 676036 126958 676088 126964
rect 676034 126440 676090 126449
rect 676034 126375 676090 126384
rect 675942 126032 675998 126041
rect 675942 125967 675998 125976
rect 675850 125216 675906 125225
rect 675850 125151 675906 125160
rect 675864 124438 675892 125151
rect 675956 124506 675984 125967
rect 675944 124500 675996 124506
rect 675944 124442 675996 124448
rect 675852 124432 675904 124438
rect 675852 124374 675904 124380
rect 675942 124400 675998 124409
rect 675942 124335 675998 124344
rect 675956 124302 675984 124335
rect 675944 124296 675996 124302
rect 675944 124238 675996 124244
rect 676048 124234 676076 126375
rect 676126 125352 676182 125361
rect 676126 125287 676182 125296
rect 676140 124370 676168 125287
rect 676128 124364 676180 124370
rect 676128 124306 676180 124312
rect 676036 124228 676088 124234
rect 676036 124170 676088 124176
rect 676034 123992 676090 124001
rect 676034 123927 676090 123936
rect 675942 123584 675998 123593
rect 675942 123519 675998 123528
rect 675956 121514 675984 123519
rect 676048 123282 676076 123927
rect 676036 123276 676088 123282
rect 676036 123218 676088 123224
rect 676034 123176 676090 123185
rect 676034 123111 676036 123120
rect 676088 123111 676090 123120
rect 676036 123082 676088 123088
rect 676034 122768 676090 122777
rect 676034 122703 676036 122712
rect 676088 122703 676090 122712
rect 676036 122674 676088 122680
rect 676034 121952 676090 121961
rect 676034 121887 676036 121896
rect 676088 121887 676090 121896
rect 676036 121858 676088 121864
rect 675944 121508 675996 121514
rect 675944 121450 675996 121456
rect 675760 115796 675812 115802
rect 675760 115738 675812 115744
rect 675760 115592 675812 115598
rect 675760 115534 675812 115540
rect 675772 115124 675800 115534
rect 675208 115048 675260 115054
rect 675208 114990 675260 114996
rect 675392 115048 675444 115054
rect 675392 114990 675444 114996
rect 675404 114479 675432 114990
rect 675392 114232 675444 114238
rect 675392 114174 675444 114180
rect 675404 113832 675432 114174
rect 675392 112396 675444 112402
rect 675392 112338 675444 112344
rect 675404 111996 675432 112338
rect 675392 111920 675444 111926
rect 675392 111862 675444 111868
rect 675404 111452 675432 111862
rect 675392 111172 675444 111178
rect 675392 111114 675444 111120
rect 675404 110772 675432 111114
rect 675116 110696 675168 110702
rect 675116 110638 675168 110644
rect 675392 110696 675444 110702
rect 675392 110638 675444 110644
rect 675404 110160 675432 110638
rect 675484 108248 675536 108254
rect 675484 108190 675536 108196
rect 675496 107644 675524 108190
rect 675392 107568 675444 107574
rect 675392 107510 675444 107516
rect 675404 107100 675432 107510
rect 675392 107024 675444 107030
rect 675392 106966 675444 106972
rect 675404 106488 675432 106966
rect 675392 106412 675444 106418
rect 675392 106354 675444 106360
rect 675404 105808 675432 106354
rect 674472 105188 674524 105194
rect 674472 105130 674524 105136
rect 675484 105188 675536 105194
rect 675484 105130 675536 105136
rect 675496 104652 675524 105130
rect 675758 103320 675814 103329
rect 675758 103255 675814 103264
rect 675772 102816 675800 103255
rect 671986 102504 672042 102513
rect 671986 102439 672042 102448
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 670882 100872 670938 100881
rect 670882 100807 670938 100816
rect 666558 48512 666614 48521
rect 666558 48447 666614 48456
rect 665178 47424 665234 47433
rect 665178 47359 665234 47368
rect 661130 46240 661186 46249
rect 661130 46175 661186 46184
rect 642824 45620 642876 45626
rect 642824 45562 642876 45568
rect 639328 45552 639380 45558
rect 639328 45494 639380 45500
rect 631876 43308 631928 43314
rect 631876 43250 631928 43256
rect 587990 41576 588046 41585
rect 587990 41511 588046 41520
rect 530214 41304 530270 41313
rect 530214 41239 530270 41248
rect 543002 41304 543058 41313
rect 543002 41239 543058 41248
rect 514024 38616 514076 38622
rect 514024 38558 514076 38564
rect 475568 38548 475620 38554
rect 475568 38490 475620 38496
rect 505652 38548 505704 38554
rect 505652 38490 505704 38496
rect 229376 6520 229428 6526
rect 229376 6462 229428 6468
rect 233148 6520 233200 6526
rect 233148 6462 233200 6468
rect 229388 6225 229416 6462
rect 229374 6216 229430 6225
rect 229374 6151 229430 6160
<< via2 >>
rect 154578 1007428 154580 1007448
rect 154580 1007428 154632 1007448
rect 154632 1007428 154634 1007448
rect 109314 1005372 109370 1005408
rect 109314 1005352 109316 1005372
rect 109316 1005352 109368 1005372
rect 109368 1005352 109370 1005372
rect 87786 995696 87842 995752
rect 85302 995560 85358 995616
rect 82358 995424 82414 995480
rect 81622 995288 81678 995344
rect 80702 995152 80758 995208
rect 84474 994064 84530 994120
rect 80150 993792 80206 993848
rect 78310 993656 78366 993712
rect 106462 1005116 106464 1005136
rect 106464 1005116 106516 1005136
rect 106516 1005116 106518 1005136
rect 106462 1005080 106518 1005116
rect 108026 1004844 108028 1004864
rect 108028 1004844 108080 1004864
rect 108080 1004844 108082 1004864
rect 108026 1004808 108082 1004844
rect 108854 1004828 108910 1004864
rect 108854 1004808 108856 1004828
rect 108856 1004808 108908 1004828
rect 108908 1004808 108910 1004828
rect 92774 995152 92830 995208
rect 41786 968768 41842 968824
rect 41786 965096 41842 965152
rect 41786 963328 41842 963384
rect 35806 949456 35862 949512
rect 41510 943880 41566 943936
rect 41786 943084 41842 943120
rect 41786 943064 41788 943084
rect 41788 943064 41840 943084
rect 41840 943064 41842 943084
rect 41786 942692 41788 942712
rect 41788 942692 41840 942712
rect 41840 942692 41842 942712
rect 41786 942656 41842 942692
rect 41878 942248 41934 942304
rect 41786 941468 41788 941488
rect 41788 941468 41840 941488
rect 41840 941468 41842 941488
rect 41786 941432 41842 941468
rect 41694 940480 41750 940536
rect 41970 941840 42026 941896
rect 41878 941024 41934 941080
rect 41786 936536 41842 936592
rect 35806 934904 35862 934960
rect 35714 934496 35770 934552
rect 35622 934088 35678 934144
rect 41970 940208 42026 940264
rect 41970 938440 42026 938496
rect 42338 938984 42394 939040
rect 42246 938168 42302 938224
rect 41786 933272 41842 933328
rect 41786 932068 41842 932104
rect 41786 932048 41788 932068
rect 41788 932048 41840 932068
rect 41840 932048 41842 932068
rect 41786 817692 41842 817728
rect 41786 817672 41788 817692
rect 41788 817672 41840 817692
rect 41840 817672 41842 817692
rect 41786 817300 41788 817320
rect 41788 817300 41840 817320
rect 41840 817300 41842 817320
rect 41786 817264 41842 817300
rect 42798 938576 42854 938632
rect 42982 939800 43038 939856
rect 42890 933680 42946 933736
rect 42798 921984 42854 922040
rect 41694 815768 41750 815824
rect 41878 816448 41934 816504
rect 41786 814408 41842 814464
rect 42706 816040 42762 816096
rect 42338 814816 42394 814872
rect 41878 814136 41934 814192
rect 41786 813592 41842 813648
rect 41786 811552 41842 811608
rect 41878 811144 41934 811200
rect 41786 808308 41842 808344
rect 41786 808288 41788 808308
rect 41788 808288 41840 808308
rect 41840 808288 41842 808308
rect 41786 807880 41842 807936
rect 41970 807472 42026 807528
rect 41970 806248 42026 806304
rect 41510 774732 41512 774752
rect 41512 774732 41564 774752
rect 41564 774732 41566 774752
rect 41510 774696 41566 774732
rect 41510 774288 41566 774344
rect 41510 773916 41512 773936
rect 41512 773916 41564 773936
rect 41564 773916 41566 773936
rect 41510 773880 41566 773916
rect 42062 773200 42118 773256
rect 41878 767896 41934 767952
rect 41510 764088 41566 764144
rect 41510 762884 41566 762920
rect 41510 762864 41512 762884
rect 41512 762864 41564 762884
rect 41564 762864 41566 762884
rect 41786 757016 41842 757072
rect 41970 766672 42026 766728
rect 42154 771976 42210 772032
rect 42430 769528 42486 769584
rect 41970 757016 42026 757072
rect 42706 767080 42762 767136
rect 42614 755248 42670 755304
rect 41878 754024 41934 754080
rect 39762 731040 39818 731096
rect 39762 730224 39818 730280
rect 43166 937760 43222 937816
rect 43074 937352 43130 937408
rect 43350 936128 43406 936184
rect 43258 935720 43314 935776
rect 43810 927152 43866 927208
rect 43718 815224 43774 815280
rect 43350 814000 43406 814056
rect 42982 813184 43038 813240
rect 42890 812776 42946 812832
rect 43166 810328 43222 810384
rect 43074 809512 43130 809568
rect 43258 809104 43314 809160
rect 43442 812368 43498 812424
rect 43534 811960 43590 812016
rect 43626 808696 43682 808752
rect 43350 772384 43406 772440
rect 43718 771160 43774 771216
rect 42890 770344 42946 770400
rect 43258 769120 43314 769176
rect 43166 768304 43222 768360
rect 43074 766264 43130 766320
rect 42890 764632 42946 764688
rect 42798 730088 42854 730144
rect 43442 768712 43498 768768
rect 43258 765856 43314 765912
rect 43166 765040 43222 765096
rect 43074 752936 43130 752992
rect 42982 729680 43038 729736
rect 43626 767488 43682 767544
rect 43902 810736 43958 810792
rect 43994 809920 44050 809976
rect 44086 770752 44142 770808
rect 43994 769936 44050 769992
rect 43718 765448 43774 765504
rect 43626 757696 43682 757752
rect 41510 729408 41566 729464
rect 41786 728884 41842 728920
rect 41786 728864 41788 728884
rect 41788 728864 41840 728884
rect 41840 728864 41842 728884
rect 39762 728184 39818 728240
rect 44178 730088 44234 730144
rect 43626 728456 43682 728512
rect 42522 727232 42578 727288
rect 43534 726824 43590 726880
rect 42890 726416 42946 726472
rect 41878 724784 41934 724840
rect 41326 723696 41382 723752
rect 41510 720840 41566 720896
rect 41510 719636 41566 719672
rect 41510 719616 41512 719636
rect 41512 719616 41564 719636
rect 41564 719616 41566 719636
rect 42798 723152 42854 723208
rect 43258 726008 43314 726064
rect 42982 724376 43038 724432
rect 43074 723560 43130 723616
rect 41510 688372 41512 688392
rect 41512 688372 41564 688392
rect 41564 688372 41566 688392
rect 41510 688336 41566 688372
rect 41786 687692 41788 687712
rect 41788 687692 41840 687712
rect 41840 687692 41842 687712
rect 41786 687656 41842 687692
rect 41694 687520 41750 687576
rect 43166 721520 43222 721576
rect 43442 725600 43498 725656
rect 43350 725192 43406 725248
rect 43902 722744 43958 722800
rect 43810 721928 43866 721984
rect 43994 722336 44050 722392
rect 44270 727640 44326 727696
rect 44178 686432 44234 686488
rect 43166 685616 43222 685672
rect 42982 684800 43038 684856
rect 42798 684392 42854 684448
rect 41694 681808 41750 681864
rect 43074 682760 43130 682816
rect 42982 682352 43038 682408
rect 41878 681536 41934 681592
rect 41786 678680 41842 678736
rect 41786 677864 41842 677920
rect 41786 676660 41842 676696
rect 41786 676640 41788 676660
rect 41788 676640 41840 676660
rect 41840 676640 41842 676660
rect 41970 678272 42026 678328
rect 41510 645124 41512 645144
rect 41512 645124 41564 645144
rect 41564 645124 41566 645144
rect 41510 645088 41566 645124
rect 41786 644512 41788 644532
rect 41788 644512 41840 644532
rect 41840 644512 41842 644532
rect 41786 644476 41842 644512
rect 41510 644272 41566 644328
rect 43350 685208 43406 685264
rect 43258 680720 43314 680776
rect 43166 643048 43222 643104
rect 44362 686024 44418 686080
rect 44270 683984 44326 684040
rect 43626 683576 43682 683632
rect 43442 680312 43498 680368
rect 43534 679496 43590 679552
rect 43902 683168 43958 683224
rect 43810 681128 43866 681184
rect 43718 679904 43774 679960
rect 43994 679088 44050 679144
rect 44086 643456 44142 643512
rect 43350 641824 43406 641880
rect 42798 641008 42854 641064
rect 43350 640328 43406 640384
rect 42798 639376 42854 639432
rect 41786 638356 41842 638412
rect 30286 634888 30342 634944
rect 41510 634480 41566 634536
rect 41510 633276 41566 633312
rect 41510 633256 41512 633276
rect 41512 633256 41564 633276
rect 41564 633256 41566 633276
rect 42982 637744 43038 637800
rect 42890 637608 42946 637664
rect 43074 636520 43130 636576
rect 43258 636112 43314 636168
rect 43166 635296 43222 635352
rect 43718 639784 43774 639840
rect 43534 638968 43590 639024
rect 43442 636928 43498 636984
rect 43902 638560 43958 638616
rect 43810 635704 43866 635760
rect 41510 601876 41512 601896
rect 41512 601876 41564 601896
rect 41564 601876 41566 601896
rect 41510 601840 41566 601876
rect 42430 600480 42486 600536
rect 44822 642232 44878 642288
rect 44362 641960 44418 642016
rect 44178 600072 44234 600128
rect 43442 599256 43498 599312
rect 41878 595176 41934 595232
rect 41142 594088 41198 594144
rect 41510 591232 41566 591288
rect 41510 590028 41566 590064
rect 41510 590008 41512 590028
rect 41512 590008 41564 590028
rect 41564 590008 41566 590028
rect 43258 597216 43314 597272
rect 42890 596808 42946 596864
rect 42798 593544 42854 593600
rect 43074 596400 43130 596456
rect 42982 594768 43038 594824
rect 41510 558764 41512 558784
rect 41512 558764 41564 558784
rect 41564 558764 41566 558784
rect 41510 558728 41566 558764
rect 41510 558320 41566 558376
rect 41418 557912 41474 557968
rect 43166 593952 43222 594008
rect 43350 595584 43406 595640
rect 42798 556824 42854 556880
rect 44638 641144 44694 641200
rect 44362 598440 44418 598496
rect 43994 598032 44050 598088
rect 43810 595992 43866 596048
rect 43718 593136 43774 593192
rect 43626 592320 43682 592376
rect 43534 591912 43590 591968
rect 43902 592728 43958 592784
rect 44822 599664 44878 599720
rect 44638 597624 44694 597680
rect 43442 556416 43498 556472
rect 43258 554376 43314 554432
rect 43810 553968 43866 554024
rect 42706 553560 42762 553616
rect 41786 551928 41842 551984
rect 41510 548936 41566 548992
rect 41510 548528 41566 548584
rect 41602 548120 41658 548176
rect 41602 546916 41658 546952
rect 41602 546896 41604 546916
rect 41604 546896 41656 546916
rect 41656 546896 41658 546916
rect 43166 553152 43222 553208
rect 43074 551112 43130 551168
rect 42982 550296 43038 550352
rect 42890 540912 42946 540968
rect 43350 552744 43406 552800
rect 43258 549888 43314 549944
rect 43626 552336 43682 552392
rect 43442 551520 43498 551576
rect 43994 550704 44050 550760
rect 43902 549480 43958 549536
rect 44086 540776 44142 540832
rect 42890 450744 42946 450800
rect 41786 430888 41842 430944
rect 43074 430616 43130 430672
rect 43626 429664 43682 429720
rect 43074 429256 43130 429312
rect 41786 426808 41842 426864
rect 42890 426400 42946 426456
rect 42798 425992 42854 426048
rect 42338 424360 42394 424416
rect 41878 421504 41934 421560
rect 41786 420688 41842 420744
rect 41786 419484 41842 419520
rect 41786 419464 41788 419484
rect 41788 419464 41840 419484
rect 41840 419464 41842 419484
rect 42522 421096 42578 421152
rect 42798 411212 42854 411268
rect 41142 389000 41198 389056
rect 41510 387948 41512 387968
rect 41512 387948 41564 387968
rect 41564 387948 41566 387968
rect 41510 387912 41566 387948
rect 41510 387504 41566 387560
rect 41510 387132 41512 387152
rect 41512 387132 41564 387152
rect 41564 387132 41566 387152
rect 41510 387096 41566 387132
rect 41142 386688 41198 386744
rect 43258 425584 43314 425640
rect 42982 422728 43038 422784
rect 43166 422320 43222 422376
rect 43350 425176 43406 425232
rect 43442 424768 43498 424824
rect 43534 423136 43590 423192
rect 43810 428440 43866 428496
rect 43718 423544 43774 423600
rect 43626 411440 43682 411496
rect 43902 423952 43958 424008
rect 43994 421912 44050 421968
rect 42798 386008 42854 386064
rect 43810 385600 43866 385656
rect 43534 385192 43590 385248
rect 41142 384648 41198 384704
rect 43350 383152 43406 383208
rect 42798 382744 42854 382800
rect 42338 381112 42394 381168
rect 41510 377712 41566 377768
rect 41602 377304 41658 377360
rect 41602 376100 41658 376136
rect 41602 376080 41604 376100
rect 41604 376080 41656 376100
rect 41656 376080 41658 376100
rect 42982 381928 43038 381984
rect 42890 379480 42946 379536
rect 43166 379072 43222 379128
rect 43074 378256 43130 378312
rect 43258 378664 43314 378720
rect 43442 380704 43498 380760
rect 41786 355680 41842 355736
rect 33046 351872 33102 351928
rect 43902 381520 43958 381576
rect 43626 380296 43682 380352
rect 43718 379888 43774 379944
rect 33046 343032 33102 343088
rect 41786 344528 41842 344584
rect 41602 344292 41604 344312
rect 41604 344292 41656 344312
rect 41656 344292 41658 344312
rect 41602 344256 41658 344292
rect 41602 343884 41604 343904
rect 41604 343884 41656 343904
rect 41656 343884 41658 343904
rect 41602 343848 41658 343884
rect 41786 343340 41788 343360
rect 41788 343340 41840 343360
rect 41840 343340 41842 343360
rect 41786 343304 41842 343340
rect 41510 342624 41566 342680
rect 43258 342080 43314 342136
rect 32678 339768 32734 339824
rect 32770 338136 32826 338192
rect 33046 337728 33102 337784
rect 32862 336096 32918 336152
rect 32954 335688 33010 335744
rect 43074 335552 43130 335608
rect 42982 335144 43038 335200
rect 41510 334056 41566 334112
rect 41510 332852 41566 332888
rect 41510 332832 41512 332852
rect 41512 332832 41564 332852
rect 41564 332832 41566 332852
rect 32770 329704 32826 329760
rect 41786 319912 41842 319968
rect 43166 334736 43222 334792
rect 42154 316920 42210 316976
rect 42154 316240 42210 316296
rect 41970 315560 42026 315616
rect 41878 313792 41934 313848
rect 41786 312976 41842 313032
rect 42154 312296 42210 312352
rect 41510 301588 41512 301608
rect 41512 301588 41564 301608
rect 41564 301588 41566 301608
rect 41510 301552 41566 301588
rect 41786 300908 41788 300928
rect 41788 300908 41840 300928
rect 41840 300908 41842 300928
rect 41786 300872 41842 300908
rect 44270 341672 44326 341728
rect 44362 340856 44418 340912
rect 44270 339904 44326 339960
rect 44178 299648 44234 299704
rect 43074 299240 43130 299296
rect 43442 298832 43498 298888
rect 32586 296792 32642 296848
rect 32678 296384 32734 296440
rect 32954 295976 33010 296032
rect 32862 295160 32918 295216
rect 32770 292304 32826 292360
rect 32586 285640 32642 285696
rect 41878 294752 41934 294808
rect 33046 294344 33102 294400
rect 41786 293936 41842 293992
rect 41786 291896 41842 291952
rect 41786 291488 41842 291544
rect 42430 293528 42486 293584
rect 33046 285912 33102 285968
rect 32954 285776 33010 285832
rect 43074 293120 43130 293176
rect 43258 292712 43314 292768
rect 41970 272312 42026 272368
rect 42154 270408 42210 270464
rect 42154 270000 42210 270056
rect 42154 269320 42210 269376
rect 41510 258340 41512 258360
rect 41512 258340 41564 258360
rect 41564 258340 41566 258360
rect 41510 258304 41566 258340
rect 41510 257896 41566 257952
rect 41510 257524 41512 257544
rect 41512 257524 41564 257544
rect 41564 257524 41566 257544
rect 41510 257488 41566 257524
rect 41786 256844 41788 256864
rect 41788 256844 41840 256864
rect 41840 256844 41842 256864
rect 41786 256808 41842 256844
rect 44362 339496 44418 339552
rect 44270 298016 44326 298072
rect 44362 297200 44418 297256
rect 45374 289856 45430 289912
rect 43442 255992 43498 256048
rect 43442 255584 43498 255640
rect 42706 253544 42762 253600
rect 31666 253000 31722 253056
rect 33046 251776 33102 251832
rect 32770 250552 32826 250608
rect 32862 250144 32918 250200
rect 32954 249736 33010 249792
rect 38290 248104 38346 248160
rect 41510 247716 41566 247752
rect 41510 247696 41512 247716
rect 41512 247696 41564 247716
rect 41564 247696 41566 247716
rect 41510 247308 41566 247344
rect 41510 247288 41512 247308
rect 41512 247288 41564 247308
rect 41564 247288 41566 247308
rect 41510 246492 41566 246528
rect 41510 246472 41512 246492
rect 41512 246472 41564 246492
rect 41564 246472 41566 246492
rect 42798 252320 42854 252376
rect 43258 249464 43314 249520
rect 43166 248648 43222 248704
rect 43350 249056 43406 249112
rect 41970 225936 42026 225992
rect 29182 204448 29238 204504
rect 41510 215056 41566 215112
rect 41602 214648 41658 214704
rect 41418 214240 41474 214296
rect 43810 251504 43866 251560
rect 43902 251096 43958 251152
rect 41418 213868 41420 213888
rect 41420 213868 41472 213888
rect 41472 213868 41474 213888
rect 41418 213832 41474 213868
rect 41510 213016 41566 213072
rect 45926 255176 45982 255232
rect 45742 254360 45798 254416
rect 46202 339904 46258 339960
rect 46110 298424 46166 298480
rect 46110 290672 46166 290728
rect 46478 683984 46534 684040
rect 46386 339496 46442 339552
rect 46386 291080 46442 291136
rect 46570 598440 46626 598496
rect 46754 597624 46810 597680
rect 58438 975976 58494 976032
rect 57978 962920 58034 962976
rect 58438 949864 58494 949920
rect 58438 936944 58494 937000
rect 58438 923752 58494 923808
rect 48318 300056 48374 300112
rect 48226 297608 48282 297664
rect 59174 910696 59230 910752
rect 48594 730904 48650 730960
rect 51262 731312 51318 731368
rect 51078 730496 51134 730552
rect 58438 897776 58494 897832
rect 58438 884720 58494 884776
rect 58438 871664 58494 871720
rect 58438 858608 58494 858664
rect 58438 845552 58494 845608
rect 57978 832496 58034 832552
rect 53838 816856 53894 816912
rect 59174 819440 59230 819496
rect 58438 806520 58494 806576
rect 58070 793464 58126 793520
rect 58438 780408 58494 780464
rect 58438 767372 58494 767408
rect 58438 767352 58440 767372
rect 58440 767352 58492 767372
rect 58492 767352 58494 767372
rect 58346 754296 58402 754352
rect 58438 741240 58494 741296
rect 58438 728184 58494 728240
rect 58438 715264 58494 715320
rect 58622 702208 58678 702264
rect 58438 689152 58494 689208
rect 58438 676096 58494 676152
rect 58438 663040 58494 663096
rect 59174 649984 59230 650040
rect 51078 601296 51134 601352
rect 58438 637064 58494 637120
rect 58438 624008 58494 624064
rect 58438 610952 58494 611008
rect 53838 600888 53894 600944
rect 59174 597896 59230 597952
rect 58438 584840 58494 584896
rect 58438 571784 58494 571840
rect 58346 558728 58402 558784
rect 58346 545808 58402 545864
rect 51262 430480 51318 430536
rect 59266 532752 59322 532808
rect 58438 519696 58494 519752
rect 58438 506640 58494 506696
rect 57978 493584 58034 493640
rect 58438 480528 58494 480584
rect 58714 467472 58770 467528
rect 53838 430072 53894 430128
rect 59174 454552 59230 454608
rect 58438 441496 58494 441552
rect 58254 428440 58310 428496
rect 58438 415384 58494 415440
rect 58438 402328 58494 402384
rect 57978 389272 58034 389328
rect 62118 386280 62174 386336
rect 62302 939392 62358 939448
rect 62210 383424 62266 383480
rect 62026 383016 62082 383072
rect 58438 376216 58494 376272
rect 58438 363296 58494 363352
rect 58438 350240 58494 350296
rect 58438 337184 58494 337240
rect 58162 324128 58218 324184
rect 53838 300464 53894 300520
rect 59266 311072 59322 311128
rect 46938 212472 46994 212528
rect 45650 212064 45706 212120
rect 45466 211248 45522 211304
rect 32954 209752 33010 209808
rect 31666 203632 31722 203688
rect 33046 208120 33102 208176
rect 42890 206760 42946 206816
rect 42798 205128 42854 205184
rect 43074 206352 43130 206408
rect 42982 205536 43038 205592
rect 48226 204720 48282 204776
rect 42154 190168 42210 190224
rect 41878 187584 41934 187640
rect 42154 187040 42210 187096
rect 41970 186360 42026 186416
rect 42154 185816 42210 185872
rect 42154 184184 42210 184240
rect 41786 183640 41842 183696
rect 41786 182688 41842 182744
rect 57610 227704 57666 227760
rect 56046 227568 56102 227624
rect 55126 224984 55182 225040
rect 54390 222128 54446 222184
rect 56874 224848 56930 224904
rect 59358 298152 59414 298208
rect 59450 285096 59506 285152
rect 62486 938440 62542 938496
rect 62302 278296 62358 278352
rect 62578 596128 62634 596184
rect 62578 430616 62634 430672
rect 98274 1004692 98330 1004728
rect 98274 1004672 98276 1004692
rect 98276 1004672 98328 1004692
rect 98328 1004672 98330 1004692
rect 99102 1004692 99158 1004728
rect 99102 1004672 99104 1004692
rect 99104 1004672 99156 1004692
rect 99156 1004672 99158 1004692
rect 105634 1004708 105636 1004728
rect 105636 1004708 105688 1004728
rect 105688 1004708 105690 1004728
rect 105634 1004672 105690 1004708
rect 102782 999796 102838 999832
rect 102782 999776 102784 999796
rect 102784 999776 102836 999796
rect 102836 999776 102838 999796
rect 104346 999812 104348 999832
rect 104348 999812 104400 999832
rect 104400 999812 104402 999832
rect 104346 999776 104402 999812
rect 100666 999676 100668 999696
rect 100668 999676 100720 999696
rect 100720 999676 100722 999696
rect 100666 999640 100722 999676
rect 102322 999660 102378 999696
rect 102322 999640 102324 999660
rect 102324 999640 102376 999660
rect 102376 999640 102378 999660
rect 101494 999524 101550 999560
rect 101494 999504 101496 999524
rect 101496 999504 101548 999524
rect 101548 999504 101550 999524
rect 101954 999540 101956 999560
rect 101956 999540 102008 999560
rect 102008 999540 102010 999560
rect 101954 999504 102010 999540
rect 95698 996376 95754 996432
rect 95514 995560 95570 995616
rect 97354 995560 97410 995616
rect 95330 995424 95386 995480
rect 95146 995288 95202 995344
rect 99470 999388 99526 999424
rect 99470 999368 99472 999388
rect 99472 999368 99524 999388
rect 99524 999368 99526 999388
rect 103150 999404 103152 999424
rect 103152 999404 103204 999424
rect 103204 999404 103206 999424
rect 103150 999368 103206 999404
rect 100298 999252 100354 999288
rect 100298 999232 100300 999252
rect 100300 999232 100352 999252
rect 100352 999232 100354 999252
rect 101126 999268 101128 999288
rect 101128 999268 101180 999288
rect 101180 999268 101182 999288
rect 101126 999232 101182 999268
rect 99930 999132 99932 999152
rect 99932 999132 99984 999152
rect 99984 999132 99986 999152
rect 99930 999096 99986 999132
rect 107658 997212 107714 997248
rect 107658 997192 107660 997212
rect 107660 997192 107712 997212
rect 107712 997192 107714 997212
rect 115938 997212 115994 997248
rect 115938 997192 115940 997212
rect 115940 997192 115992 997212
rect 115992 997192 115994 997212
rect 108486 996124 108542 996160
rect 108486 996104 108488 996124
rect 108488 996104 108540 996124
rect 108540 996104 108542 996124
rect 113270 995832 113326 995888
rect 110418 995696 110474 995752
rect 104162 995560 104218 995616
rect 104346 995560 104402 995616
rect 97906 994064 97962 994120
rect 97354 993792 97410 993848
rect 104346 993656 104402 993712
rect 110510 995560 110566 995616
rect 110602 995424 110658 995480
rect 143814 1005080 143870 1005136
rect 143722 1004944 143778 1005000
rect 142802 995696 142858 995752
rect 143998 997192 144054 997248
rect 137374 995560 137430 995616
rect 133694 995424 133750 995480
rect 143998 995424 144054 995480
rect 154578 1007392 154634 1007428
rect 501326 1007256 501382 1007312
rect 424690 1006052 424746 1006088
rect 424690 1006032 424692 1006052
rect 424692 1006032 424744 1006052
rect 424744 1006032 424746 1006052
rect 423862 1005916 423918 1005952
rect 423862 1005896 423864 1005916
rect 423864 1005896 423916 1005916
rect 423916 1005896 423918 1005916
rect 424322 1005796 424324 1005816
rect 424324 1005796 424376 1005816
rect 424376 1005796 424378 1005816
rect 424322 1005760 424378 1005796
rect 356058 1005660 356060 1005680
rect 356060 1005660 356112 1005680
rect 356112 1005660 356114 1005680
rect 356058 1005624 356114 1005660
rect 356518 1005644 356574 1005680
rect 356518 1005624 356520 1005644
rect 356520 1005624 356572 1005644
rect 356572 1005624 356574 1005644
rect 160282 1005508 160338 1005544
rect 207202 1005524 207204 1005544
rect 207204 1005524 207256 1005544
rect 207256 1005524 207258 1005544
rect 160282 1005488 160284 1005508
rect 160284 1005488 160336 1005508
rect 160336 1005488 160338 1005508
rect 153750 1005372 153806 1005408
rect 153750 1005352 153752 1005372
rect 153752 1005352 153804 1005372
rect 153804 1005352 153806 1005372
rect 154946 1005388 154948 1005408
rect 154948 1005388 155000 1005408
rect 155000 1005388 155002 1005408
rect 154946 1005352 155002 1005388
rect 151266 1005236 151322 1005272
rect 151266 1005216 151268 1005236
rect 151268 1005216 151320 1005236
rect 151320 1005216 151322 1005236
rect 153290 1005252 153292 1005272
rect 153292 1005252 153344 1005272
rect 153344 1005252 153346 1005272
rect 153290 1005216 153346 1005252
rect 148874 1005080 148930 1005136
rect 149702 1005100 149758 1005136
rect 149702 1005080 149704 1005100
rect 149704 1005080 149756 1005100
rect 149756 1005080 149758 1005100
rect 150438 1005100 150494 1005136
rect 150438 1005080 150440 1005100
rect 150440 1005080 150492 1005100
rect 150492 1005080 150494 1005100
rect 148874 1004980 148876 1005000
rect 148876 1004980 148928 1005000
rect 148928 1004980 148930 1005000
rect 148874 1004944 148930 1004980
rect 150898 1004980 150900 1005000
rect 150900 1004980 150952 1005000
rect 150952 1004980 150954 1005000
rect 150898 1004944 150954 1004980
rect 154118 1004964 154174 1005000
rect 154118 1004944 154120 1004964
rect 154120 1004944 154172 1004964
rect 154172 1004944 154174 1004964
rect 159454 1004964 159510 1005000
rect 159454 1004944 159456 1004964
rect 159456 1004944 159508 1004964
rect 159508 1004944 159510 1004964
rect 147586 1004808 147642 1004864
rect 147770 1004672 147826 1004728
rect 148874 1004844 148876 1004864
rect 148876 1004844 148928 1004864
rect 148928 1004844 148930 1004864
rect 148874 1004808 148930 1004844
rect 152094 1004844 152096 1004864
rect 152096 1004844 152148 1004864
rect 152148 1004844 152150 1004864
rect 152094 1004808 152150 1004844
rect 152922 1004828 152978 1004864
rect 152922 1004808 152924 1004828
rect 152924 1004808 152976 1004828
rect 152976 1004808 152978 1004828
rect 156970 1004828 157026 1004864
rect 156970 1004808 156972 1004828
rect 156972 1004808 157024 1004828
rect 157024 1004808 157026 1004828
rect 148874 1004708 148876 1004728
rect 148876 1004708 148928 1004728
rect 148928 1004708 148930 1004728
rect 148874 1004672 148930 1004708
rect 151726 1004708 151728 1004728
rect 151728 1004708 151780 1004728
rect 151780 1004708 151782 1004728
rect 151726 1004672 151782 1004708
rect 152554 1004692 152610 1004728
rect 157798 1004708 157800 1004728
rect 157800 1004708 157852 1004728
rect 157852 1004708 157854 1004728
rect 152554 1004672 152556 1004692
rect 152556 1004672 152608 1004692
rect 152608 1004672 152610 1004692
rect 157798 1004672 157854 1004708
rect 160650 1004692 160706 1004728
rect 160650 1004672 160652 1004692
rect 160652 1004672 160704 1004692
rect 160704 1004672 160706 1004692
rect 148138 996376 148194 996432
rect 147586 995560 147642 995616
rect 155774 999540 155776 999560
rect 155776 999540 155828 999560
rect 155828 999540 155830 999560
rect 155774 999504 155830 999540
rect 159086 999524 159142 999560
rect 159086 999504 159088 999524
rect 159088 999504 159140 999524
rect 159140 999504 159142 999524
rect 155774 999132 155776 999152
rect 155776 999132 155828 999152
rect 155828 999132 155830 999152
rect 155774 999096 155830 999132
rect 158258 999116 158314 999152
rect 158258 999096 158260 999116
rect 158260 999096 158312 999116
rect 158312 999096 158314 999116
rect 156142 997756 156198 997792
rect 156142 997736 156144 997756
rect 156144 997736 156196 997756
rect 156196 997736 156198 997756
rect 156970 996099 157026 996155
rect 157798 996135 157800 996155
rect 157800 996135 157852 996155
rect 157852 996135 157854 996155
rect 157798 996099 157854 996135
rect 159454 996119 159510 996155
rect 159454 996099 159456 996119
rect 159456 996099 159508 996119
rect 159508 996099 159510 996119
rect 168858 997056 168914 997112
rect 162950 995696 163006 995752
rect 162858 995560 162914 995616
rect 168378 993672 168434 993728
rect 195150 997192 195206 997248
rect 195334 997056 195390 997112
rect 187606 995696 187662 995752
rect 192482 995560 192538 995616
rect 207202 1005488 207258 1005524
rect 209594 1005508 209650 1005544
rect 209594 1005488 209596 1005508
rect 209596 1005488 209648 1005508
rect 209648 1005488 209650 1005508
rect 361026 1005508 361082 1005544
rect 361026 1005488 361028 1005508
rect 361028 1005488 361080 1005508
rect 361080 1005488 361082 1005508
rect 263852 1005408 263908 1005464
rect 259826 1005252 259828 1005272
rect 259828 1005252 259880 1005272
rect 259880 1005252 259882 1005272
rect 259826 1005216 259882 1005252
rect 260194 1005236 260250 1005272
rect 260194 1005216 260196 1005236
rect 260196 1005216 260248 1005236
rect 260248 1005216 260250 1005236
rect 208398 1005100 208454 1005136
rect 261850 1005116 261852 1005136
rect 261852 1005116 261904 1005136
rect 261904 1005116 261906 1005136
rect 208398 1005080 208400 1005100
rect 208400 1005080 208452 1005100
rect 208452 1005080 208454 1005100
rect 209226 1004964 209282 1005000
rect 209226 1004944 209228 1004964
rect 209228 1004944 209280 1004964
rect 209280 1004944 209282 1004964
rect 211618 1004980 211620 1005000
rect 211620 1004980 211672 1005000
rect 211672 1004980 211674 1005000
rect 211618 1004944 211674 1004980
rect 201038 1004708 201040 1004728
rect 201040 1004708 201092 1004728
rect 201092 1004708 201094 1004728
rect 201038 1004672 201094 1004708
rect 201866 1004708 201868 1004728
rect 201868 1004708 201920 1004728
rect 201920 1004708 201922 1004728
rect 201866 1004672 201922 1004708
rect 203890 999660 203946 999696
rect 203890 999640 203892 999660
rect 203892 999640 203944 999660
rect 203944 999640 203946 999660
rect 203522 999540 203524 999560
rect 203524 999540 203576 999560
rect 203576 999540 203578 999560
rect 203522 999504 203578 999540
rect 202234 999388 202290 999424
rect 202234 999368 202236 999388
rect 202236 999368 202288 999388
rect 202288 999368 202290 999388
rect 202694 999252 202750 999288
rect 202694 999232 202696 999252
rect 202696 999232 202748 999252
rect 202748 999232 202750 999252
rect 203062 999132 203064 999152
rect 203064 999132 203116 999152
rect 203116 999132 203118 999152
rect 203062 999096 203118 999132
rect 191838 993656 191894 993712
rect 206374 1004828 206430 1004864
rect 206374 1004808 206376 1004828
rect 206376 1004808 206428 1004828
rect 206428 1004808 206430 1004828
rect 210882 1004844 210884 1004864
rect 210884 1004844 210936 1004864
rect 210936 1004844 210938 1004864
rect 210882 1004808 210938 1004844
rect 205914 1004692 205970 1004728
rect 205914 1004672 205916 1004692
rect 205916 1004672 205968 1004692
rect 205968 1004672 205970 1004692
rect 212458 1004672 212514 1004728
rect 205546 999676 205548 999696
rect 205548 999676 205600 999696
rect 205600 999676 205602 999696
rect 205546 999640 205602 999676
rect 204350 999524 204406 999560
rect 204350 999504 204352 999524
rect 204352 999504 204404 999524
rect 204404 999504 204406 999524
rect 204718 999404 204720 999424
rect 204720 999404 204772 999424
rect 204772 999404 204774 999424
rect 204718 999368 204774 999404
rect 208858 999404 208860 999424
rect 208860 999404 208912 999424
rect 208912 999404 208914 999424
rect 208858 999368 208914 999404
rect 210422 999388 210478 999424
rect 210422 999368 210424 999388
rect 210424 999368 210476 999388
rect 210476 999368 210478 999388
rect 205178 999268 205180 999288
rect 205180 999268 205232 999288
rect 205232 999268 205234 999288
rect 205178 999232 205234 999268
rect 209594 999268 209596 999288
rect 209596 999268 209648 999288
rect 209648 999268 209650 999288
rect 209594 999232 209650 999268
rect 211710 999252 211766 999288
rect 211710 999232 211712 999252
rect 211712 999232 211764 999252
rect 211764 999232 211766 999252
rect 207570 999096 207626 999152
rect 211250 999132 211252 999152
rect 211252 999132 211304 999152
rect 211304 999132 211306 999152
rect 211250 999096 211306 999132
rect 218970 997192 219026 997248
rect 261850 1005080 261906 1005116
rect 263046 1005100 263102 1005136
rect 263046 1005080 263048 1005100
rect 263048 1005080 263100 1005100
rect 263100 1005080 263102 1005100
rect 260654 1004980 260656 1005000
rect 260656 1004980 260708 1005000
rect 260708 1004980 260710 1005000
rect 260654 1004944 260710 1004980
rect 262678 1004964 262734 1005000
rect 262678 1004944 262680 1004964
rect 262680 1004944 262732 1004964
rect 262732 1004944 262734 1004964
rect 261022 1004844 261024 1004864
rect 261024 1004844 261076 1004864
rect 261076 1004844 261078 1004864
rect 261022 1004808 261078 1004844
rect 262218 1004828 262274 1004864
rect 262218 1004808 262220 1004828
rect 262220 1004808 262272 1004828
rect 262272 1004808 262274 1004828
rect 252466 1004692 252522 1004728
rect 252466 1004672 252468 1004692
rect 252468 1004672 252520 1004692
rect 252520 1004672 252522 1004692
rect 253294 1004692 253350 1004728
rect 253294 1004672 253296 1004692
rect 253296 1004672 253348 1004692
rect 253348 1004672 253350 1004692
rect 261482 1004708 261484 1004728
rect 261484 1004708 261536 1004728
rect 261536 1004708 261538 1004728
rect 261482 1004672 261538 1004708
rect 263506 1004672 263562 1004728
rect 258630 999932 258686 999968
rect 258630 999912 258632 999932
rect 258632 999912 258684 999932
rect 258684 999912 258686 999932
rect 235262 995696 235318 995752
rect 235906 995696 235962 995752
rect 242070 995696 242126 995752
rect 256974 999796 257030 999832
rect 256974 999776 256976 999796
rect 256976 999776 257028 999796
rect 257028 999776 257030 999796
rect 257342 999812 257344 999832
rect 257344 999812 257396 999832
rect 257396 999812 257398 999832
rect 257342 999776 257398 999812
rect 240046 995560 240102 995616
rect 232226 994064 232282 994120
rect 236550 995424 236606 995480
rect 234388 995288 234444 995344
rect 232870 993928 232926 993984
rect 254858 999660 254914 999696
rect 254858 999640 254860 999660
rect 254860 999640 254912 999660
rect 254912 999640 254914 999660
rect 257802 999676 257804 999696
rect 257804 999676 257856 999696
rect 257856 999676 257858 999696
rect 257802 999640 257858 999676
rect 247958 997192 248014 997248
rect 249706 995560 249762 995616
rect 255686 999524 255742 999560
rect 255686 999504 255688 999524
rect 255688 999504 255740 999524
rect 255740 999504 255742 999524
rect 256146 999540 256148 999560
rect 256148 999540 256200 999560
rect 256200 999540 256202 999560
rect 256146 999504 256202 999540
rect 253662 999388 253718 999424
rect 253662 999368 253664 999388
rect 253664 999368 253716 999388
rect 253716 999368 253718 999388
rect 255318 999404 255320 999424
rect 255320 999404 255372 999424
rect 255372 999404 255374 999424
rect 255318 999368 255374 999404
rect 254490 999268 254492 999288
rect 254492 999268 254544 999288
rect 254544 999268 254546 999288
rect 254490 999232 254546 999268
rect 256514 999252 256570 999288
rect 256514 999232 256516 999252
rect 256516 999232 256568 999252
rect 256568 999232 256570 999252
rect 250442 995968 250498 996024
rect 250258 995832 250314 995888
rect 250074 995696 250130 995752
rect 249890 995424 249946 995480
rect 246854 995288 246910 995344
rect 254122 999132 254124 999152
rect 254124 999132 254176 999152
rect 254176 999132 254178 999152
rect 254122 999096 254178 999132
rect 258538 999132 258540 999152
rect 258540 999132 258592 999152
rect 258592 999132 258594 999152
rect 258538 999096 258594 999132
rect 252466 994064 252522 994120
rect 243266 993792 243322 993848
rect 248326 993656 248382 993712
rect 265534 1005100 265590 1005136
rect 265534 1005080 265536 1005100
rect 265536 1005080 265588 1005100
rect 265588 1005080 265590 1005100
rect 265534 1004964 265590 1005000
rect 265534 1004944 265536 1004964
rect 265536 1004944 265588 1004964
rect 265588 1004944 265590 1004964
rect 266630 1004944 266686 1005000
rect 265474 1004672 265530 1004728
rect 266538 1004672 266594 1004728
rect 360198 1005372 360254 1005408
rect 360198 1005352 360200 1005372
rect 360200 1005352 360252 1005372
rect 360252 1005352 360254 1005372
rect 267010 1005080 267066 1005136
rect 270466 997192 270522 997248
rect 359738 1005236 359794 1005272
rect 359738 1005216 359740 1005236
rect 359740 1005216 359792 1005236
rect 359792 1005216 359794 1005236
rect 358174 1005100 358230 1005136
rect 358174 1005080 358176 1005100
rect 358176 1005080 358228 1005100
rect 358228 1005080 358230 1005100
rect 356886 1004980 356888 1005000
rect 356888 1004980 356940 1005000
rect 356940 1004980 356942 1005000
rect 356886 1004944 356942 1004980
rect 358542 1004964 358598 1005000
rect 358542 1004944 358544 1004964
rect 358544 1004944 358596 1004964
rect 358596 1004944 358598 1004964
rect 357346 1004844 357348 1004864
rect 357348 1004844 357400 1004864
rect 357400 1004844 357402 1004864
rect 357346 1004808 357402 1004844
rect 357714 1004828 357770 1004864
rect 357714 1004808 357716 1004828
rect 357716 1004808 357768 1004828
rect 357768 1004808 357770 1004828
rect 315118 1004692 315174 1004728
rect 315118 1004672 315120 1004692
rect 315120 1004672 315172 1004692
rect 315172 1004672 315174 1004692
rect 350446 1004672 350502 1004728
rect 353666 1004672 353722 1004728
rect 354034 1004672 354090 1004728
rect 354494 1004672 354550 1004728
rect 355230 1004672 355286 1004728
rect 360566 1004708 360568 1004728
rect 360568 1004708 360620 1004728
rect 360620 1004708 360622 1004728
rect 360566 1004672 360622 1004708
rect 361394 1004692 361450 1004728
rect 361394 1004672 361396 1004692
rect 361396 1004672 361448 1004692
rect 361448 1004672 361450 1004692
rect 310150 999796 310206 999832
rect 310150 999776 310152 999796
rect 310152 999776 310204 999796
rect 310204 999776 310206 999796
rect 312174 999812 312176 999832
rect 312176 999812 312228 999832
rect 312228 999812 312230 999832
rect 312174 999776 312230 999812
rect 311438 999676 311440 999696
rect 311440 999676 311492 999696
rect 311492 999676 311494 999696
rect 311438 999640 311494 999676
rect 313830 999660 313886 999696
rect 313830 999640 313832 999660
rect 313832 999640 313884 999660
rect 313884 999640 313886 999660
rect 312634 999540 312636 999560
rect 312636 999540 312688 999560
rect 312688 999540 312690 999560
rect 312634 999504 312690 999540
rect 314658 999504 314714 999560
rect 312634 999116 312690 999152
rect 312634 999096 312636 999116
rect 312636 999096 312688 999116
rect 312688 999096 312690 999116
rect 298742 997192 298798 997248
rect 288070 995696 288126 995752
rect 292486 995696 292542 995752
rect 300766 995832 300822 995888
rect 291106 995560 291162 995616
rect 300214 995560 300270 995616
rect 290554 995424 290610 995480
rect 297270 995424 297326 995480
rect 294510 993656 294566 993712
rect 305734 996260 305790 996296
rect 305734 996240 305736 996260
rect 305736 996240 305788 996260
rect 305788 996240 305790 996260
rect 308126 996276 308128 996296
rect 308128 996276 308180 996296
rect 308180 996276 308182 996296
rect 308126 996240 308182 996276
rect 305274 996104 305330 996160
rect 306470 996104 306526 996160
rect 306930 996104 306986 996160
rect 307298 996104 307354 996160
rect 307758 996104 307814 996160
rect 309322 996104 309378 996160
rect 310150 996104 310206 996160
rect 310610 996104 310666 996160
rect 311806 996104 311862 996160
rect 314290 996140 314292 996160
rect 314292 996140 314344 996160
rect 314344 996140 314346 996160
rect 314290 996104 314346 996140
rect 305274 995560 305330 995616
rect 316774 993792 316830 993848
rect 321466 993524 321522 993580
rect 358910 1000492 358912 1000512
rect 358912 1000492 358964 1000512
rect 358964 1000492 358966 1000512
rect 358910 1000456 358966 1000492
rect 361854 999676 361856 999696
rect 361856 999676 361908 999696
rect 361908 999676 361910 999696
rect 361854 999640 361910 999676
rect 362590 999660 362646 999696
rect 362590 999640 362592 999660
rect 362592 999640 362644 999660
rect 362644 999640 362646 999660
rect 363418 999540 363420 999560
rect 363420 999540 363472 999560
rect 363472 999540 363474 999560
rect 363418 999504 363474 999540
rect 362222 999404 362224 999424
rect 362224 999404 362276 999424
rect 362276 999404 362278 999424
rect 362222 999368 362278 999404
rect 364246 999252 364302 999288
rect 364246 999232 364248 999252
rect 364248 999232 364300 999252
rect 364300 999232 364302 999252
rect 358910 999132 358912 999152
rect 358912 999132 358964 999152
rect 358964 999132 358966 999152
rect 358910 999096 358966 999132
rect 363050 999132 363052 999152
rect 363052 999132 363104 999152
rect 363104 999132 363106 999152
rect 363050 999096 363106 999132
rect 371330 1004672 371386 1004728
rect 365074 999524 365130 999560
rect 365074 999504 365076 999524
rect 365076 999504 365128 999524
rect 365128 999504 365130 999524
rect 364706 999388 364762 999424
rect 364706 999368 364708 999388
rect 364708 999368 364760 999388
rect 364760 999368 364762 999388
rect 365442 999268 365444 999288
rect 365444 999268 365496 999288
rect 365496 999268 365498 999288
rect 365442 999232 365498 999268
rect 366178 993656 366234 993712
rect 368938 997192 368994 997248
rect 423494 1005372 423550 1005408
rect 423494 1005352 423496 1005372
rect 423496 1005352 423548 1005372
rect 423548 1005352 423550 1005372
rect 428370 1005252 428372 1005272
rect 428372 1005252 428424 1005272
rect 428424 1005252 428426 1005272
rect 428370 1005216 428426 1005252
rect 428830 1005100 428886 1005136
rect 428830 1005080 428832 1005100
rect 428832 1005080 428884 1005100
rect 428884 1005080 428886 1005100
rect 425518 1004980 425520 1005000
rect 425520 1004980 425572 1005000
rect 425572 1004980 425574 1005000
rect 425518 1004944 425574 1004980
rect 426806 1004964 426862 1005000
rect 426806 1004944 426808 1004964
rect 426808 1004944 426860 1004964
rect 426860 1004944 426862 1004964
rect 427174 1004844 427176 1004864
rect 427176 1004844 427228 1004864
rect 427228 1004844 427230 1004864
rect 427174 1004808 427230 1004844
rect 427542 1004828 427598 1004864
rect 427542 1004808 427544 1004828
rect 427544 1004808 427596 1004828
rect 427596 1004808 427598 1004828
rect 421838 1004708 421840 1004728
rect 421840 1004708 421892 1004728
rect 421892 1004708 421894 1004728
rect 383096 996376 383152 996432
rect 399942 997192 399998 997248
rect 388166 995696 388222 995752
rect 378138 993792 378194 993848
rect 375194 993656 375250 993712
rect 396998 993792 397054 993848
rect 395158 993656 395214 993712
rect 421838 1004672 421894 1004708
rect 422666 1004708 422668 1004728
rect 422668 1004708 422720 1004728
rect 422720 1004708 422722 1004728
rect 422666 1004672 422722 1004708
rect 425150 1004708 425152 1004728
rect 425152 1004708 425204 1004728
rect 425204 1004708 425206 1004728
rect 425150 1004672 425206 1004708
rect 426346 1000612 426402 1000648
rect 426346 1000592 426348 1000612
rect 426348 1000592 426400 1000612
rect 426400 1000592 426402 1000612
rect 428002 1000628 428004 1000648
rect 428004 1000628 428056 1000648
rect 428056 1000628 428058 1000648
rect 428002 1000592 428058 1000628
rect 425978 1000492 425980 1000512
rect 425980 1000492 426032 1000512
rect 426032 1000492 426034 1000512
rect 425978 1000456 426034 1000492
rect 430854 999812 430856 999832
rect 430856 999812 430908 999832
rect 430908 999812 430910 999832
rect 430854 999776 430910 999812
rect 431682 999796 431738 999832
rect 431682 999776 431684 999796
rect 431684 999776 431736 999796
rect 431736 999776 431738 999796
rect 429198 999676 429200 999696
rect 429200 999676 429252 999696
rect 429252 999676 429254 999696
rect 429198 999640 429254 999676
rect 430026 999660 430082 999696
rect 430026 999640 430028 999660
rect 430028 999640 430080 999660
rect 430080 999640 430082 999660
rect 431222 999540 431224 999560
rect 431224 999540 431276 999560
rect 431276 999540 431278 999560
rect 431222 999504 431278 999540
rect 432418 999524 432474 999560
rect 432418 999504 432420 999524
rect 432420 999504 432472 999524
rect 432472 999504 432474 999524
rect 429658 999388 429714 999424
rect 429658 999368 429660 999388
rect 429660 999368 429712 999388
rect 429712 999368 429714 999388
rect 432878 999404 432880 999424
rect 432880 999404 432932 999424
rect 432932 999404 432934 999424
rect 432878 999368 432934 999404
rect 430394 999268 430396 999288
rect 430396 999268 430448 999288
rect 430448 999268 430450 999288
rect 430394 999232 430450 999268
rect 432050 999252 432106 999288
rect 432050 999232 432052 999252
rect 432052 999232 432104 999252
rect 432104 999232 432106 999252
rect 437386 999096 437442 999152
rect 439822 997192 439878 997248
rect 502982 1005780 503038 1005816
rect 502982 1005760 502984 1005780
rect 502984 1005760 503036 1005780
rect 503036 1005760 503038 1005780
rect 503350 1005796 503352 1005816
rect 503352 1005796 503404 1005816
rect 503404 1005796 503406 1005816
rect 503350 1005760 503406 1005796
rect 502522 1005660 502524 1005680
rect 502524 1005660 502576 1005680
rect 502576 1005660 502578 1005680
rect 502522 1005624 502578 1005660
rect 504546 1005644 504602 1005680
rect 504546 1005624 504548 1005644
rect 504548 1005624 504600 1005644
rect 504600 1005624 504602 1005644
rect 505374 1005508 505430 1005544
rect 505374 1005488 505376 1005508
rect 505376 1005488 505428 1005508
rect 505428 1005488 505430 1005508
rect 505834 1005524 505836 1005544
rect 505836 1005524 505888 1005544
rect 505888 1005524 505890 1005544
rect 505834 1005488 505890 1005524
rect 447322 995696 447378 995752
rect 447138 993656 447194 993712
rect 504178 1005116 504180 1005136
rect 504180 1005116 504232 1005136
rect 504232 1005116 504234 1005136
rect 504178 1005080 504234 1005116
rect 505006 1004964 505062 1005000
rect 505006 1004944 505008 1004964
rect 505008 1004944 505060 1004964
rect 505060 1004944 505062 1004964
rect 500498 1004828 500554 1004864
rect 500498 1004808 500500 1004828
rect 500500 1004808 500552 1004828
rect 500552 1004808 500554 1004828
rect 498842 1004708 498844 1004728
rect 498844 1004708 498896 1004728
rect 498896 1004708 498898 1004728
rect 488906 997192 488962 997248
rect 481454 995696 481510 995752
rect 478602 993656 478658 993712
rect 485318 989440 485374 989496
rect 498842 1004672 498898 1004708
rect 499670 1004708 499672 1004728
rect 499672 1004708 499724 1004728
rect 499724 1004708 499726 1004728
rect 499670 1004672 499726 1004708
rect 501694 1004708 501696 1004728
rect 501696 1004708 501748 1004728
rect 501748 1004708 501750 1004728
rect 501694 1004672 501750 1004708
rect 502154 1004692 502210 1004728
rect 502154 1004672 502156 1004692
rect 502156 1004672 502208 1004692
rect 502208 1004672 502210 1004692
rect 508686 999796 508742 999832
rect 508686 999776 508688 999796
rect 508688 999776 508740 999796
rect 508740 999776 508742 999796
rect 506202 999676 506204 999696
rect 506204 999676 506256 999696
rect 506256 999676 506258 999696
rect 506202 999640 506258 999676
rect 508226 999660 508282 999696
rect 508226 999640 508228 999660
rect 508228 999640 508280 999660
rect 508280 999640 508282 999660
rect 507030 999540 507032 999560
rect 507032 999540 507084 999560
rect 507084 999540 507086 999560
rect 507030 999504 507086 999540
rect 507858 999524 507914 999560
rect 507858 999504 507860 999524
rect 507860 999504 507912 999524
rect 507912 999504 507914 999524
rect 506662 999404 506664 999424
rect 506664 999404 506716 999424
rect 506716 999404 506718 999424
rect 506662 999368 506718 999404
rect 509054 999388 509110 999424
rect 509054 999368 509056 999388
rect 509056 999368 509108 999388
rect 509108 999368 509110 999388
rect 500866 999252 500922 999288
rect 500866 999232 500868 999252
rect 500868 999232 500920 999252
rect 500920 999232 500922 999252
rect 507398 999268 507400 999288
rect 507400 999268 507452 999288
rect 507452 999268 507454 999288
rect 507398 999232 507454 999268
rect 503350 999132 503352 999152
rect 503352 999132 503404 999152
rect 503404 999132 503406 999152
rect 503350 999096 503406 999132
rect 509514 999252 509570 999288
rect 509514 999232 509516 999252
rect 509516 999232 509568 999252
rect 509568 999232 509570 999252
rect 509882 999132 509884 999152
rect 509884 999132 509936 999152
rect 509936 999132 509938 999152
rect 509882 999096 509938 999132
rect 513629 999096 513685 999152
rect 511446 989440 511502 989496
rect 517242 999096 517298 999152
rect 520002 999232 520058 999288
rect 520186 995696 520242 995752
rect 517610 995560 517666 995616
rect 551926 1005100 551982 1005136
rect 551926 1005080 551928 1005100
rect 551928 1005080 551980 1005100
rect 551980 1005080 551982 1005100
rect 554778 1004964 554834 1005000
rect 554778 1004944 554780 1004964
rect 554780 1004944 554832 1004964
rect 554832 1004944 554834 1004964
rect 520370 995424 520426 995480
rect 546406 1004672 546462 1004728
rect 549442 1004708 549444 1004728
rect 549444 1004708 549496 1004728
rect 549496 1004708 549498 1004728
rect 549442 1004672 549498 1004708
rect 550270 1004708 550272 1004728
rect 550272 1004708 550324 1004728
rect 550324 1004708 550326 1004728
rect 550270 1004672 550326 1004708
rect 551098 1004708 551100 1004728
rect 551100 1004708 551152 1004728
rect 551152 1004708 551154 1004728
rect 551098 1004672 551154 1004708
rect 523866 999232 523922 999288
rect 524050 999096 524106 999152
rect 523866 996512 523922 996568
rect 524050 996376 524106 996432
rect 525430 995696 525486 995752
rect 528006 995696 528062 995752
rect 528558 995696 528614 995752
rect 526074 995560 526130 995616
rect 532146 995424 532202 995480
rect 517426 993656 517482 993712
rect 537390 993656 537446 993712
rect 553122 1004844 553124 1004864
rect 553124 1004844 553176 1004864
rect 553176 1004844 553178 1004864
rect 553122 1004808 553178 1004844
rect 553950 1004828 554006 1004864
rect 553950 1004808 553952 1004828
rect 553952 1004808 554004 1004828
rect 554004 1004808 554006 1004828
rect 552754 1004708 552756 1004728
rect 552756 1004708 552808 1004728
rect 552808 1004708 552810 1004728
rect 552754 1004672 552810 1004708
rect 553490 1003484 553492 1003504
rect 553492 1003484 553544 1003504
rect 553544 1003484 553546 1003504
rect 553490 1003448 553546 1003484
rect 555146 1004672 555202 1004728
rect 567474 1004808 567530 1004864
rect 554318 1003212 554320 1003232
rect 554320 1003212 554372 1003232
rect 554372 1003212 554374 1003232
rect 554318 1003176 554374 1003212
rect 555974 1000068 556030 1000104
rect 555974 1000048 555976 1000068
rect 555976 1000048 556028 1000068
rect 556028 1000048 556030 1000068
rect 558458 999932 558514 999968
rect 558458 999912 558460 999932
rect 558460 999912 558512 999932
rect 558512 999912 558514 999932
rect 556342 999796 556398 999832
rect 556342 999776 556344 999796
rect 556344 999776 556396 999796
rect 556396 999776 556398 999796
rect 560850 999812 560852 999832
rect 560852 999812 560904 999832
rect 560904 999812 560906 999832
rect 560850 999776 560906 999812
rect 559194 999660 559250 999696
rect 559194 999640 559196 999660
rect 559196 999640 559248 999660
rect 559248 999640 559250 999660
rect 560482 999676 560484 999696
rect 560484 999676 560536 999696
rect 560536 999676 560538 999696
rect 560482 999640 560538 999676
rect 557998 999524 558054 999560
rect 557998 999504 558000 999524
rect 558000 999504 558052 999524
rect 558052 999504 558054 999524
rect 560022 999540 560024 999560
rect 560024 999540 560076 999560
rect 560076 999540 560078 999560
rect 560022 999504 560078 999540
rect 556802 999404 556804 999424
rect 556804 999404 556856 999424
rect 556856 999404 556858 999424
rect 556802 999368 556858 999404
rect 557170 999388 557226 999424
rect 557170 999368 557172 999388
rect 557172 999368 557224 999388
rect 557224 999368 557226 999388
rect 554318 999252 554374 999288
rect 554318 999232 554320 999252
rect 554320 999232 554372 999252
rect 554372 999232 554374 999252
rect 558826 999268 558828 999288
rect 558828 999268 558880 999288
rect 558880 999268 558882 999288
rect 558826 999232 558882 999268
rect 559654 999252 559710 999288
rect 559654 999232 559656 999252
rect 559656 999232 559708 999252
rect 559708 999232 559710 999252
rect 561310 999232 561366 999288
rect 551926 999132 551928 999152
rect 551928 999132 551980 999152
rect 551980 999132 551982 999152
rect 551926 999096 551982 999132
rect 557630 999132 557632 999152
rect 557632 999132 557684 999152
rect 557684 999132 557686 999152
rect 557630 999096 557686 999132
rect 561770 993656 561826 993712
rect 561034 985768 561090 985824
rect 561586 985768 561642 985824
rect 564438 985904 564494 985960
rect 567014 993688 567070 993744
rect 571338 994064 571394 994120
rect 569958 993792 570014 993848
rect 575570 994200 575626 994256
rect 629666 993928 629722 993984
rect 634818 994200 634874 994256
rect 638544 995152 638600 995208
rect 637026 994064 637082 994120
rect 635186 993792 635242 993848
rect 638866 993656 638922 993712
rect 641166 990528 641222 990584
rect 62854 814136 62910 814192
rect 62670 278160 62726 278216
rect 62486 278024 62542 278080
rect 63038 730224 63094 730280
rect 62946 427896 63002 427952
rect 62854 277888 62910 277944
rect 63130 684256 63186 684312
rect 63222 386688 63278 386744
rect 63314 383696 63370 383752
rect 63038 277752 63094 277808
rect 70582 271768 70638 271824
rect 69386 269048 69442 269104
rect 76470 271904 76526 271960
rect 78862 269320 78918 269376
rect 77666 269184 77722 269240
rect 83554 272040 83610 272096
rect 85946 272176 86002 272232
rect 87142 269592 87198 269648
rect 84750 269456 84806 269512
rect 91834 272312 91890 272368
rect 90638 269728 90694 269784
rect 97722 272720 97778 272776
rect 100114 272584 100170 272640
rect 98918 272448 98974 272504
rect 101310 270000 101366 270056
rect 96618 269864 96674 269920
rect 107198 272992 107254 273048
rect 106002 272856 106058 272912
rect 108394 270272 108450 270328
rect 103702 270136 103758 270192
rect 111982 273128 112038 273184
rect 115478 271632 115534 271688
rect 122562 271496 122618 271552
rect 121366 270408 121422 270464
rect 128542 268912 128598 268968
rect 127346 268776 127402 268832
rect 142710 268640 142766 268696
rect 153290 268504 153346 268560
rect 184938 268368 184994 268424
rect 194138 271768 194194 271824
rect 194506 271788 194562 271824
rect 194506 271768 194508 271788
rect 194508 271768 194560 271788
rect 194560 271768 194562 271788
rect 193678 269048 193734 269104
rect 196346 271904 196402 271960
rect 196806 269184 196862 269240
rect 199106 272040 199162 272096
rect 199934 272176 199990 272232
rect 199014 269456 199070 269512
rect 197726 269320 197782 269376
rect 200394 269592 200450 269648
rect 201314 272720 201370 272776
rect 202142 272312 202198 272368
rect 201682 269728 201738 269784
rect 203522 272992 203578 273048
rect 203062 268368 203118 268424
rect 204810 272448 204866 272504
rect 204350 269864 204406 269920
rect 203522 268096 203578 268152
rect 205730 272584 205786 272640
rect 205270 270000 205326 270056
rect 207478 272856 207534 272912
rect 207018 270136 207074 270192
rect 208490 271768 208546 271824
rect 207938 270272 207994 270328
rect 208398 268096 208454 268152
rect 209226 273128 209282 273184
rect 210606 271632 210662 271688
rect 213274 271496 213330 271552
rect 213734 270408 213790 270464
rect 215482 268776 215538 268832
rect 216402 268912 216458 268968
rect 221738 268640 221794 268696
rect 225786 268504 225842 268560
rect 353942 268232 353998 268288
rect 356610 268368 356666 268424
rect 358910 268640 358966 268696
rect 359370 268504 359426 268560
rect 362038 268776 362094 268832
rect 363326 271360 363382 271416
rect 364246 268912 364302 268968
rect 365994 271632 366050 271688
rect 365534 271496 365590 271552
rect 366914 270408 366970 270464
rect 368662 273128 368718 273184
rect 369582 270272 369638 270328
rect 371238 272992 371294 273048
rect 371330 272856 371386 272912
rect 372250 270136 372306 270192
rect 373998 272720 374054 272776
rect 378046 270000 378102 270056
rect 379334 272584 379390 272640
rect 383382 269864 383438 269920
rect 385130 266056 385186 266112
rect 386970 267552 387026 267608
rect 386510 266192 386566 266248
rect 388258 275848 388314 275904
rect 387798 267688 387854 267744
rect 389638 267416 389694 267472
rect 391294 275712 391350 275768
rect 390466 267280 390522 267336
rect 391386 269728 391442 269784
rect 392766 272448 392822 272504
rect 391846 267144 391902 267200
rect 393134 267008 393190 267064
rect 393594 275576 393650 275632
rect 394514 266872 394570 266928
rect 396262 275440 396318 275496
rect 395802 266736 395858 266792
rect 397182 266600 397238 266656
rect 398930 275304 398986 275360
rect 398102 272312 398158 272368
rect 398470 266464 398526 266520
rect 399850 266328 399906 266384
rect 401690 275168 401746 275224
rect 402702 274896 402758 274952
rect 402058 269592 402114 269648
rect 403438 272176 403494 272232
rect 404266 275032 404322 275088
rect 405462 274760 405518 274816
rect 404726 269456 404782 269512
rect 405646 265920 405702 265976
rect 406934 274624 406990 274680
rect 408222 274488 408278 274544
rect 407394 269320 407450 269376
rect 408314 265784 408370 265840
rect 408774 272040 408830 272096
rect 410522 271904 410578 271960
rect 409602 269184 409658 269240
rect 410062 269048 410118 269104
rect 410890 271768 410946 271824
rect 466274 265920 466330 265976
rect 459466 265784 459522 265840
rect 494978 268232 495034 268288
rect 502062 268368 502118 268424
rect 507950 268640 508006 268696
rect 509146 268504 509202 268560
rect 516230 268776 516286 268832
rect 519818 271360 519874 271416
rect 522210 268912 522266 268968
rect 526902 271632 526958 271688
rect 525706 271496 525762 271552
rect 529294 270408 529350 270464
rect 533986 273128 534042 273184
rect 536378 270272 536434 270328
rect 539874 272992 539930 273048
rect 541070 272856 541126 272912
rect 543462 270136 543518 270192
rect 548154 272720 548210 272776
rect 558826 270000 558882 270056
rect 562414 272584 562470 272640
rect 572994 269864 573050 269920
rect 586058 275848 586114 275904
rect 584862 267688 584918 267744
rect 582470 267552 582526 267608
rect 589554 267416 589610 267472
rect 593142 275712 593198 275768
rect 594338 269728 594394 269784
rect 591946 267280 592002 267336
rect 595442 267144 595498 267200
rect 597834 272448 597890 272504
rect 600226 275576 600282 275632
rect 599030 267008 599086 267064
rect 602526 266872 602582 266928
rect 607310 275440 607366 275496
rect 606114 266736 606170 266792
rect 612002 272312 612058 272368
rect 609702 266600 609758 266656
rect 614394 275304 614450 275360
rect 613198 266464 613254 266520
rect 621478 275168 621534 275224
rect 623870 274896 623926 274952
rect 628562 275032 628618 275088
rect 626170 272176 626226 272232
rect 622674 269592 622730 269648
rect 630954 274760 631010 274816
rect 635646 274624 635702 274680
rect 629758 269456 629814 269512
rect 638038 274488 638094 274544
rect 640430 272040 640486 272096
rect 636842 269320 636898 269376
rect 642730 269184 642786 269240
rect 645122 271904 645178 271960
rect 646318 271768 646374 271824
rect 643926 269048 643982 269104
rect 616786 266328 616842 266384
rect 581274 266192 581330 266248
rect 577778 266056 577834 266112
rect 416778 262268 416834 262304
rect 416778 262248 416780 262268
rect 416780 262248 416832 262268
rect 416832 262248 416834 262268
rect 416778 259120 416834 259176
rect 184938 258576 184994 258632
rect 416778 255856 416834 255912
rect 416778 252728 416834 252784
rect 416778 249464 416834 249520
rect 184938 247968 184994 248024
rect 416778 246336 416834 246392
rect 418066 243072 418122 243128
rect 184938 237396 184940 237416
rect 184940 237396 184992 237416
rect 184992 237396 184994 237416
rect 184938 237360 184994 237396
rect 93030 228928 93086 228984
rect 84658 228792 84714 228848
rect 82726 228384 82782 228440
rect 76286 228248 76342 228304
rect 71226 228112 71282 228168
rect 69478 227976 69534 228032
rect 62762 227840 62818 227896
rect 61106 222264 61162 222320
rect 63406 225120 63462 225176
rect 66994 225256 67050 225312
rect 67822 222400 67878 222456
rect 70398 225392 70454 225448
rect 72882 222672 72938 222728
rect 74446 222536 74502 222592
rect 77114 225528 77170 225584
rect 80426 225800 80482 225856
rect 79598 222808 79654 222864
rect 81254 222944 81310 223000
rect 83830 225664 83886 225720
rect 86314 228656 86370 228712
rect 88062 228520 88118 228576
rect 92202 225936 92258 225992
rect 89718 223080 89774 223136
rect 94778 227432 94834 227488
rect 101494 227296 101550 227352
rect 99838 227160 99894 227216
rect 98918 226208 98974 226264
rect 97262 224712 97318 224768
rect 96434 223216 96490 223272
rect 98090 223352 98146 223408
rect 106554 227024 106610 227080
rect 102046 226072 102102 226128
rect 103150 221992 103206 222048
rect 104806 223488 104862 223544
rect 113086 226888 113142 226944
rect 109038 224576 109094 224632
rect 112442 224440 112498 224496
rect 110694 224168 110750 224224
rect 109866 221856 109922 221912
rect 111614 221720 111670 221776
rect 114926 226752 114982 226808
rect 115754 224304 115810 224360
rect 118330 221448 118386 221504
rect 120814 224032 120870 224088
rect 121366 221584 121422 221640
rect 192574 224984 192630 225040
rect 193678 224848 193734 224904
rect 193310 222128 193366 222184
rect 194782 227704 194838 227760
rect 194414 227568 194470 227624
rect 197266 227840 197322 227896
rect 196530 225120 196586 225176
rect 196162 222264 196218 222320
rect 198002 225256 198058 225312
rect 198738 222400 198794 222456
rect 200486 228112 200542 228168
rect 200118 227976 200174 228032
rect 199382 225392 199438 225448
rect 201498 222672 201554 222728
rect 202970 228248 203026 228304
rect 202234 225528 202290 225584
rect 201866 222536 201922 222592
rect 203706 225800 203762 225856
rect 205086 225664 205142 225720
rect 204718 222944 204774 223000
rect 204350 222808 204406 222864
rect 206190 228792 206246 228848
rect 205822 228384 205878 228440
rect 207202 228656 207258 228712
rect 207570 228520 207626 228576
rect 208306 225936 208362 225992
rect 208674 223080 208730 223136
rect 210054 228928 210110 228984
rect 210422 227432 210478 227488
rect 210790 227704 210846 227760
rect 210514 224712 210570 224768
rect 211158 226208 211214 226264
rect 211526 223216 211582 223272
rect 212354 227568 212410 227624
rect 211894 223352 211950 223408
rect 213274 227296 213330 227352
rect 212906 227160 212962 227216
rect 212538 226072 212594 226128
rect 214470 223488 214526 223544
rect 214378 221992 214434 222048
rect 215758 227024 215814 227080
rect 215390 224576 215446 224632
rect 216494 224168 216550 224224
rect 216862 224440 216918 224496
rect 217230 221856 217286 221912
rect 217598 227840 217654 227896
rect 217322 221720 217378 221776
rect 218610 226888 218666 226944
rect 219254 227976 219310 228032
rect 218978 226752 219034 226808
rect 218242 224304 218298 224360
rect 220726 228112 220782 228168
rect 220450 221448 220506 221504
rect 220818 224032 220874 224088
rect 221830 221584 221886 221640
rect 225970 228248 226026 228304
rect 235538 228384 235594 228440
rect 237102 228520 237158 228576
rect 246946 228792 247002 228848
rect 256698 228928 256754 228984
rect 259642 228520 259698 228576
rect 260010 227704 260066 227760
rect 260378 227568 260434 227624
rect 261758 228928 261814 228984
rect 261390 228792 261446 228848
rect 262494 228384 262550 228440
rect 263230 227976 263286 228032
rect 262862 227840 262918 227896
rect 264242 228112 264298 228168
rect 266082 228248 266138 228304
rect 330942 222808 330998 222864
rect 332690 222944 332746 223000
rect 332322 222536 332378 222592
rect 333794 222400 333850 222456
rect 335818 222672 335874 222728
rect 335910 222128 335966 222184
rect 338762 222264 338818 222320
rect 369398 224440 369454 224496
rect 370870 224576 370926 224632
rect 372250 226208 372306 226264
rect 373722 224712 373778 224768
rect 375102 221992 375158 222048
rect 375838 227160 375894 227216
rect 376942 223488 376998 223544
rect 377310 223352 377366 223408
rect 378322 227296 378378 227352
rect 379794 223216 379850 223272
rect 380162 223080 380218 223136
rect 381542 228792 381598 228848
rect 381174 227432 381230 227488
rect 381082 222808 381138 222864
rect 381818 222944 381874 223000
rect 382646 222808 382702 222864
rect 383658 228928 383714 228984
rect 384302 222536 384358 222592
rect 384762 222944 384818 223000
rect 385866 228656 385922 228712
rect 387982 228520 388038 228576
rect 389086 228384 389142 228440
rect 388534 222672 388590 222728
rect 387706 222400 387762 222456
rect 386878 221720 386934 221776
rect 391202 228248 391258 228304
rect 390466 225664 390522 225720
rect 391570 225392 391626 225448
rect 390098 222672 390154 222728
rect 390190 222128 390246 222184
rect 393318 228112 393374 228168
rect 392582 225528 392638 225584
rect 392214 222536 392270 222592
rect 394422 222128 394478 222184
rect 395434 227840 395490 227896
rect 395986 224304 396042 224360
rect 397642 227976 397698 228032
rect 396538 222400 396594 222456
rect 396906 222264 396962 222320
rect 397918 225256 397974 225312
rect 400126 225120 400182 225176
rect 397458 221856 397514 221912
rect 402978 227704 403034 227760
rect 403346 224984 403402 225040
rect 405094 227568 405150 227624
rect 404358 224848 404414 224904
rect 408314 226072 408370 226128
rect 408406 225936 408462 225992
rect 410062 227024 410118 227080
rect 409786 222672 409842 222728
rect 411166 225800 411222 225856
rect 409786 221720 409842 221776
rect 418158 239944 418214 240000
rect 418434 236680 418490 236736
rect 418526 233552 418582 233608
rect 471978 224440 472034 224496
rect 478510 226208 478566 226264
rect 475106 224576 475162 224632
rect 486054 227160 486110 227216
rect 481914 224712 481970 224768
rect 480258 224304 480314 224360
rect 483570 221992 483626 222048
rect 504546 228928 504602 228984
rect 499670 228792 499726 228848
rect 496818 227432 496874 227488
rect 492310 227296 492366 227352
rect 488630 223488 488686 223544
rect 489458 223352 489514 223408
rect 488630 221176 488686 221232
rect 491390 221856 491446 221912
rect 491390 220904 491446 220960
rect 495346 223216 495402 223272
rect 494058 223080 494114 223136
rect 494058 221040 494114 221096
rect 493046 220904 493102 220960
rect 496818 221312 496874 221368
rect 496450 221040 496506 221096
rect 499302 221312 499358 221368
rect 502706 222808 502762 222864
rect 502706 221584 502762 221640
rect 509882 228656 509938 228712
rect 507122 222944 507178 223000
rect 507122 221448 507178 221504
rect 514666 228520 514722 228576
rect 513470 226072 513526 226128
rect 510618 222672 510674 222728
rect 510618 221720 510674 221776
rect 512458 221720 512514 221776
rect 516138 227024 516194 227080
rect 517242 228384 517298 228440
rect 518714 225936 518770 225992
rect 522486 228248 522542 228304
rect 520830 225664 520886 225720
rect 519726 222536 519782 222592
rect 527546 228112 527602 228168
rect 525798 225528 525854 225584
rect 523406 225392 523462 225448
rect 522486 221856 522542 221912
rect 525062 222400 525118 222456
rect 535458 227976 535514 228032
rect 532698 227840 532754 227896
rect 530674 225800 530730 225856
rect 529938 222128 529994 222184
rect 534906 222264 534962 222320
rect 538862 225256 538918 225312
rect 543554 225120 543610 225176
rect 550270 227704 550326 227760
rect 549350 224984 549406 225040
rect 552018 224848 552074 224904
rect 555054 227568 555110 227624
rect 580170 216144 580226 216200
rect 582286 214648 582342 214704
rect 580262 213152 580318 213208
rect 581642 211656 581698 211712
rect 580538 210160 580594 210216
rect 579710 208664 579766 208720
rect 582286 207052 582342 207088
rect 582286 207032 582288 207052
rect 582288 207032 582340 207052
rect 582340 207032 582342 207052
rect 582286 205536 582342 205592
rect 599766 209480 599822 209536
rect 627090 221856 627146 221912
rect 625250 221720 625306 221776
rect 623410 221584 623466 221640
rect 622950 221312 623006 221368
rect 621478 221176 621534 221232
rect 624330 221448 624386 221504
rect 637394 221040 637450 221096
rect 636934 220904 636990 220960
rect 654874 922664 654930 922720
rect 654874 909472 654930 909528
rect 654874 896144 654930 896200
rect 655150 882816 655206 882872
rect 654690 856296 654746 856352
rect 655058 842968 655114 843024
rect 654138 816448 654194 816504
rect 655058 789928 655114 789984
rect 654782 763272 654838 763328
rect 654874 750080 654930 750136
rect 654782 736752 654838 736808
rect 654690 696904 654746 696960
rect 654874 683576 654930 683632
rect 654874 643728 654930 643784
rect 655058 630536 655114 630592
rect 654598 617208 654654 617264
rect 654322 603880 654378 603936
rect 655058 577360 655114 577416
rect 654322 564032 654378 564088
rect 654690 550840 654746 550896
rect 654874 537512 654930 537568
rect 654138 524184 654194 524240
rect 654874 510992 654930 511048
rect 654874 484336 654930 484392
rect 654874 471144 654930 471200
rect 654230 457816 654286 457872
rect 654414 444508 654470 444544
rect 654414 444488 654416 444508
rect 654416 444488 654468 444508
rect 654468 444488 654470 444508
rect 654690 431296 654746 431352
rect 655058 417968 655114 418024
rect 654874 404640 654930 404696
rect 654322 391448 654378 391504
rect 654874 351600 654930 351656
rect 655058 338272 655114 338328
rect 654874 324944 654930 325000
rect 654138 311752 654194 311808
rect 655518 975840 655574 975896
rect 655702 962512 655758 962568
rect 655794 949320 655850 949376
rect 655610 936128 655666 936184
rect 656806 869644 656862 869680
rect 656806 869624 656808 869644
rect 656808 869624 656860 869644
rect 656860 869624 656862 869644
rect 655518 829776 655574 829832
rect 656806 803276 656862 803312
rect 656806 803256 656808 803276
rect 656808 803256 656860 803276
rect 656860 803256 656862 803276
rect 655518 776600 655574 776656
rect 655518 723424 655574 723480
rect 655978 710232 656034 710288
rect 655518 670384 655574 670440
rect 656162 657076 656218 657112
rect 656162 657056 656164 657076
rect 656164 657056 656216 657076
rect 656216 657056 656218 657076
rect 656806 590708 656862 590744
rect 656806 590688 656808 590708
rect 656808 590688 656860 590708
rect 656860 590688 656862 590708
rect 656806 497684 656862 497720
rect 656806 497664 656808 497684
rect 656808 497664 656860 497684
rect 656860 497664 656862 497684
rect 656806 378156 656808 378176
rect 656808 378156 656860 378176
rect 656860 378156 656862 378176
rect 656806 378120 656862 378156
rect 656806 364792 656862 364848
rect 655610 298424 655666 298480
rect 655334 285232 655390 285288
rect 658186 262384 658242 262440
rect 599950 208528 600006 208584
rect 599858 207440 599914 207496
rect 600042 206488 600098 206544
rect 599122 205400 599178 205456
rect 580722 204040 580778 204096
rect 581090 202544 581146 202600
rect 601514 204448 601570 204504
rect 601422 203360 601478 203416
rect 599950 202408 600006 202464
rect 598938 201320 598994 201376
rect 581090 201048 581146 201104
rect 599950 200368 600006 200424
rect 582286 199552 582342 199608
rect 599950 199280 600006 199336
rect 599122 198328 599178 198384
rect 582286 197920 582342 197976
rect 580722 196424 580778 196480
rect 599950 197276 599952 197296
rect 599952 197276 600004 197296
rect 600004 197276 600006 197296
rect 599950 197240 600006 197276
rect 599858 196288 599914 196344
rect 599950 195200 600006 195256
rect 582286 194928 582342 194984
rect 599122 194248 599178 194304
rect 582194 193432 582250 193488
rect 599950 193160 600006 193216
rect 599122 192208 599178 192264
rect 582286 191936 582342 191992
rect 599858 191120 599914 191176
rect 582194 190440 582250 190496
rect 600962 190168 601018 190224
rect 579802 188808 579858 188864
rect 601606 189080 601662 189136
rect 601422 188128 601478 188184
rect 582286 187312 582342 187368
rect 599950 187040 600006 187096
rect 582194 185816 582250 185872
rect 599858 185000 599914 185056
rect 580906 184320 580962 184376
rect 599766 184048 599822 184104
rect 580262 182824 580318 182880
rect 580630 181328 580686 181384
rect 580538 179696 580594 179752
rect 600042 186088 600098 186144
rect 599950 182960 600006 183016
rect 599858 179968 599914 180024
rect 599674 178880 599730 178936
rect 581090 178200 581146 178256
rect 598938 176840 598994 176896
rect 580722 176704 580778 176760
rect 579710 172216 579766 172272
rect 580538 170584 580594 170640
rect 579894 161472 579950 161528
rect 579710 158480 579766 158536
rect 580170 156984 580226 157040
rect 581458 175208 581514 175264
rect 582286 173748 582288 173768
rect 582288 173748 582340 173768
rect 582340 173748 582342 173768
rect 582286 173712 582342 173748
rect 582010 169088 582066 169144
rect 580998 167592 581054 167648
rect 580814 164600 580870 164656
rect 580354 152360 580410 152416
rect 580538 146376 580594 146432
rect 579710 122032 579766 122088
rect 579802 112920 579858 112976
rect 579894 108432 579950 108488
rect 580078 111424 580134 111480
rect 580170 106800 580226 106856
rect 579986 105304 580042 105360
rect 580262 102312 580318 102368
rect 580354 100816 580410 100872
rect 580814 141752 580870 141808
rect 580998 147872 581054 147928
rect 581826 163104 581882 163160
rect 581274 153992 581330 154048
rect 581458 149368 581514 149424
rect 581182 144880 581238 144936
rect 581090 143248 581146 143304
rect 580906 140256 580962 140312
rect 580722 138760 580778 138816
rect 580630 128152 580686 128208
rect 580538 97688 580594 97744
rect 580446 96192 580502 96248
rect 187606 41792 187662 41848
rect 194414 41792 194470 41848
rect 209778 41248 209834 41304
rect 212446 41248 212502 41304
rect 281446 48184 281502 48240
rect 230570 12144 230626 12200
rect 230938 16632 230994 16688
rect 230846 15136 230902 15192
rect 230754 13640 230810 13696
rect 230662 10648 230718 10704
rect 230478 9152 230534 9208
rect 230386 7656 230442 7712
rect 307298 41792 307354 41848
rect 362038 41792 362094 41848
rect 415490 41792 415546 41848
rect 470052 41928 470108 41984
rect 518806 44240 518862 44296
rect 520462 42064 520518 42120
rect 526166 44104 526222 44160
rect 552018 41792 552074 41848
rect 580722 99320 580778 99376
rect 580998 115912 581054 115968
rect 580906 103808 580962 103864
rect 580814 94696 580870 94752
rect 580630 93200 580686 93256
rect 579618 82628 579620 82648
rect 579620 82628 579672 82648
rect 579672 82628 579674 82648
rect 579618 82592 579674 82628
rect 580538 65864 580594 65920
rect 579618 59744 579674 59800
rect 579618 58248 579674 58304
rect 581366 126656 581422 126712
rect 581550 125024 581606 125080
rect 581458 123528 581514 123584
rect 581274 120536 581330 120592
rect 581182 114416 581238 114472
rect 581090 109928 581146 109984
rect 580998 70352 581054 70408
rect 581274 77968 581330 78024
rect 581918 150864 581974 150920
rect 581826 131144 581882 131200
rect 599766 177928 599822 177984
rect 600042 182008 600098 182064
rect 600134 180920 600190 180976
rect 599950 174800 600006 174856
rect 600318 175888 600374 175944
rect 599858 172760 599914 172816
rect 599950 171808 600006 171864
rect 599950 170720 600006 170776
rect 599766 169768 599822 169824
rect 599030 168680 599086 168736
rect 601146 173848 601202 173904
rect 599858 167728 599914 167784
rect 582286 166096 582342 166152
rect 600042 166640 600098 166696
rect 599950 165688 600006 165744
rect 599858 164600 599914 164656
rect 599950 163648 600006 163704
rect 599858 162560 599914 162616
rect 600042 161608 600098 161664
rect 599950 160520 600006 160576
rect 582194 159976 582250 160032
rect 598938 159568 598994 159624
rect 599858 158480 599914 158536
rect 599950 157548 600006 157584
rect 599950 157528 599952 157548
rect 599952 157528 600004 157548
rect 600004 157528 600006 157548
rect 599858 156440 599914 156496
rect 582102 155488 582158 155544
rect 582010 137264 582066 137320
rect 599950 155488 600006 155544
rect 600042 154400 600098 154456
rect 599858 153448 599914 153504
rect 599950 152360 600006 152416
rect 582194 135768 582250 135824
rect 582102 134136 582158 134192
rect 598938 151408 598994 151464
rect 599858 150320 599914 150376
rect 599950 149368 600006 149424
rect 599858 148280 599914 148336
rect 599950 147328 600006 147384
rect 600042 146240 600098 146296
rect 599858 145288 599914 145344
rect 599950 144200 600006 144256
rect 599858 143248 599914 143304
rect 599306 141208 599362 141264
rect 599950 142160 600006 142216
rect 599858 140120 599914 140176
rect 599766 139168 599822 139224
rect 599950 138116 599952 138136
rect 599952 138116 600004 138136
rect 600004 138116 600006 138136
rect 599950 138080 600006 138116
rect 599858 137128 599914 137184
rect 599950 136040 600006 136096
rect 600042 135088 600098 135144
rect 599858 134000 599914 134056
rect 582286 132640 582342 132696
rect 599950 133048 600006 133104
rect 599858 131960 599914 132016
rect 599766 131008 599822 131064
rect 599950 129920 600006 129976
rect 581918 129648 581974 129704
rect 599858 128968 599914 129024
rect 599950 127880 600006 127936
rect 599766 126928 599822 126984
rect 581734 119040 581790 119096
rect 581642 117544 581698 117600
rect 581550 81096 581606 81152
rect 581458 76472 581514 76528
rect 582010 90208 582066 90264
rect 600042 125840 600098 125896
rect 599950 124888 600006 124944
rect 600042 123800 600098 123856
rect 599858 122848 599914 122904
rect 599950 121760 600006 121816
rect 600042 120808 600098 120864
rect 599950 119720 600006 119776
rect 582286 91704 582342 91760
rect 582194 88576 582250 88632
rect 582102 87080 582158 87136
rect 581918 85584 581974 85640
rect 581826 84088 581882 84144
rect 581734 79464 581790 79520
rect 581642 74976 581698 75032
rect 581366 71984 581422 72040
rect 581182 67360 581238 67416
rect 581090 64368 581146 64424
rect 582010 62872 582066 62928
rect 581918 56752 581974 56808
rect 599858 118768 599914 118824
rect 599858 117680 599914 117736
rect 599950 116728 600006 116784
rect 599858 115640 599914 115696
rect 599950 114688 600006 114744
rect 599950 112648 600006 112704
rect 599766 111560 599822 111616
rect 600226 110608 600282 110664
rect 599950 109520 600006 109576
rect 599950 107480 600006 107536
rect 599950 100408 600006 100464
rect 582286 68856 582342 68912
rect 582194 61240 582250 61296
rect 600318 108568 600374 108624
rect 600594 106528 600650 106584
rect 600410 105440 600466 105496
rect 600502 103400 600558 103456
rect 600686 104488 600742 104544
rect 600870 102448 600926 102504
rect 600778 101360 600834 101416
rect 582102 55256 582158 55312
rect 580906 53760 580962 53816
rect 571338 41928 571394 41984
rect 563610 41656 563666 41712
rect 622122 85992 622178 86048
rect 623134 88848 623190 88904
rect 623226 87896 623282 87952
rect 622674 85040 622730 85096
rect 621938 84088 621994 84144
rect 623778 90616 623834 90672
rect 628286 95920 628342 95976
rect 640522 95684 640524 95704
rect 640524 95684 640576 95704
rect 640576 95684 640578 95704
rect 640522 95648 640578 95684
rect 627918 94424 627974 94480
rect 627274 93472 627330 93528
rect 626446 92520 626502 92576
rect 625894 91568 625950 91624
rect 623962 89664 624018 89720
rect 623502 86944 623558 87000
rect 623318 83136 623374 83192
rect 622306 82184 622362 82240
rect 622490 81368 622546 81424
rect 642730 92656 642786 92712
rect 645950 89664 646006 89720
rect 646042 87080 646098 87136
rect 652758 92520 652814 92576
rect 655334 93336 655390 93392
rect 654046 91432 654102 91488
rect 652942 90616 652998 90672
rect 656990 90344 657046 90400
rect 662234 95512 662290 95568
rect 657358 94696 657414 94752
rect 663246 93744 663302 93800
rect 663338 93064 663394 93120
rect 663430 92248 663486 92304
rect 663246 91024 663302 91080
rect 663430 89528 663486 89584
rect 663706 90344 663762 90400
rect 662142 88712 662198 88768
rect 646134 84632 646190 84688
rect 645858 82184 645914 82240
rect 661130 47504 661186 47560
rect 666650 183776 666706 183832
rect 666650 180376 666706 180432
rect 666650 178744 666706 178800
rect 669134 985632 669190 985688
rect 669042 983048 669098 983104
rect 666650 175344 666706 175400
rect 666650 173576 666706 173632
rect 666650 170176 666706 170232
rect 666650 168544 666706 168600
rect 666650 165144 666706 165200
rect 666650 163512 666706 163568
rect 666650 160112 666706 160168
rect 666650 158344 666706 158400
rect 666650 154944 666706 155000
rect 666650 153312 666706 153368
rect 666650 149912 666706 149968
rect 666650 148144 666706 148200
rect 666650 144880 666706 144936
rect 666650 143112 666706 143168
rect 666650 139712 666706 139768
rect 666650 132912 666706 132968
rect 670422 985496 670478 985552
rect 669778 759056 669834 759112
rect 672538 985360 672594 985416
rect 670422 621560 670478 621616
rect 670422 619520 670478 619576
rect 671066 209208 671122 209264
rect 671066 205808 671122 205864
rect 670974 204176 671030 204232
rect 670974 200776 671030 200832
rect 670882 199008 670938 199064
rect 670882 195608 670938 195664
rect 670790 193976 670846 194032
rect 670790 190576 670846 190632
rect 670698 188944 670754 189000
rect 670698 185544 670754 185600
rect 670698 138080 670754 138136
rect 670698 134680 670754 134736
rect 666650 129512 666706 129568
rect 666650 127880 666706 127936
rect 666650 124480 666706 124536
rect 666650 122848 666706 122904
rect 666650 119448 666706 119504
rect 670790 104080 670846 104136
rect 671802 173576 671858 173632
rect 672078 183776 672134 183832
rect 672170 178744 672226 178800
rect 671618 110880 671674 110936
rect 671158 107480 671214 107536
rect 672354 168544 672410 168600
rect 672170 117680 672226 117736
rect 672078 114280 672134 114336
rect 672630 982912 672686 982968
rect 675666 938712 675722 938768
rect 676310 939664 676366 939720
rect 676126 939256 676182 939312
rect 676218 938868 676274 938904
rect 676218 938848 676220 938868
rect 676220 938848 676272 938868
rect 676272 938848 676274 938868
rect 678978 937624 679034 937680
rect 676218 936400 676274 936456
rect 676034 935856 676090 935912
rect 675942 935468 675998 935504
rect 675942 935448 675944 935468
rect 675944 935448 675996 935468
rect 675996 935448 675998 935468
rect 675850 934632 675906 934688
rect 676034 935040 676090 935096
rect 675942 934224 675998 934280
rect 676126 933952 676182 934008
rect 676034 933408 676090 933464
rect 675758 933000 675814 933056
rect 676126 932764 676128 932784
rect 676128 932764 676180 932784
rect 676180 932764 676182 932784
rect 676126 932728 676182 932764
rect 676126 932320 676182 932376
rect 676034 931776 676090 931832
rect 676034 931368 676090 931424
rect 675942 930960 675998 931016
rect 676126 930688 676182 930744
rect 676034 930144 676090 930200
rect 678978 929464 679034 929520
rect 678978 928648 679034 928704
rect 675758 877240 675814 877296
rect 675666 876560 675722 876616
rect 675482 875880 675538 875936
rect 675390 873976 675446 874032
rect 673550 760280 673606 760336
rect 673550 759056 673606 759112
rect 675758 872208 675814 872264
rect 674286 797680 674342 797736
rect 674194 791968 674250 792024
rect 674378 777416 674434 777472
rect 675390 787752 675446 787808
rect 675390 787208 675446 787264
rect 675390 786800 675446 786856
rect 675390 784080 675446 784136
rect 675482 783808 675538 783864
rect 673826 699760 673882 699816
rect 673734 699488 673790 699544
rect 672446 163512 672502 163568
rect 675574 754160 675630 754216
rect 675482 744096 675538 744152
rect 675758 773336 675814 773392
rect 679070 772656 679126 772712
rect 678978 761232 679034 761288
rect 676218 760824 676274 760880
rect 676126 760416 676182 760472
rect 676310 759600 676366 759656
rect 676034 759092 676036 759112
rect 676036 759092 676088 759112
rect 676088 759092 676090 759112
rect 676034 759056 676090 759092
rect 679070 759600 679126 759656
rect 678978 758376 679034 758432
rect 676310 757968 676366 758024
rect 676126 757560 676182 757616
rect 676034 756608 676090 756664
rect 676218 757152 676274 757208
rect 676126 755520 676182 755576
rect 676034 754976 676090 755032
rect 675758 753752 675814 753808
rect 676034 753344 676090 753400
rect 676034 752936 676090 752992
rect 678978 751032 679034 751088
rect 678978 750216 679034 750272
rect 675666 743960 675722 744016
rect 675758 742872 675814 742928
rect 675758 742464 675814 742520
rect 675482 741648 675538 741704
rect 675390 739744 675446 739800
rect 675390 739064 675446 739120
rect 675666 738520 675722 738576
rect 675758 737976 675814 738032
rect 674010 699624 674066 699680
rect 672538 158344 672594 158400
rect 672630 153312 672686 153368
rect 676034 716488 676090 716544
rect 675942 716116 675944 716136
rect 675944 716116 675996 716136
rect 675996 716116 675998 716136
rect 675942 716080 675998 716116
rect 675942 715708 675944 715728
rect 675944 715708 675996 715728
rect 675996 715708 675998 715728
rect 675942 715672 675998 715708
rect 675942 715300 675944 715320
rect 675944 715300 675996 715320
rect 675996 715300 675998 715320
rect 675942 715264 675998 715300
rect 676034 714876 676090 714912
rect 676034 714856 676036 714876
rect 676036 714856 676088 714876
rect 676088 714856 676090 714876
rect 678978 714448 679034 714504
rect 676034 714060 676090 714096
rect 676034 714040 676036 714060
rect 676036 714040 676088 714060
rect 676088 714040 676090 714060
rect 676034 713668 676036 713688
rect 676036 713668 676088 713688
rect 676088 713668 676090 713688
rect 676034 713632 676090 713668
rect 676034 713244 676090 713280
rect 676034 713224 676036 713244
rect 676036 713224 676088 713244
rect 676088 713224 676090 713244
rect 676034 712836 676090 712872
rect 676034 712816 676036 712836
rect 676036 712816 676088 712836
rect 676088 712816 676090 712836
rect 676034 712428 676090 712464
rect 676034 712408 676036 712428
rect 676036 712408 676088 712428
rect 676088 712408 676090 712428
rect 675758 711592 675814 711648
rect 675850 710776 675906 710832
rect 675942 710368 675998 710424
rect 676310 711830 676366 711886
rect 676954 711830 677010 711886
rect 676034 709960 676090 710016
rect 676034 708328 676090 708384
rect 676034 707920 676090 707976
rect 676034 707512 676090 707568
rect 676310 707104 676366 707160
rect 676034 706696 676090 706752
rect 676034 706288 676090 706344
rect 676034 705100 676036 705120
rect 676036 705100 676088 705120
rect 676088 705100 676090 705120
rect 676034 705064 676090 705100
rect 675482 698128 675538 698184
rect 675390 697176 675446 697232
rect 675390 696632 675446 696688
rect 675390 695000 675446 695056
rect 675482 694184 675538 694240
rect 675390 693640 675446 693696
rect 675758 692960 675814 693016
rect 675758 690104 675814 690160
rect 676218 671508 676220 671528
rect 676220 671508 676272 671528
rect 676272 671508 676274 671528
rect 676218 671472 676274 671508
rect 676034 670928 676090 670984
rect 676034 670556 676036 670576
rect 676036 670556 676088 670576
rect 676088 670556 676090 670576
rect 676034 670520 676090 670556
rect 676218 670284 676220 670304
rect 676220 670284 676272 670304
rect 676272 670284 676274 670304
rect 676218 670248 676274 670284
rect 676034 669740 676036 669760
rect 676036 669740 676088 669760
rect 676088 669740 676090 669760
rect 676034 669704 676090 669740
rect 678978 669432 679034 669488
rect 676034 668888 676090 668944
rect 675942 668092 675998 668128
rect 675942 668072 675944 668092
rect 675944 668072 675996 668092
rect 675996 668072 675998 668092
rect 676218 668652 676220 668672
rect 676220 668652 676272 668672
rect 676272 668652 676274 668672
rect 676218 668616 676274 668652
rect 675942 667700 675944 667720
rect 675944 667700 675996 667720
rect 675996 667700 675998 667720
rect 675942 667664 675998 667700
rect 676126 666576 676182 666632
rect 676034 665216 676090 665272
rect 676034 664808 676090 664864
rect 676034 663176 676090 663232
rect 678978 660864 679034 660920
rect 678978 660048 679034 660104
rect 675390 652568 675446 652624
rect 675482 652160 675538 652216
rect 675390 651616 675446 651672
rect 675758 649168 675814 649224
rect 675666 648624 675722 648680
rect 674378 607688 674434 607744
rect 678978 626048 679034 626104
rect 676218 625640 676274 625696
rect 676034 625096 676090 625152
rect 676126 624416 676182 624472
rect 676034 623908 676036 623928
rect 676036 623908 676088 623928
rect 676088 623908 676090 623928
rect 676034 623872 676090 623908
rect 676310 625232 676366 625288
rect 679070 624416 679126 624472
rect 679162 623600 679218 623656
rect 678978 623192 679034 623248
rect 676218 621968 676274 622024
rect 676034 621424 676090 621480
rect 676126 620336 676182 620392
rect 676034 619792 676090 619848
rect 676034 618196 676036 618216
rect 676036 618196 676088 618216
rect 676088 618196 676090 618216
rect 676034 618160 676090 618196
rect 676218 617924 676220 617944
rect 676220 617924 676272 617944
rect 676272 617924 676274 617944
rect 676218 617888 676274 617924
rect 676218 616700 676220 616720
rect 676220 616700 676272 616720
rect 676272 616700 676274 616720
rect 676218 616664 676274 616700
rect 678978 615848 679034 615904
rect 678978 615032 679034 615088
rect 675482 607552 675538 607608
rect 674746 607416 674802 607472
rect 675758 607280 675814 607336
rect 675390 606464 675446 606520
rect 675390 604696 675446 604752
rect 675390 604288 675446 604344
rect 675482 603472 675538 603528
rect 675758 602928 675814 602984
rect 674654 564440 674710 564496
rect 676310 580896 676366 580952
rect 676126 580488 676182 580544
rect 676218 580080 676274 580136
rect 676034 579808 676090 579864
rect 676218 579284 676274 579320
rect 676218 579264 676220 579284
rect 676220 579264 676272 579284
rect 676272 579264 676274 579284
rect 678978 579264 679034 579320
rect 676218 578468 676274 578504
rect 676218 578448 676220 578468
rect 676220 578448 676272 578468
rect 676272 578448 676274 578468
rect 676218 577652 676274 577688
rect 676218 577632 676220 577652
rect 676220 577632 676272 577652
rect 676272 577632 676274 577652
rect 676218 577224 676274 577280
rect 676034 576952 676090 577008
rect 675942 576136 675998 576192
rect 675942 574912 675998 574968
rect 676126 575592 676182 575648
rect 676034 574504 676090 574560
rect 676034 572872 676090 572928
rect 676034 572464 676090 572520
rect 675666 572056 675722 572112
rect 678978 570696 679034 570752
rect 678978 569880 679034 569936
rect 675758 562400 675814 562456
rect 675758 561992 675814 562048
rect 675482 561176 675538 561232
rect 675390 558728 675446 558784
rect 675758 558320 675814 558376
rect 675758 557504 675814 557560
rect 676218 535880 676274 535936
rect 676034 535676 676090 535732
rect 678978 535064 679034 535120
rect 676034 534896 676036 534916
rect 676036 534896 676088 534916
rect 676088 534896 676090 534916
rect 676034 534860 676090 534896
rect 676126 534248 676182 534304
rect 676034 533264 676036 533284
rect 676036 533264 676088 533284
rect 676088 533264 676090 533284
rect 676034 533228 676090 533264
rect 675942 532820 675998 532876
rect 679070 534248 679126 534304
rect 679070 533432 679126 533488
rect 676218 532636 676274 532672
rect 676218 532616 676220 532636
rect 676220 532616 676272 532636
rect 676272 532616 676274 532636
rect 676126 531800 676182 531856
rect 676034 531188 676090 531244
rect 676034 529964 676090 530020
rect 676034 529556 676090 529612
rect 676034 527924 676090 527980
rect 676034 527516 676090 527572
rect 676034 526292 676090 526348
rect 678978 525680 679034 525736
rect 678978 524864 679034 524920
rect 676034 492088 676090 492144
rect 675942 491680 675998 491736
rect 676034 491272 676090 491328
rect 676034 490864 676090 490920
rect 675942 490456 675998 490512
rect 675850 489232 675906 489288
rect 675850 488824 675906 488880
rect 675574 488416 675630 488472
rect 675666 486376 675722 486432
rect 674010 483520 674066 483576
rect 675666 482704 675722 482760
rect 676034 490048 676090 490104
rect 676034 489640 676090 489696
rect 675942 488008 675998 488064
rect 676034 487192 676090 487248
rect 676034 485968 676090 486024
rect 676034 485560 676090 485616
rect 676034 483928 676090 483984
rect 676034 482296 676090 482352
rect 676034 481888 676090 481944
rect 676034 480700 676036 480720
rect 676036 480700 676088 480720
rect 676088 480700 676090 480720
rect 676034 480664 676090 480700
rect 675758 402192 675814 402248
rect 675666 401376 675722 401432
rect 675574 400968 675630 401024
rect 672722 148144 672778 148200
rect 672354 116048 672410 116104
rect 672262 109248 672318 109304
rect 675298 396888 675354 396944
rect 675942 403008 675998 403064
rect 675850 401784 675906 401840
rect 676218 403688 676274 403744
rect 676218 403300 676274 403336
rect 676218 403280 676220 403300
rect 676220 403280 676272 403300
rect 676272 403280 676274 403300
rect 676126 402872 676182 402928
rect 676126 400444 676182 400480
rect 676126 400424 676128 400444
rect 676128 400424 676180 400444
rect 676180 400424 676182 400444
rect 676034 400152 676090 400208
rect 676034 399744 676090 399800
rect 676034 399336 676090 399392
rect 675850 398520 675906 398576
rect 676126 398792 676182 398848
rect 676034 398112 676090 398168
rect 675942 397704 675998 397760
rect 676034 397296 676090 397352
rect 676034 396480 676090 396536
rect 675942 395664 675998 395720
rect 675942 395256 675998 395312
rect 676126 395936 676182 395992
rect 676034 394848 676090 394904
rect 676034 394440 676090 394496
rect 676126 393896 676182 393952
rect 679070 393488 679126 393544
rect 679070 392672 679126 392728
rect 672906 143112 672962 143168
rect 675850 358672 675906 358728
rect 675758 357448 675814 357504
rect 675758 357060 675814 357096
rect 675758 357040 675760 357060
rect 675760 357040 675812 357060
rect 675812 357040 675814 357060
rect 675666 356632 675722 356688
rect 675942 358264 675998 358320
rect 676034 357856 676090 357912
rect 676034 356224 676090 356280
rect 675298 355816 675354 355872
rect 676034 355428 676090 355464
rect 676034 355408 676036 355428
rect 676036 355408 676088 355428
rect 676088 355408 676090 355428
rect 674746 355000 674802 355056
rect 676034 354612 676090 354648
rect 676034 354592 676036 354612
rect 676036 354592 676088 354612
rect 676088 354592 676090 354612
rect 676034 354184 676090 354240
rect 676034 353368 676090 353424
rect 676034 352960 676090 353016
rect 675942 352552 675998 352608
rect 675298 351736 675354 351792
rect 676034 351328 676090 351384
rect 675942 350920 675998 350976
rect 676034 350104 676090 350160
rect 676034 349696 676090 349752
rect 675942 349288 675998 349344
rect 675942 348880 675998 348936
rect 676034 347268 676090 347304
rect 676034 347248 676036 347268
rect 676036 347248 676088 347268
rect 676088 347248 676090 347268
rect 675666 330520 675722 330576
rect 675758 328344 675814 328400
rect 675758 326848 675814 326904
rect 676034 313692 676036 313712
rect 676036 313692 676088 313712
rect 676088 313692 676090 313712
rect 676034 313656 676090 313692
rect 676218 313112 676274 313168
rect 676034 312876 676036 312896
rect 676036 312876 676088 312896
rect 676088 312876 676090 312896
rect 676034 312840 676090 312876
rect 676034 312468 676036 312488
rect 676036 312468 676088 312488
rect 676088 312468 676090 312488
rect 676034 312432 676090 312468
rect 676034 312060 676036 312080
rect 676036 312060 676088 312080
rect 676088 312060 676090 312080
rect 676034 312024 676090 312060
rect 676034 311652 676036 311672
rect 676036 311652 676088 311672
rect 676088 311652 676090 311672
rect 676034 311616 676090 311652
rect 676034 311208 676090 311264
rect 672998 138080 673054 138136
rect 676034 310836 676036 310856
rect 676036 310836 676088 310856
rect 676088 310836 676090 310856
rect 676034 310800 676090 310836
rect 676034 310428 676036 310448
rect 676036 310428 676088 310448
rect 676088 310428 676090 310448
rect 676034 310392 676090 310428
rect 676034 310020 676036 310040
rect 676036 310020 676088 310040
rect 676088 310020 676090 310040
rect 676034 309984 676090 310020
rect 676034 309612 676036 309632
rect 676036 309612 676088 309632
rect 676088 309612 676090 309632
rect 676034 309576 676090 309612
rect 676034 309188 676090 309224
rect 676034 309168 676036 309188
rect 676036 309168 676088 309188
rect 676088 309168 676090 309188
rect 676034 308760 676090 308816
rect 675758 308352 675814 308408
rect 675482 306720 675538 306776
rect 676034 307944 676090 308000
rect 675942 307128 675998 307184
rect 676126 307400 676182 307456
rect 676034 306312 676090 306368
rect 676126 305360 676182 305416
rect 676126 304952 676182 305008
rect 676126 304544 676182 304600
rect 675942 304272 675998 304328
rect 675850 303884 675906 303920
rect 675850 303864 675852 303884
rect 675852 303864 675904 303884
rect 675904 303864 675906 303884
rect 678978 303320 679034 303376
rect 678978 302504 679034 302560
rect 675758 291624 675814 291680
rect 676126 268504 676182 268560
rect 676034 267824 676090 267880
rect 676218 268116 676274 268152
rect 676218 268096 676220 268116
rect 676220 268096 676272 268116
rect 676272 268096 676274 268116
rect 675942 267452 675944 267472
rect 675944 267452 675996 267472
rect 675996 267452 675998 267472
rect 675942 267416 675998 267452
rect 675758 267008 675814 267064
rect 675666 265376 675722 265432
rect 675574 260480 675630 260536
rect 675574 260072 675630 260128
rect 676034 266600 676090 266656
rect 676034 266192 676090 266248
rect 676218 266092 676220 266112
rect 676220 266092 676272 266112
rect 676272 266092 676274 266112
rect 676218 266056 676274 266092
rect 676218 264832 676274 264888
rect 676034 264152 676090 264208
rect 675850 263336 675906 263392
rect 676126 263608 676182 263664
rect 676034 262928 676090 262984
rect 676126 262384 676182 262440
rect 676034 262112 676090 262168
rect 676034 261704 676090 261760
rect 675942 260888 675998 260944
rect 676126 261160 676182 261216
rect 676126 259548 676182 259584
rect 676126 259528 676128 259548
rect 676128 259528 676180 259548
rect 676180 259528 676182 259548
rect 676034 259256 676090 259312
rect 676126 258712 676182 258768
rect 678978 258304 679034 258360
rect 678978 257488 679034 257544
rect 673090 132912 673146 132968
rect 672814 127880 672870 127936
rect 674470 204992 674526 205048
rect 675666 223080 675722 223136
rect 675758 222264 675814 222320
rect 675758 221856 675814 221912
rect 675942 223488 675998 223544
rect 675850 221448 675906 221504
rect 676034 222672 676090 222728
rect 675758 221040 675814 221096
rect 675574 220632 675630 220688
rect 675390 215328 675446 215384
rect 676034 220224 676090 220280
rect 676034 219408 676090 219464
rect 676034 219000 676090 219056
rect 675942 218592 675998 218648
rect 676034 218184 676090 218240
rect 676034 217776 676090 217832
rect 675942 217368 675998 217424
rect 675942 216960 675998 217016
rect 676034 216552 676090 216608
rect 675942 216144 675998 216200
rect 675850 215736 675906 215792
rect 676034 214920 676090 214976
rect 676034 214512 676090 214568
rect 675942 214104 675998 214160
rect 676034 213696 676090 213752
rect 676034 212084 676090 212120
rect 676034 212064 676036 212084
rect 676036 212064 676088 212084
rect 676088 212064 676090 212084
rect 675574 205944 675630 206000
rect 675758 178472 675814 178528
rect 675942 178064 675998 178120
rect 675850 177248 675906 177304
rect 676034 177656 676090 177712
rect 675942 176876 675944 176896
rect 675944 176876 675996 176896
rect 675996 176876 675998 176896
rect 675942 176840 675998 176876
rect 676034 176432 676090 176488
rect 675942 176044 675998 176080
rect 675942 176024 675944 176044
rect 675944 176024 675996 176044
rect 675996 176024 675998 176044
rect 676034 175616 676090 175672
rect 675942 175244 675944 175264
rect 675944 175244 675996 175264
rect 675996 175244 675998 175264
rect 675942 175208 675998 175244
rect 676034 174800 676090 174856
rect 676034 174428 676036 174448
rect 676036 174428 676088 174448
rect 676088 174428 676090 174448
rect 676034 174392 676090 174428
rect 676034 173984 676090 174040
rect 675758 173168 675814 173224
rect 676034 172760 676090 172816
rect 675942 172352 675998 172408
rect 676034 171536 676090 171592
rect 675942 171164 675944 171184
rect 675944 171164 675996 171184
rect 675996 171164 675998 171184
rect 675942 171128 675998 171164
rect 675942 170312 675998 170368
rect 675942 169904 675998 169960
rect 676034 169496 676090 169552
rect 675942 169088 675998 169144
rect 675850 168680 675906 168736
rect 676034 168292 676090 168328
rect 676034 168272 676036 168292
rect 676036 168272 676088 168292
rect 676088 168272 676090 168292
rect 676034 167884 676090 167920
rect 676034 167864 676036 167884
rect 676036 167864 676088 167884
rect 676088 167864 676090 167884
rect 676034 167068 676090 167104
rect 676034 167048 676036 167068
rect 676036 167048 676088 167068
rect 676088 167048 676090 167068
rect 675758 156440 675814 156496
rect 675758 148416 675814 148472
rect 675758 146240 675814 146296
rect 676126 133048 676182 133104
rect 676034 132912 676090 132968
rect 676218 132640 676274 132696
rect 676218 132268 676220 132288
rect 676220 132268 676272 132288
rect 676272 132268 676274 132288
rect 676218 132232 676274 132268
rect 676034 131708 676090 131744
rect 676034 131688 676036 131708
rect 676036 131688 676088 131708
rect 676088 131688 676090 131708
rect 676218 131452 676220 131472
rect 676220 131452 676272 131472
rect 676272 131452 676274 131472
rect 676218 131416 676274 131452
rect 676034 130892 676090 130928
rect 676034 130872 676036 130892
rect 676036 130872 676088 130892
rect 676088 130872 676090 130892
rect 676218 130636 676220 130656
rect 676220 130636 676272 130656
rect 676272 130636 676274 130656
rect 676218 130600 676274 130636
rect 676034 130076 676090 130112
rect 676034 130056 676036 130076
rect 676036 130056 676088 130076
rect 676088 130056 676090 130076
rect 676034 129684 676036 129704
rect 676036 129684 676088 129704
rect 676088 129684 676090 129704
rect 676034 129648 676090 129684
rect 676218 129412 676220 129432
rect 676220 129412 676272 129432
rect 676272 129412 676274 129432
rect 676218 129376 676274 129412
rect 676034 128832 676090 128888
rect 675758 128016 675814 128072
rect 673182 122848 673238 122904
rect 672906 112648 672962 112704
rect 672446 105848 672502 105904
rect 675666 124752 675722 124808
rect 676034 127608 676090 127664
rect 675942 127200 675998 127256
rect 676034 126384 676090 126440
rect 675942 125976 675998 126032
rect 675850 125160 675906 125216
rect 675942 124344 675998 124400
rect 676126 125296 676182 125352
rect 676034 123936 676090 123992
rect 675942 123528 675998 123584
rect 676034 123140 676090 123176
rect 676034 123120 676036 123140
rect 676036 123120 676088 123140
rect 676088 123120 676090 123140
rect 676034 122732 676090 122768
rect 676034 122712 676036 122732
rect 676036 122712 676088 122732
rect 676088 122712 676090 122732
rect 676034 121916 676090 121952
rect 676034 121896 676036 121916
rect 676036 121896 676088 121916
rect 676088 121896 676090 121916
rect 675758 103264 675814 103320
rect 671986 102448 672042 102504
rect 675758 101360 675814 101416
rect 670882 100816 670938 100872
rect 666558 48456 666614 48512
rect 665178 47368 665234 47424
rect 661130 46184 661186 46240
rect 587990 41520 588046 41576
rect 530214 41248 530270 41304
rect 543002 41248 543058 41304
rect 229374 6160 229430 6216
<< metal3 >>
rect 154573 1007450 154639 1007453
rect 154573 1007448 154836 1007450
rect 154573 1007392 154578 1007448
rect 154634 1007392 154836 1007448
rect 154573 1007390 154836 1007392
rect 154573 1007387 154639 1007390
rect 501321 1007314 501387 1007317
rect 501124 1007312 501387 1007314
rect 501124 1007256 501326 1007312
rect 501382 1007256 501387 1007312
rect 501124 1007254 501387 1007256
rect 501321 1007251 501387 1007254
rect 424685 1006090 424751 1006093
rect 424580 1006088 424751 1006090
rect 424580 1006032 424690 1006088
rect 424746 1006032 424751 1006088
rect 424580 1006030 424751 1006032
rect 424685 1006027 424751 1006030
rect 423857 1005954 423923 1005957
rect 423752 1005952 423923 1005954
rect 423752 1005896 423862 1005952
rect 423918 1005896 423923 1005952
rect 423752 1005894 423923 1005896
rect 423857 1005891 423923 1005894
rect 424317 1005818 424383 1005821
rect 502977 1005818 503043 1005821
rect 503345 1005818 503411 1005821
rect 424120 1005816 424383 1005818
rect 424120 1005760 424322 1005816
rect 424378 1005760 424383 1005816
rect 424120 1005758 424383 1005760
rect 502780 1005816 503043 1005818
rect 502780 1005760 502982 1005816
rect 503038 1005760 503043 1005816
rect 502780 1005758 503043 1005760
rect 503148 1005816 503411 1005818
rect 503148 1005760 503350 1005816
rect 503406 1005760 503411 1005816
rect 503148 1005758 503411 1005760
rect 424317 1005755 424383 1005758
rect 502977 1005755 503043 1005758
rect 503345 1005755 503411 1005758
rect 356053 1005682 356119 1005685
rect 356513 1005682 356579 1005685
rect 502517 1005682 502583 1005685
rect 504541 1005682 504607 1005685
rect 355948 1005680 356119 1005682
rect 355948 1005624 356058 1005680
rect 356114 1005624 356119 1005680
rect 355948 1005622 356119 1005624
rect 356316 1005680 356579 1005682
rect 356316 1005624 356518 1005680
rect 356574 1005624 356579 1005680
rect 356316 1005622 356579 1005624
rect 502412 1005680 502583 1005682
rect 502412 1005624 502522 1005680
rect 502578 1005624 502583 1005680
rect 502412 1005622 502583 1005624
rect 504436 1005680 504607 1005682
rect 504436 1005624 504546 1005680
rect 504602 1005624 504607 1005680
rect 504436 1005622 504607 1005624
rect 356053 1005619 356119 1005622
rect 356513 1005619 356579 1005622
rect 502517 1005619 502583 1005622
rect 504541 1005619 504607 1005622
rect 160277 1005546 160343 1005549
rect 207197 1005546 207263 1005549
rect 160277 1005544 160540 1005546
rect 160277 1005488 160282 1005544
rect 160338 1005488 160540 1005544
rect 160277 1005486 160540 1005488
rect 207000 1005544 207263 1005546
rect 207000 1005488 207202 1005544
rect 207258 1005488 207263 1005544
rect 207000 1005486 207263 1005488
rect 160277 1005483 160343 1005486
rect 207197 1005483 207263 1005486
rect 209589 1005546 209655 1005549
rect 361021 1005546 361087 1005549
rect 505369 1005546 505435 1005549
rect 505829 1005546 505895 1005549
rect 209589 1005544 209852 1005546
rect 209589 1005488 209594 1005544
rect 209650 1005488 209852 1005544
rect 209589 1005486 209852 1005488
rect 360824 1005544 361087 1005546
rect 360824 1005488 361026 1005544
rect 361082 1005488 361087 1005544
rect 360824 1005486 361087 1005488
rect 505172 1005544 505435 1005546
rect 505172 1005488 505374 1005544
rect 505430 1005488 505435 1005544
rect 505172 1005486 505435 1005488
rect 505632 1005544 505895 1005546
rect 505632 1005488 505834 1005544
rect 505890 1005488 505895 1005544
rect 505632 1005486 505895 1005488
rect 209589 1005483 209655 1005486
rect 361021 1005483 361087 1005486
rect 505369 1005483 505435 1005486
rect 505829 1005483 505895 1005486
rect 263847 1005466 263913 1005469
rect 263664 1005464 263913 1005466
rect 109309 1005410 109375 1005413
rect 153745 1005410 153811 1005413
rect 154941 1005410 155007 1005413
rect 109309 1005408 109480 1005410
rect 109309 1005352 109314 1005408
rect 109370 1005352 109480 1005408
rect 109309 1005350 109480 1005352
rect 153745 1005408 153916 1005410
rect 153745 1005352 153750 1005408
rect 153806 1005352 153916 1005408
rect 153745 1005350 153916 1005352
rect 154941 1005408 155204 1005410
rect 154941 1005352 154946 1005408
rect 155002 1005352 155204 1005408
rect 263664 1005408 263852 1005464
rect 263908 1005408 263913 1005464
rect 360193 1005410 360259 1005413
rect 423489 1005410 423555 1005413
rect 263664 1005406 263913 1005408
rect 263847 1005403 263913 1005406
rect 359996 1005408 360259 1005410
rect 154941 1005350 155204 1005352
rect 359996 1005352 360198 1005408
rect 360254 1005352 360259 1005408
rect 359996 1005350 360259 1005352
rect 423292 1005408 423555 1005410
rect 423292 1005352 423494 1005408
rect 423550 1005352 423555 1005408
rect 423292 1005350 423555 1005352
rect 109309 1005347 109375 1005350
rect 153745 1005347 153811 1005350
rect 154941 1005347 155007 1005350
rect 360193 1005347 360259 1005350
rect 423489 1005347 423555 1005350
rect 151261 1005274 151327 1005277
rect 153285 1005274 153351 1005277
rect 259821 1005274 259887 1005277
rect 260189 1005274 260255 1005277
rect 359733 1005274 359799 1005277
rect 428365 1005274 428431 1005277
rect 151261 1005272 151524 1005274
rect 151261 1005216 151266 1005272
rect 151322 1005216 151524 1005272
rect 151261 1005214 151524 1005216
rect 153285 1005272 153548 1005274
rect 153285 1005216 153290 1005272
rect 153346 1005216 153548 1005272
rect 153285 1005214 153548 1005216
rect 259624 1005272 259887 1005274
rect 259624 1005216 259826 1005272
rect 259882 1005216 259887 1005272
rect 259624 1005214 259887 1005216
rect 260084 1005272 260255 1005274
rect 260084 1005216 260194 1005272
rect 260250 1005216 260255 1005272
rect 260084 1005214 260255 1005216
rect 359628 1005272 359799 1005274
rect 359628 1005216 359738 1005272
rect 359794 1005216 359799 1005272
rect 359628 1005214 359799 1005216
rect 428260 1005272 428431 1005274
rect 428260 1005216 428370 1005272
rect 428426 1005216 428431 1005272
rect 428260 1005214 428431 1005216
rect 151261 1005211 151327 1005214
rect 153285 1005211 153351 1005214
rect 259821 1005211 259887 1005214
rect 260189 1005211 260255 1005214
rect 359733 1005211 359799 1005214
rect 428365 1005211 428431 1005214
rect 106457 1005138 106523 1005141
rect 106260 1005136 106523 1005138
rect 106260 1005080 106462 1005136
rect 106518 1005080 106523 1005136
rect 106260 1005078 106523 1005080
rect 106457 1005075 106523 1005078
rect 143809 1005138 143875 1005141
rect 148869 1005138 148935 1005141
rect 149697 1005138 149763 1005141
rect 143809 1005136 148935 1005138
rect 143809 1005080 143814 1005136
rect 143870 1005080 148874 1005136
rect 148930 1005080 148935 1005136
rect 143809 1005078 148935 1005080
rect 149500 1005136 149763 1005138
rect 149500 1005080 149702 1005136
rect 149758 1005080 149763 1005136
rect 149500 1005078 149763 1005080
rect 143809 1005075 143875 1005078
rect 148869 1005075 148935 1005078
rect 149697 1005075 149763 1005078
rect 150433 1005138 150499 1005141
rect 208393 1005138 208459 1005141
rect 261845 1005138 261911 1005141
rect 263041 1005138 263107 1005141
rect 150433 1005136 150696 1005138
rect 150433 1005080 150438 1005136
rect 150494 1005080 150696 1005136
rect 150433 1005078 150696 1005080
rect 208196 1005136 208459 1005138
rect 208196 1005080 208398 1005136
rect 208454 1005080 208459 1005136
rect 208196 1005078 208459 1005080
rect 261648 1005136 261911 1005138
rect 261648 1005080 261850 1005136
rect 261906 1005080 261911 1005136
rect 261648 1005078 261911 1005080
rect 262844 1005136 263107 1005138
rect 262844 1005080 263046 1005136
rect 263102 1005080 263107 1005136
rect 262844 1005078 263107 1005080
rect 150433 1005075 150499 1005078
rect 208393 1005075 208459 1005078
rect 261845 1005075 261911 1005078
rect 263041 1005075 263107 1005078
rect 265529 1005138 265595 1005141
rect 267005 1005138 267071 1005141
rect 358169 1005138 358235 1005141
rect 428825 1005138 428891 1005141
rect 504173 1005138 504239 1005141
rect 551921 1005138 551987 1005141
rect 265529 1005136 267071 1005138
rect 265529 1005080 265534 1005136
rect 265590 1005080 267010 1005136
rect 267066 1005080 267071 1005136
rect 265529 1005078 267071 1005080
rect 357972 1005136 358235 1005138
rect 357972 1005080 358174 1005136
rect 358230 1005080 358235 1005136
rect 357972 1005078 358235 1005080
rect 428628 1005136 428891 1005138
rect 428628 1005080 428830 1005136
rect 428886 1005080 428891 1005136
rect 428628 1005078 428891 1005080
rect 503976 1005136 504239 1005138
rect 503976 1005080 504178 1005136
rect 504234 1005080 504239 1005136
rect 503976 1005078 504239 1005080
rect 551724 1005136 551987 1005138
rect 551724 1005080 551926 1005136
rect 551982 1005080 551987 1005136
rect 551724 1005078 551987 1005080
rect 265529 1005075 265595 1005078
rect 267005 1005075 267071 1005078
rect 358169 1005075 358235 1005078
rect 428825 1005075 428891 1005078
rect 504173 1005075 504239 1005078
rect 551921 1005075 551987 1005078
rect 143717 1005002 143783 1005005
rect 148869 1005002 148935 1005005
rect 143717 1005000 148935 1005002
rect 143717 1004944 143722 1005000
rect 143778 1004944 148874 1005000
rect 148930 1004944 148935 1005000
rect 143717 1004942 148935 1004944
rect 143717 1004939 143783 1004942
rect 148869 1004939 148935 1004942
rect 150893 1005002 150959 1005005
rect 154113 1005002 154179 1005005
rect 159449 1005002 159515 1005005
rect 209221 1005002 209287 1005005
rect 150893 1005000 151156 1005002
rect 150893 1004944 150898 1005000
rect 150954 1004944 151156 1005000
rect 150893 1004942 151156 1004944
rect 154113 1005000 154376 1005002
rect 154113 1004944 154118 1005000
rect 154174 1004944 154376 1005000
rect 154113 1004942 154376 1004944
rect 159252 1005000 159515 1005002
rect 159252 1004944 159454 1005000
rect 159510 1004944 159515 1005000
rect 159252 1004942 159515 1004944
rect 209024 1005000 209287 1005002
rect 209024 1004944 209226 1005000
rect 209282 1004944 209287 1005000
rect 209024 1004942 209287 1004944
rect 150893 1004939 150959 1004942
rect 154113 1004939 154179 1004942
rect 159449 1004939 159515 1004942
rect 209221 1004939 209287 1004942
rect 211613 1005002 211679 1005005
rect 260649 1005002 260715 1005005
rect 262673 1005002 262739 1005005
rect 211613 1005000 211876 1005002
rect 211613 1004944 211618 1005000
rect 211674 1004944 211876 1005000
rect 211613 1004942 211876 1004944
rect 260452 1005000 260715 1005002
rect 260452 1004944 260654 1005000
rect 260710 1004944 260715 1005000
rect 260452 1004942 260715 1004944
rect 262476 1005000 262739 1005002
rect 262476 1004944 262678 1005000
rect 262734 1004944 262739 1005000
rect 262476 1004942 262739 1004944
rect 211613 1004939 211679 1004942
rect 260649 1004939 260715 1004942
rect 262673 1004939 262739 1004942
rect 265529 1005002 265595 1005005
rect 266625 1005002 266691 1005005
rect 356881 1005002 356947 1005005
rect 358537 1005002 358603 1005005
rect 425513 1005002 425579 1005005
rect 426801 1005002 426867 1005005
rect 505001 1005002 505067 1005005
rect 265529 1005000 266691 1005002
rect 265529 1004944 265534 1005000
rect 265590 1004944 266630 1005000
rect 266686 1004944 266691 1005000
rect 265529 1004942 266691 1004944
rect 356684 1005000 356947 1005002
rect 356684 1004944 356886 1005000
rect 356942 1004944 356947 1005000
rect 356684 1004942 356947 1004944
rect 358340 1005000 358603 1005002
rect 358340 1004944 358542 1005000
rect 358598 1004944 358603 1005000
rect 358340 1004942 358603 1004944
rect 425316 1005000 425579 1005002
rect 425316 1004944 425518 1005000
rect 425574 1004944 425579 1005000
rect 425316 1004942 425579 1004944
rect 426604 1005000 426867 1005002
rect 426604 1004944 426806 1005000
rect 426862 1004944 426867 1005000
rect 426604 1004942 426867 1004944
rect 504804 1005000 505067 1005002
rect 504804 1004944 505006 1005000
rect 505062 1004944 505067 1005000
rect 504804 1004942 505067 1004944
rect 265529 1004939 265595 1004942
rect 266625 1004939 266691 1004942
rect 356881 1004939 356947 1004942
rect 358537 1004939 358603 1004942
rect 425513 1004939 425579 1004942
rect 426801 1004939 426867 1004942
rect 505001 1004939 505067 1004942
rect 554773 1005002 554839 1005005
rect 554773 1005000 555036 1005002
rect 554773 1004944 554778 1005000
rect 554834 1004944 555036 1005000
rect 554773 1004942 555036 1004944
rect 554773 1004939 554839 1004942
rect 108021 1004866 108087 1004869
rect 107916 1004864 108087 1004866
rect 107916 1004808 108026 1004864
rect 108082 1004808 108087 1004864
rect 107916 1004806 108087 1004808
rect 108021 1004803 108087 1004806
rect 108849 1004866 108915 1004869
rect 147581 1004866 147647 1004869
rect 148869 1004866 148935 1004869
rect 108849 1004864 109112 1004866
rect 108849 1004808 108854 1004864
rect 108910 1004808 109112 1004864
rect 108849 1004806 109112 1004808
rect 147581 1004864 148935 1004866
rect 147581 1004808 147586 1004864
rect 147642 1004808 148874 1004864
rect 148930 1004808 148935 1004864
rect 147581 1004806 148935 1004808
rect 108849 1004803 108915 1004806
rect 147581 1004803 147647 1004806
rect 148869 1004803 148935 1004806
rect 152089 1004866 152155 1004869
rect 152917 1004866 152983 1004869
rect 156965 1004866 157031 1004869
rect 152089 1004864 152352 1004866
rect 152089 1004808 152094 1004864
rect 152150 1004808 152352 1004864
rect 152089 1004806 152352 1004808
rect 152917 1004864 153180 1004866
rect 152917 1004808 152922 1004864
rect 152978 1004808 153180 1004864
rect 152917 1004806 153180 1004808
rect 156860 1004864 157031 1004866
rect 156860 1004808 156970 1004864
rect 157026 1004808 157031 1004864
rect 156860 1004806 157031 1004808
rect 152089 1004803 152155 1004806
rect 152917 1004803 152983 1004806
rect 156965 1004803 157031 1004806
rect 206369 1004866 206435 1004869
rect 210877 1004866 210943 1004869
rect 261017 1004866 261083 1004869
rect 262213 1004866 262279 1004869
rect 357341 1004866 357407 1004869
rect 357709 1004866 357775 1004869
rect 427169 1004866 427235 1004869
rect 427537 1004866 427603 1004869
rect 500493 1004866 500559 1004869
rect 553117 1004866 553183 1004869
rect 553945 1004866 554011 1004869
rect 567469 1004866 567535 1004869
rect 206369 1004864 206540 1004866
rect 206369 1004808 206374 1004864
rect 206430 1004808 206540 1004864
rect 206369 1004806 206540 1004808
rect 210680 1004864 210943 1004866
rect 210680 1004808 210882 1004864
rect 210938 1004808 210943 1004864
rect 210680 1004806 210943 1004808
rect 260820 1004864 261083 1004866
rect 260820 1004808 261022 1004864
rect 261078 1004808 261083 1004864
rect 260820 1004806 261083 1004808
rect 262108 1004864 262279 1004866
rect 262108 1004808 262218 1004864
rect 262274 1004808 262279 1004864
rect 262108 1004806 262279 1004808
rect 357144 1004864 357407 1004866
rect 357144 1004808 357346 1004864
rect 357402 1004808 357407 1004864
rect 357144 1004806 357407 1004808
rect 357604 1004864 357775 1004866
rect 357604 1004808 357714 1004864
rect 357770 1004808 357775 1004864
rect 357604 1004806 357775 1004808
rect 426972 1004864 427235 1004866
rect 426972 1004808 427174 1004864
rect 427230 1004808 427235 1004864
rect 426972 1004806 427235 1004808
rect 427340 1004864 427603 1004866
rect 427340 1004808 427542 1004864
rect 427598 1004808 427603 1004864
rect 427340 1004806 427603 1004808
rect 500296 1004864 500559 1004866
rect 500296 1004808 500498 1004864
rect 500554 1004808 500559 1004864
rect 500296 1004806 500559 1004808
rect 552920 1004864 553183 1004866
rect 552920 1004808 553122 1004864
rect 553178 1004808 553183 1004864
rect 552920 1004806 553183 1004808
rect 553748 1004864 554011 1004866
rect 553748 1004808 553950 1004864
rect 554006 1004808 554011 1004864
rect 553748 1004806 554011 1004808
rect 561476 1004864 567535 1004866
rect 561476 1004808 567474 1004864
rect 567530 1004808 567535 1004864
rect 561476 1004806 567535 1004808
rect 206369 1004803 206435 1004806
rect 210877 1004803 210943 1004806
rect 261017 1004803 261083 1004806
rect 262213 1004803 262279 1004806
rect 357341 1004803 357407 1004806
rect 357709 1004803 357775 1004806
rect 427169 1004803 427235 1004806
rect 427537 1004803 427603 1004806
rect 500493 1004803 500559 1004806
rect 553117 1004803 553183 1004806
rect 553945 1004803 554011 1004806
rect 567469 1004803 567535 1004806
rect 98269 1004730 98335 1004733
rect 99097 1004730 99163 1004733
rect 105629 1004730 105695 1004733
rect 98072 1004728 98335 1004730
rect 98072 1004672 98274 1004728
rect 98330 1004672 98335 1004728
rect 98072 1004670 98335 1004672
rect 98532 1004670 98900 1004730
rect 99097 1004728 99268 1004730
rect 99097 1004672 99102 1004728
rect 99158 1004672 99268 1004728
rect 99097 1004670 99268 1004672
rect 105432 1004728 105695 1004730
rect 105432 1004672 105634 1004728
rect 105690 1004672 105695 1004728
rect 105432 1004670 105695 1004672
rect 98269 1004667 98335 1004670
rect 99097 1004667 99163 1004670
rect 105629 1004667 105695 1004670
rect 147765 1004730 147831 1004733
rect 148869 1004730 148935 1004733
rect 151721 1004730 151787 1004733
rect 152549 1004730 152615 1004733
rect 157793 1004730 157859 1004733
rect 147765 1004728 148935 1004730
rect 147765 1004672 147770 1004728
rect 147826 1004672 148874 1004728
rect 148930 1004672 148935 1004728
rect 147765 1004670 148935 1004672
rect 149868 1004670 150328 1004730
rect 151721 1004728 151892 1004730
rect 151721 1004672 151726 1004728
rect 151782 1004672 151892 1004728
rect 151721 1004670 151892 1004672
rect 152549 1004728 152720 1004730
rect 152549 1004672 152554 1004728
rect 152610 1004672 152720 1004728
rect 152549 1004670 152720 1004672
rect 157596 1004728 157859 1004730
rect 157596 1004672 157798 1004728
rect 157854 1004672 157859 1004728
rect 157596 1004670 157859 1004672
rect 147765 1004667 147831 1004670
rect 148869 1004667 148935 1004670
rect 151721 1004667 151787 1004670
rect 152549 1004667 152615 1004670
rect 157793 1004667 157859 1004670
rect 160645 1004730 160711 1004733
rect 201033 1004730 201099 1004733
rect 201861 1004730 201927 1004733
rect 205909 1004730 205975 1004733
rect 212453 1004730 212519 1004733
rect 252461 1004730 252527 1004733
rect 253289 1004730 253355 1004733
rect 261477 1004730 261543 1004733
rect 263501 1004730 263567 1004733
rect 160645 1004728 160908 1004730
rect 160645 1004672 160650 1004728
rect 160706 1004672 160908 1004728
rect 160645 1004670 160908 1004672
rect 200836 1004728 201099 1004730
rect 200836 1004672 201038 1004728
rect 201094 1004672 201099 1004728
rect 200836 1004670 201099 1004672
rect 201296 1004670 201756 1004730
rect 201861 1004728 202124 1004730
rect 201861 1004672 201866 1004728
rect 201922 1004672 202124 1004728
rect 201861 1004670 202124 1004672
rect 205909 1004728 206172 1004730
rect 205909 1004672 205914 1004728
rect 205970 1004672 206172 1004728
rect 205909 1004670 206172 1004672
rect 212336 1004728 212519 1004730
rect 212336 1004672 212458 1004728
rect 212514 1004672 212519 1004728
rect 212336 1004670 212519 1004672
rect 252264 1004728 252527 1004730
rect 252264 1004672 252466 1004728
rect 252522 1004672 252527 1004728
rect 252264 1004670 252527 1004672
rect 252724 1004670 253092 1004730
rect 253289 1004728 253460 1004730
rect 253289 1004672 253294 1004728
rect 253350 1004672 253460 1004728
rect 253289 1004670 253460 1004672
rect 261280 1004728 261543 1004730
rect 261280 1004672 261482 1004728
rect 261538 1004672 261543 1004728
rect 261280 1004670 261543 1004672
rect 263304 1004728 263567 1004730
rect 263304 1004672 263506 1004728
rect 263562 1004672 263567 1004728
rect 263304 1004670 263567 1004672
rect 160645 1004667 160711 1004670
rect 201033 1004667 201099 1004670
rect 201861 1004667 201927 1004670
rect 205909 1004667 205975 1004670
rect 212453 1004667 212519 1004670
rect 252461 1004667 252527 1004670
rect 253289 1004667 253355 1004670
rect 261477 1004667 261543 1004670
rect 263501 1004667 263567 1004670
rect 265469 1004730 265535 1004733
rect 266533 1004730 266599 1004733
rect 315113 1004730 315179 1004733
rect 265469 1004728 266599 1004730
rect 265469 1004672 265474 1004728
rect 265530 1004672 266538 1004728
rect 266594 1004672 266599 1004728
rect 265469 1004670 266599 1004672
rect 304244 1004670 304704 1004730
rect 314916 1004728 315179 1004730
rect 314916 1004672 315118 1004728
rect 315174 1004672 315179 1004728
rect 314916 1004670 315179 1004672
rect 265469 1004667 265535 1004670
rect 266533 1004667 266599 1004670
rect 315113 1004667 315179 1004670
rect 350441 1004730 350507 1004733
rect 353661 1004730 353727 1004733
rect 350441 1004728 353727 1004730
rect 350441 1004672 350446 1004728
rect 350502 1004672 353666 1004728
rect 353722 1004672 353727 1004728
rect 350441 1004670 353727 1004672
rect 350441 1004667 350507 1004670
rect 353661 1004667 353727 1004670
rect 354029 1004730 354095 1004733
rect 354489 1004730 354555 1004733
rect 355225 1004730 355291 1004733
rect 360561 1004730 360627 1004733
rect 361389 1004730 361455 1004733
rect 371325 1004730 371391 1004733
rect 421833 1004730 421899 1004733
rect 422661 1004730 422727 1004733
rect 425145 1004730 425211 1004733
rect 498837 1004730 498903 1004733
rect 499665 1004730 499731 1004733
rect 501689 1004730 501755 1004733
rect 502149 1004730 502215 1004733
rect 354029 1004728 354555 1004730
rect 354029 1004672 354034 1004728
rect 354090 1004672 354494 1004728
rect 354550 1004672 354555 1004728
rect 354029 1004670 354555 1004672
rect 354660 1004670 355120 1004730
rect 355225 1004728 355488 1004730
rect 355225 1004672 355230 1004728
rect 355286 1004672 355488 1004728
rect 355225 1004670 355488 1004672
rect 360364 1004728 360627 1004730
rect 360364 1004672 360566 1004728
rect 360622 1004672 360627 1004728
rect 360364 1004670 360627 1004672
rect 361192 1004728 361455 1004730
rect 361192 1004672 361394 1004728
rect 361450 1004672 361455 1004728
rect 361192 1004670 361455 1004672
rect 365700 1004728 371391 1004730
rect 365700 1004672 371330 1004728
rect 371386 1004672 371391 1004728
rect 365700 1004670 371391 1004672
rect 421636 1004728 421899 1004730
rect 421636 1004672 421838 1004728
rect 421894 1004672 421899 1004728
rect 421636 1004670 421899 1004672
rect 422096 1004670 422556 1004730
rect 422661 1004728 422924 1004730
rect 422661 1004672 422666 1004728
rect 422722 1004672 422924 1004728
rect 422661 1004670 422924 1004672
rect 424948 1004728 425211 1004730
rect 424948 1004672 425150 1004728
rect 425206 1004672 425211 1004728
rect 424948 1004670 425211 1004672
rect 498732 1004728 498903 1004730
rect 498732 1004672 498842 1004728
rect 498898 1004672 498903 1004728
rect 498732 1004670 498903 1004672
rect 499100 1004670 499468 1004730
rect 499665 1004728 499928 1004730
rect 499665 1004672 499670 1004728
rect 499726 1004672 499928 1004728
rect 499665 1004670 499928 1004672
rect 501492 1004728 501755 1004730
rect 501492 1004672 501694 1004728
rect 501750 1004672 501755 1004728
rect 501492 1004670 501755 1004672
rect 501952 1004728 502215 1004730
rect 501952 1004672 502154 1004728
rect 502210 1004672 502215 1004728
rect 501952 1004670 502215 1004672
rect 354029 1004667 354095 1004670
rect 354489 1004667 354555 1004670
rect 355225 1004667 355291 1004670
rect 360561 1004667 360627 1004670
rect 361389 1004667 361455 1004670
rect 371325 1004667 371391 1004670
rect 421833 1004667 421899 1004670
rect 422661 1004667 422727 1004670
rect 425145 1004667 425211 1004670
rect 498837 1004667 498903 1004670
rect 499665 1004667 499731 1004670
rect 501689 1004667 501755 1004670
rect 502149 1004667 502215 1004670
rect 546401 1004730 546467 1004733
rect 549437 1004730 549503 1004733
rect 550265 1004730 550331 1004733
rect 551093 1004730 551159 1004733
rect 552749 1004730 552815 1004733
rect 546401 1004728 549503 1004730
rect 546401 1004672 546406 1004728
rect 546462 1004672 549442 1004728
rect 549498 1004672 549503 1004728
rect 546401 1004670 549503 1004672
rect 550068 1004728 550331 1004730
rect 550068 1004672 550270 1004728
rect 550326 1004672 550331 1004728
rect 550068 1004670 550331 1004672
rect 550436 1004670 550896 1004730
rect 551093 1004728 551356 1004730
rect 551093 1004672 551098 1004728
rect 551154 1004672 551356 1004728
rect 551093 1004670 551356 1004672
rect 552552 1004728 552815 1004730
rect 552552 1004672 552754 1004728
rect 552810 1004672 552815 1004728
rect 552552 1004670 552815 1004672
rect 546401 1004667 546467 1004670
rect 549437 1004667 549503 1004670
rect 550265 1004667 550331 1004670
rect 551093 1004667 551159 1004670
rect 552749 1004667 552815 1004670
rect 555141 1004730 555207 1004733
rect 555141 1004728 555404 1004730
rect 555141 1004672 555146 1004728
rect 555202 1004672 555404 1004728
rect 555141 1004670 555404 1004672
rect 555141 1004667 555207 1004670
rect 553485 1003506 553551 1003509
rect 553380 1003504 553551 1003506
rect 553380 1003448 553490 1003504
rect 553546 1003448 553551 1003504
rect 553380 1003446 553551 1003448
rect 553485 1003443 553551 1003446
rect 554313 1003234 554379 1003237
rect 554116 1003232 554379 1003234
rect 554116 1003176 554318 1003232
rect 554374 1003176 554379 1003232
rect 554116 1003174 554379 1003176
rect 554313 1003171 554379 1003174
rect 426341 1000650 426407 1000653
rect 427997 1000650 428063 1000653
rect 426144 1000648 426407 1000650
rect 426144 1000592 426346 1000648
rect 426402 1000592 426407 1000648
rect 426144 1000590 426407 1000592
rect 427800 1000648 428063 1000650
rect 427800 1000592 428002 1000648
rect 428058 1000592 428063 1000648
rect 427800 1000590 428063 1000592
rect 426341 1000587 426407 1000590
rect 427997 1000587 428063 1000590
rect 358905 1000514 358971 1000517
rect 425973 1000514 426039 1000517
rect 358800 1000512 358971 1000514
rect 358800 1000456 358910 1000512
rect 358966 1000456 358971 1000512
rect 358800 1000454 358971 1000456
rect 425776 1000512 426039 1000514
rect 425776 1000456 425978 1000512
rect 426034 1000456 426039 1000512
rect 425776 1000454 426039 1000456
rect 358905 1000451 358971 1000454
rect 425973 1000451 426039 1000454
rect 555969 1000106 556035 1000109
rect 555772 1000104 556035 1000106
rect 555772 1000048 555974 1000104
rect 556030 1000048 556035 1000104
rect 555772 1000046 556035 1000048
rect 555969 1000043 556035 1000046
rect 258625 999970 258691 999973
rect 558453 999970 558519 999973
rect 258625 999968 258796 999970
rect 258625 999912 258630 999968
rect 258686 999912 258796 999968
rect 258625 999910 258796 999912
rect 558256 999968 558519 999970
rect 558256 999912 558458 999968
rect 558514 999912 558519 999968
rect 558256 999910 558519 999912
rect 258625 999907 258691 999910
rect 558453 999907 558519 999910
rect 102777 999834 102843 999837
rect 104341 999834 104407 999837
rect 256969 999834 257035 999837
rect 257337 999834 257403 999837
rect 310145 999834 310211 999837
rect 312169 999834 312235 999837
rect 430849 999834 430915 999837
rect 431677 999834 431743 999837
rect 508681 999834 508747 999837
rect 556337 999834 556403 999837
rect 560845 999834 560911 999837
rect 102777 999832 102948 999834
rect 102777 999776 102782 999832
rect 102838 999776 102948 999832
rect 102777 999774 102948 999776
rect 104341 999832 104604 999834
rect 104341 999776 104346 999832
rect 104402 999776 104604 999832
rect 104341 999774 104604 999776
rect 256969 999832 257140 999834
rect 256969 999776 256974 999832
rect 257030 999776 257140 999832
rect 256969 999774 257140 999776
rect 257337 999832 257600 999834
rect 257337 999776 257342 999832
rect 257398 999776 257600 999832
rect 257337 999774 257600 999776
rect 309948 999832 310211 999834
rect 309948 999776 310150 999832
rect 310206 999776 310211 999832
rect 309948 999774 310211 999776
rect 312064 999832 312235 999834
rect 312064 999776 312174 999832
rect 312230 999776 312235 999832
rect 312064 999774 312235 999776
rect 430652 999832 430915 999834
rect 430652 999776 430854 999832
rect 430910 999776 430915 999832
rect 430652 999774 430915 999776
rect 431480 999832 431743 999834
rect 431480 999776 431682 999832
rect 431738 999776 431743 999832
rect 431480 999774 431743 999776
rect 508484 999832 508747 999834
rect 508484 999776 508686 999832
rect 508742 999776 508747 999832
rect 508484 999774 508747 999776
rect 556232 999832 556403 999834
rect 556232 999776 556342 999832
rect 556398 999776 556403 999832
rect 556232 999774 556403 999776
rect 560740 999832 560911 999834
rect 560740 999776 560850 999832
rect 560906 999776 560911 999832
rect 560740 999774 560911 999776
rect 102777 999771 102843 999774
rect 104341 999771 104407 999774
rect 256969 999771 257035 999774
rect 257337 999771 257403 999774
rect 310145 999771 310211 999774
rect 312169 999771 312235 999774
rect 430849 999771 430915 999774
rect 431677 999771 431743 999774
rect 508681 999771 508747 999774
rect 556337 999771 556403 999774
rect 560845 999771 560911 999774
rect 100661 999698 100727 999701
rect 102317 999698 102383 999701
rect 203885 999698 203951 999701
rect 205541 999698 205607 999701
rect 254853 999698 254919 999701
rect 257797 999698 257863 999701
rect 311433 999698 311499 999701
rect 313825 999698 313891 999701
rect 361849 999698 361915 999701
rect 362585 999698 362651 999701
rect 429193 999698 429259 999701
rect 430021 999698 430087 999701
rect 506197 999698 506263 999701
rect 508221 999698 508287 999701
rect 559189 999698 559255 999701
rect 560477 999698 560543 999701
rect 100661 999696 100924 999698
rect 100661 999640 100666 999696
rect 100722 999640 100924 999696
rect 100661 999638 100924 999640
rect 102317 999696 102580 999698
rect 102317 999640 102322 999696
rect 102378 999640 102580 999696
rect 102317 999638 102580 999640
rect 203885 999696 204148 999698
rect 203885 999640 203890 999696
rect 203946 999640 204148 999696
rect 203885 999638 204148 999640
rect 205541 999696 205804 999698
rect 205541 999640 205546 999696
rect 205602 999640 205804 999696
rect 205541 999638 205804 999640
rect 254853 999696 255116 999698
rect 254853 999640 254858 999696
rect 254914 999640 255116 999696
rect 254853 999638 255116 999640
rect 257797 999696 257968 999698
rect 257797 999640 257802 999696
rect 257858 999640 257968 999696
rect 257797 999638 257968 999640
rect 311236 999696 311499 999698
rect 311236 999640 311438 999696
rect 311494 999640 311499 999696
rect 311236 999638 311499 999640
rect 313628 999696 313891 999698
rect 313628 999640 313830 999696
rect 313886 999640 313891 999696
rect 313628 999638 313891 999640
rect 361652 999696 361915 999698
rect 361652 999640 361854 999696
rect 361910 999640 361915 999696
rect 361652 999638 361915 999640
rect 362388 999696 362651 999698
rect 362388 999640 362590 999696
rect 362646 999640 362651 999696
rect 362388 999638 362651 999640
rect 428996 999696 429259 999698
rect 428996 999640 429198 999696
rect 429254 999640 429259 999696
rect 428996 999638 429259 999640
rect 429824 999696 430087 999698
rect 429824 999640 430026 999696
rect 430082 999640 430087 999696
rect 429824 999638 430087 999640
rect 506000 999696 506263 999698
rect 506000 999640 506202 999696
rect 506258 999640 506263 999696
rect 506000 999638 506263 999640
rect 508116 999696 508287 999698
rect 508116 999640 508226 999696
rect 508282 999640 508287 999696
rect 508116 999638 508287 999640
rect 559084 999696 559255 999698
rect 559084 999640 559194 999696
rect 559250 999640 559255 999696
rect 559084 999638 559255 999640
rect 560280 999696 560543 999698
rect 560280 999640 560482 999696
rect 560538 999640 560543 999696
rect 560280 999638 560543 999640
rect 100661 999635 100727 999638
rect 102317 999635 102383 999638
rect 203885 999635 203951 999638
rect 205541 999635 205607 999638
rect 254853 999635 254919 999638
rect 257797 999635 257863 999638
rect 311433 999635 311499 999638
rect 313825 999635 313891 999638
rect 361849 999635 361915 999638
rect 362585 999635 362651 999638
rect 429193 999635 429259 999638
rect 430021 999635 430087 999638
rect 506197 999635 506263 999638
rect 508221 999635 508287 999638
rect 559189 999635 559255 999638
rect 560477 999635 560543 999638
rect 101489 999562 101555 999565
rect 101949 999562 102015 999565
rect 155769 999562 155835 999565
rect 159081 999562 159147 999565
rect 101489 999560 101752 999562
rect 101489 999504 101494 999560
rect 101550 999504 101752 999560
rect 101489 999502 101752 999504
rect 101949 999560 102212 999562
rect 101949 999504 101954 999560
rect 102010 999504 102212 999560
rect 101949 999502 102212 999504
rect 155572 999560 155835 999562
rect 155572 999504 155774 999560
rect 155830 999504 155835 999560
rect 155572 999502 155835 999504
rect 158884 999560 159147 999562
rect 158884 999504 159086 999560
rect 159142 999504 159147 999560
rect 158884 999502 159147 999504
rect 101489 999499 101555 999502
rect 101949 999499 102015 999502
rect 155769 999499 155835 999502
rect 159081 999499 159147 999502
rect 203517 999562 203583 999565
rect 204345 999562 204411 999565
rect 255681 999562 255747 999565
rect 256141 999562 256207 999565
rect 312629 999562 312695 999565
rect 203517 999560 203780 999562
rect 203517 999504 203522 999560
rect 203578 999504 203780 999560
rect 203517 999502 203780 999504
rect 204345 999560 204516 999562
rect 204345 999504 204350 999560
rect 204406 999504 204516 999560
rect 204345 999502 204516 999504
rect 255681 999560 255944 999562
rect 255681 999504 255686 999560
rect 255742 999504 255944 999560
rect 255681 999502 255944 999504
rect 256141 999560 256404 999562
rect 256141 999504 256146 999560
rect 256202 999504 256404 999560
rect 256141 999502 256404 999504
rect 312432 999560 312695 999562
rect 312432 999504 312634 999560
rect 312690 999504 312695 999560
rect 312432 999502 312695 999504
rect 203517 999499 203583 999502
rect 204345 999499 204411 999502
rect 255681 999499 255747 999502
rect 256141 999499 256207 999502
rect 312629 999499 312695 999502
rect 314653 999562 314719 999565
rect 363413 999562 363479 999565
rect 365069 999562 365135 999565
rect 431217 999562 431283 999565
rect 432413 999562 432479 999565
rect 507025 999562 507091 999565
rect 507853 999562 507919 999565
rect 557993 999562 558059 999565
rect 560017 999562 560083 999565
rect 314653 999560 314762 999562
rect 314653 999504 314658 999560
rect 314714 999504 314762 999560
rect 314653 999499 314762 999504
rect 363308 999560 363479 999562
rect 363308 999504 363418 999560
rect 363474 999504 363479 999560
rect 363308 999502 363479 999504
rect 364872 999560 365135 999562
rect 364872 999504 365074 999560
rect 365130 999504 365135 999560
rect 364872 999502 365135 999504
rect 431020 999560 431283 999562
rect 431020 999504 431222 999560
rect 431278 999504 431283 999560
rect 431020 999502 431283 999504
rect 432308 999560 432479 999562
rect 432308 999504 432418 999560
rect 432474 999504 432479 999560
rect 432308 999502 432479 999504
rect 506828 999560 507091 999562
rect 506828 999504 507030 999560
rect 507086 999504 507091 999560
rect 506828 999502 507091 999504
rect 507656 999560 507919 999562
rect 507656 999504 507858 999560
rect 507914 999504 507919 999560
rect 507656 999502 507919 999504
rect 557796 999560 558059 999562
rect 557796 999504 557998 999560
rect 558054 999504 558059 999560
rect 557796 999502 558059 999504
rect 559820 999560 560083 999562
rect 559820 999504 560022 999560
rect 560078 999504 560083 999560
rect 559820 999502 560083 999504
rect 363413 999499 363479 999502
rect 365069 999499 365135 999502
rect 431217 999499 431283 999502
rect 432413 999499 432479 999502
rect 507025 999499 507091 999502
rect 507853 999499 507919 999502
rect 557993 999499 558059 999502
rect 560017 999499 560083 999502
rect 99465 999426 99531 999429
rect 103145 999426 103211 999429
rect 202229 999426 202295 999429
rect 204713 999426 204779 999429
rect 208853 999426 208919 999429
rect 210417 999426 210483 999429
rect 99465 999424 99728 999426
rect 99465 999368 99470 999424
rect 99526 999368 99728 999424
rect 99465 999366 99728 999368
rect 103145 999424 103408 999426
rect 103145 999368 103150 999424
rect 103206 999368 103408 999424
rect 103145 999366 103408 999368
rect 202229 999424 202492 999426
rect 202229 999368 202234 999424
rect 202290 999368 202492 999424
rect 202229 999366 202492 999368
rect 204713 999424 204976 999426
rect 204713 999368 204718 999424
rect 204774 999368 204976 999424
rect 204713 999366 204976 999368
rect 208656 999424 208919 999426
rect 208656 999368 208858 999424
rect 208914 999368 208919 999424
rect 208656 999366 208919 999368
rect 210220 999424 210483 999426
rect 210220 999368 210422 999424
rect 210478 999368 210483 999424
rect 210220 999366 210483 999368
rect 99465 999363 99531 999366
rect 103145 999363 103211 999366
rect 202229 999363 202295 999366
rect 204713 999363 204779 999366
rect 208853 999363 208919 999366
rect 210417 999363 210483 999366
rect 253657 999426 253723 999429
rect 255313 999426 255379 999429
rect 314702 999426 314762 999499
rect 362217 999426 362283 999429
rect 364701 999426 364767 999429
rect 429653 999426 429719 999429
rect 432873 999426 432939 999429
rect 506657 999426 506723 999429
rect 509049 999426 509115 999429
rect 556797 999426 556863 999429
rect 557165 999426 557231 999429
rect 253657 999424 253920 999426
rect 253657 999368 253662 999424
rect 253718 999368 253920 999424
rect 253657 999366 253920 999368
rect 255313 999424 255576 999426
rect 255313 999368 255318 999424
rect 255374 999368 255576 999424
rect 255313 999366 255576 999368
rect 314548 999366 314762 999426
rect 362020 999424 362283 999426
rect 362020 999368 362222 999424
rect 362278 999368 362283 999424
rect 362020 999366 362283 999368
rect 364504 999424 364767 999426
rect 364504 999368 364706 999424
rect 364762 999368 364767 999424
rect 364504 999366 364767 999368
rect 429456 999424 429719 999426
rect 429456 999368 429658 999424
rect 429714 999368 429719 999424
rect 429456 999366 429719 999368
rect 432676 999424 432939 999426
rect 432676 999368 432878 999424
rect 432934 999368 432939 999424
rect 432676 999366 432939 999368
rect 506460 999424 506723 999426
rect 506460 999368 506662 999424
rect 506718 999368 506723 999424
rect 506460 999366 506723 999368
rect 508852 999424 509115 999426
rect 508852 999368 509054 999424
rect 509110 999368 509115 999424
rect 508852 999366 509115 999368
rect 556600 999424 556863 999426
rect 556600 999368 556802 999424
rect 556858 999368 556863 999424
rect 556600 999366 556863 999368
rect 557060 999424 557231 999426
rect 557060 999368 557170 999424
rect 557226 999368 557231 999424
rect 557060 999366 557231 999368
rect 253657 999363 253723 999366
rect 255313 999363 255379 999366
rect 362217 999363 362283 999366
rect 364701 999363 364767 999366
rect 429653 999363 429719 999366
rect 432873 999363 432939 999366
rect 506657 999363 506723 999366
rect 509049 999363 509115 999366
rect 556797 999363 556863 999366
rect 557165 999363 557231 999366
rect 100293 999290 100359 999293
rect 101121 999290 101187 999293
rect 202689 999290 202755 999293
rect 205173 999290 205239 999293
rect 209589 999290 209655 999293
rect 211705 999290 211771 999293
rect 100293 999288 100556 999290
rect 100293 999232 100298 999288
rect 100354 999232 100556 999288
rect 100293 999230 100556 999232
rect 101121 999288 101292 999290
rect 101121 999232 101126 999288
rect 101182 999232 101292 999288
rect 101121 999230 101292 999232
rect 202689 999288 202952 999290
rect 202689 999232 202694 999288
rect 202750 999232 202952 999288
rect 202689 999230 202952 999232
rect 205173 999288 205344 999290
rect 205173 999232 205178 999288
rect 205234 999232 205344 999288
rect 205173 999230 205344 999232
rect 209484 999288 209655 999290
rect 209484 999232 209594 999288
rect 209650 999232 209655 999288
rect 209484 999230 209655 999232
rect 211508 999288 211771 999290
rect 211508 999232 211710 999288
rect 211766 999232 211771 999288
rect 211508 999230 211771 999232
rect 100293 999227 100359 999230
rect 101121 999227 101187 999230
rect 202689 999227 202755 999230
rect 205173 999227 205239 999230
rect 209589 999227 209655 999230
rect 211705 999227 211771 999230
rect 254485 999290 254551 999293
rect 256509 999290 256575 999293
rect 364241 999290 364307 999293
rect 365437 999290 365503 999293
rect 430389 999290 430455 999293
rect 432045 999290 432111 999293
rect 500861 999290 500927 999293
rect 507393 999290 507459 999293
rect 509509 999290 509575 999293
rect 254485 999288 254748 999290
rect 254485 999232 254490 999288
rect 254546 999232 254748 999288
rect 254485 999230 254748 999232
rect 256509 999288 256772 999290
rect 256509 999232 256514 999288
rect 256570 999232 256772 999288
rect 256509 999230 256772 999232
rect 364044 999288 364307 999290
rect 364044 999232 364246 999288
rect 364302 999232 364307 999288
rect 364044 999230 364307 999232
rect 365332 999288 365503 999290
rect 365332 999232 365442 999288
rect 365498 999232 365503 999288
rect 365332 999230 365503 999232
rect 430284 999288 430455 999290
rect 430284 999232 430394 999288
rect 430450 999232 430455 999288
rect 430284 999230 430455 999232
rect 431940 999288 432111 999290
rect 431940 999232 432050 999288
rect 432106 999232 432111 999288
rect 431940 999230 432111 999232
rect 500756 999288 500927 999290
rect 500756 999232 500866 999288
rect 500922 999232 500927 999288
rect 500756 999230 500927 999232
rect 507196 999288 507459 999290
rect 507196 999232 507398 999288
rect 507454 999232 507459 999288
rect 507196 999230 507459 999232
rect 509312 999288 509575 999290
rect 509312 999232 509514 999288
rect 509570 999232 509575 999288
rect 509312 999230 509575 999232
rect 254485 999227 254551 999230
rect 256509 999227 256575 999230
rect 364241 999227 364307 999230
rect 365437 999227 365503 999230
rect 430389 999227 430455 999230
rect 432045 999227 432111 999230
rect 500861 999227 500927 999230
rect 507393 999227 507459 999230
rect 509509 999227 509575 999230
rect 519997 999290 520063 999293
rect 523861 999290 523927 999293
rect 519997 999288 523927 999290
rect 519997 999232 520002 999288
rect 520058 999232 523866 999288
rect 523922 999232 523927 999288
rect 519997 999230 523927 999232
rect 519997 999227 520063 999230
rect 523861 999227 523927 999230
rect 554313 999290 554379 999293
rect 558821 999290 558887 999293
rect 559649 999290 559715 999293
rect 561305 999290 561371 999293
rect 554313 999288 554576 999290
rect 554313 999232 554318 999288
rect 554374 999232 554576 999288
rect 554313 999230 554576 999232
rect 558624 999288 558887 999290
rect 558624 999232 558826 999288
rect 558882 999232 558887 999288
rect 558624 999230 558887 999232
rect 559452 999288 559715 999290
rect 559452 999232 559654 999288
rect 559710 999232 559715 999288
rect 559452 999230 559715 999232
rect 561108 999288 561371 999290
rect 561108 999232 561310 999288
rect 561366 999232 561371 999288
rect 561108 999230 561371 999232
rect 554313 999227 554379 999230
rect 558821 999227 558887 999230
rect 559649 999227 559715 999230
rect 561305 999227 561371 999230
rect 99925 999154 99991 999157
rect 155769 999154 155835 999157
rect 158253 999154 158319 999157
rect 203057 999154 203123 999157
rect 207565 999154 207631 999157
rect 211245 999154 211311 999157
rect 99925 999152 100096 999154
rect 99925 999096 99930 999152
rect 99986 999096 100096 999152
rect 99925 999094 100096 999096
rect 155769 999152 156032 999154
rect 155769 999096 155774 999152
rect 155830 999096 156032 999152
rect 155769 999094 156032 999096
rect 158253 999152 158516 999154
rect 158253 999096 158258 999152
rect 158314 999096 158516 999152
rect 158253 999094 158516 999096
rect 203057 999152 203320 999154
rect 203057 999096 203062 999152
rect 203118 999096 203320 999152
rect 203057 999094 203320 999096
rect 207565 999152 207828 999154
rect 207565 999096 207570 999152
rect 207626 999096 207828 999152
rect 207565 999094 207828 999096
rect 211140 999152 211311 999154
rect 211140 999096 211250 999152
rect 211306 999096 211311 999152
rect 211140 999094 211311 999096
rect 99925 999091 99991 999094
rect 155769 999091 155835 999094
rect 158253 999091 158319 999094
rect 203057 999091 203123 999094
rect 207565 999091 207631 999094
rect 211245 999091 211311 999094
rect 254117 999154 254183 999157
rect 258533 999154 258599 999157
rect 254117 999152 254380 999154
rect 254117 999096 254122 999152
rect 254178 999096 254380 999152
rect 254117 999094 254380 999096
rect 258428 999152 258599 999154
rect 258428 999096 258538 999152
rect 258594 999096 258599 999152
rect 258428 999094 258599 999096
rect 254117 999091 254183 999094
rect 258533 999091 258599 999094
rect 312629 999154 312695 999157
rect 358905 999154 358971 999157
rect 363045 999154 363111 999157
rect 437381 999154 437447 999157
rect 312629 999152 312892 999154
rect 312629 999096 312634 999152
rect 312690 999096 312892 999152
rect 312629 999094 312892 999096
rect 358905 999152 359168 999154
rect 358905 999096 358910 999152
rect 358966 999096 359168 999152
rect 358905 999094 359168 999096
rect 362848 999152 363111 999154
rect 362848 999096 363050 999152
rect 363106 999096 363111 999152
rect 362848 999094 363111 999096
rect 433136 999152 437447 999154
rect 433136 999096 437386 999152
rect 437442 999096 437447 999152
rect 433136 999094 437447 999096
rect 312629 999091 312695 999094
rect 358905 999091 358971 999094
rect 363045 999091 363111 999094
rect 437381 999091 437447 999094
rect 503345 999154 503411 999157
rect 509877 999154 509943 999157
rect 513624 999154 513690 999157
rect 517237 999154 517303 999157
rect 524045 999154 524111 999157
rect 503345 999152 503608 999154
rect 503345 999096 503350 999152
rect 503406 999096 503608 999152
rect 503345 999094 503608 999096
rect 509680 999152 509943 999154
rect 509680 999096 509882 999152
rect 509938 999096 509943 999152
rect 509680 999094 509943 999096
rect 510140 999152 513699 999154
rect 510140 999096 513629 999152
rect 513685 999096 513699 999152
rect 510140 999094 513699 999096
rect 517237 999152 524111 999154
rect 517237 999096 517242 999152
rect 517298 999096 524050 999152
rect 524106 999096 524111 999152
rect 517237 999094 524111 999096
rect 503345 999091 503411 999094
rect 509877 999091 509943 999094
rect 513624 999091 513690 999094
rect 517237 999091 517303 999094
rect 524045 999091 524111 999094
rect 551921 999154 551987 999157
rect 557625 999154 557691 999157
rect 551921 999152 552092 999154
rect 551921 999096 551926 999152
rect 551982 999096 552092 999152
rect 551921 999094 552092 999096
rect 557428 999152 557691 999154
rect 557428 999096 557630 999152
rect 557686 999096 557691 999152
rect 557428 999094 557691 999096
rect 551921 999091 551987 999094
rect 557625 999091 557691 999094
rect 156137 997794 156203 997797
rect 156137 997792 156400 997794
rect 156137 997736 156142 997792
rect 156198 997736 156400 997792
rect 156137 997734 156400 997736
rect 156137 997731 156203 997734
rect 107653 997250 107719 997253
rect 107456 997248 107719 997250
rect 107456 997192 107658 997248
rect 107714 997192 107719 997248
rect 107456 997190 107719 997192
rect 107653 997187 107719 997190
rect 115933 997250 115999 997253
rect 143993 997250 144059 997253
rect 115933 997248 144059 997250
rect 115933 997192 115938 997248
rect 115994 997192 143998 997248
rect 144054 997192 144059 997248
rect 115933 997190 144059 997192
rect 115933 997187 115999 997190
rect 143993 997187 144059 997190
rect 187734 997188 187740 997252
rect 187804 997250 187810 997252
rect 195145 997250 195211 997253
rect 187804 997248 195211 997250
rect 187804 997192 195150 997248
rect 195206 997192 195211 997248
rect 187804 997190 195211 997192
rect 187804 997188 187810 997190
rect 195145 997187 195211 997190
rect 218965 997250 219031 997253
rect 247953 997250 248019 997253
rect 218965 997248 248019 997250
rect 218965 997192 218970 997248
rect 219026 997192 247958 997248
rect 248014 997192 248019 997248
rect 218965 997190 248019 997192
rect 218965 997187 219031 997190
rect 247953 997187 248019 997190
rect 270461 997250 270527 997253
rect 298737 997250 298803 997253
rect 270461 997248 298803 997250
rect 270461 997192 270466 997248
rect 270522 997192 298742 997248
rect 298798 997192 298803 997248
rect 270461 997190 298803 997192
rect 270461 997187 270527 997190
rect 298737 997187 298803 997190
rect 368933 997250 368999 997253
rect 399937 997250 400003 997253
rect 368933 997248 369113 997250
rect 368933 997192 368938 997248
rect 368994 997192 369113 997248
rect 368933 997187 369113 997192
rect 168853 997114 168919 997117
rect 195329 997114 195395 997117
rect 168853 997112 195395 997114
rect 168853 997056 168858 997112
rect 168914 997056 195334 997112
rect 195390 997056 195395 997112
rect 168853 997054 195395 997056
rect 168853 997051 168919 997054
rect 195329 997051 195395 997054
rect 95693 996434 95759 996437
rect 148133 996434 148199 996437
rect 87830 996432 95759 996434
rect 87830 996376 95698 996432
rect 95754 996376 95759 996432
rect 87830 996374 95759 996376
rect 87830 995757 87890 996374
rect 95693 996371 95759 996374
rect 142846 996432 148199 996434
rect 142846 996376 148138 996432
rect 148194 996376 148199 996432
rect 142846 996374 148199 996376
rect 108481 996162 108547 996165
rect 108284 996160 108547 996162
rect 87781 995752 87890 995757
rect 87781 995696 87786 995752
rect 87842 995696 87890 995752
rect 87781 995694 87890 995696
rect 87781 995691 87847 995694
rect 85297 995618 85363 995621
rect 95509 995618 95575 995621
rect 85297 995616 95575 995618
rect 85297 995560 85302 995616
rect 85358 995560 95514 995616
rect 95570 995560 95575 995616
rect 85297 995558 95575 995560
rect 85297 995555 85363 995558
rect 95509 995555 95575 995558
rect 97349 995618 97415 995621
rect 103746 995618 103806 996132
rect 104206 995621 104266 996132
rect 97349 995616 103806 995618
rect 97349 995560 97354 995616
rect 97410 995560 103806 995616
rect 97349 995558 103806 995560
rect 104157 995616 104266 995621
rect 104157 995560 104162 995616
rect 104218 995560 104266 995616
rect 104157 995558 104266 995560
rect 104341 995618 104407 995621
rect 104942 995618 105002 996132
rect 104341 995616 105002 995618
rect 104341 995560 104346 995616
rect 104402 995560 105002 995616
rect 104341 995558 105002 995560
rect 97349 995555 97415 995558
rect 104157 995555 104223 995558
rect 104341 995555 104407 995558
rect 82353 995482 82419 995485
rect 95325 995482 95391 995485
rect 82353 995480 95391 995482
rect 82353 995424 82358 995480
rect 82414 995424 95330 995480
rect 95386 995424 95391 995480
rect 82353 995422 95391 995424
rect 105862 995482 105922 996132
rect 106598 995618 106658 996132
rect 107058 995754 107118 996132
rect 108284 996104 108486 996160
rect 108542 996104 108547 996160
rect 108284 996102 108547 996104
rect 108481 996099 108547 996102
rect 108622 995890 108682 996132
rect 113265 995890 113331 995893
rect 108622 995888 113331 995890
rect 108622 995832 113270 995888
rect 113326 995832 113331 995888
rect 108622 995830 113331 995832
rect 113265 995827 113331 995830
rect 142846 995757 142906 996374
rect 148133 996371 148199 996374
rect 305729 996298 305795 996301
rect 308121 996298 308187 996301
rect 305729 996296 305900 996298
rect 305729 996240 305734 996296
rect 305790 996240 305900 996296
rect 305729 996238 305900 996240
rect 308121 996296 308384 996298
rect 308121 996240 308126 996296
rect 308182 996240 308384 996296
rect 308121 996238 308384 996240
rect 305729 996235 305795 996238
rect 308121 996235 308187 996238
rect 305269 996162 305335 996165
rect 306465 996162 306531 996165
rect 306925 996162 306991 996165
rect 307293 996162 307359 996165
rect 307753 996162 307819 996165
rect 309317 996162 309383 996165
rect 310145 996162 310211 996165
rect 310605 996162 310671 996165
rect 311801 996162 311867 996165
rect 314285 996162 314351 996165
rect 305269 996160 305532 996162
rect 156965 996157 157031 996160
rect 157793 996157 157859 996160
rect 159449 996157 159515 996160
rect 156965 996155 157228 996157
rect 156965 996099 156970 996155
rect 157026 996099 157228 996155
rect 156965 996097 157228 996099
rect 157793 996155 158056 996157
rect 157793 996099 157798 996155
rect 157854 996127 158056 996155
rect 159449 996155 159712 996157
rect 157854 996099 158086 996127
rect 157793 996097 158086 996099
rect 156965 996094 157031 996097
rect 157793 996094 157859 996097
rect 110413 995754 110479 995757
rect 107058 995752 110479 995754
rect 107058 995696 110418 995752
rect 110474 995696 110479 995752
rect 107058 995694 110479 995696
rect 110413 995691 110479 995694
rect 142797 995752 142906 995757
rect 142797 995696 142802 995752
rect 142858 995696 142906 995752
rect 142797 995694 142906 995696
rect 142797 995691 142863 995694
rect 110505 995618 110571 995621
rect 106598 995616 110571 995618
rect 106598 995560 110510 995616
rect 110566 995560 110571 995616
rect 106598 995558 110571 995560
rect 110505 995555 110571 995558
rect 137369 995618 137435 995621
rect 147581 995618 147647 995621
rect 137369 995616 147647 995618
rect 137369 995560 137374 995616
rect 137430 995560 147586 995616
rect 147642 995560 147647 995616
rect 137369 995558 147647 995560
rect 158026 995618 158086 996097
rect 159449 996099 159454 996155
rect 159510 996127 159712 996155
rect 159510 996099 159742 996127
rect 159449 996097 159742 996099
rect 159449 996094 159515 996097
rect 159682 995754 159742 996097
rect 160050 995890 160110 996127
rect 160050 995830 164059 995890
rect 162945 995754 163011 995757
rect 159682 995752 163011 995754
rect 159682 995696 162950 995752
rect 163006 995696 163011 995752
rect 159682 995694 163011 995696
rect 162945 995691 163011 995694
rect 162853 995618 162919 995621
rect 158026 995616 162919 995618
rect 158026 995560 162858 995616
rect 162914 995560 162919 995616
rect 158026 995558 162919 995560
rect 137369 995555 137435 995558
rect 147581 995555 147647 995558
rect 162853 995555 162919 995558
rect 110597 995482 110663 995485
rect 105862 995480 110663 995482
rect 105862 995424 110602 995480
rect 110658 995424 110663 995480
rect 105862 995422 110663 995424
rect 82353 995419 82419 995422
rect 95325 995419 95391 995422
rect 110597 995419 110663 995422
rect 133689 995482 133755 995485
rect 143993 995482 144059 995485
rect 133689 995480 144059 995482
rect 133689 995424 133694 995480
rect 133750 995424 143998 995480
rect 144054 995424 144059 995480
rect 133689 995422 144059 995424
rect 133689 995419 133755 995422
rect 143993 995419 144059 995422
rect 81617 995346 81683 995349
rect 95141 995346 95207 995349
rect 81617 995344 95207 995346
rect 81617 995288 81622 995344
rect 81678 995288 95146 995344
rect 95202 995288 95207 995344
rect 81617 995286 95207 995288
rect 81617 995283 81683 995286
rect 95141 995283 95207 995286
rect 80697 995210 80763 995213
rect 92769 995210 92835 995213
rect 80697 995208 92835 995210
rect 80697 995152 80702 995208
rect 80758 995152 92774 995208
rect 92830 995152 92835 995208
rect 80697 995150 92835 995152
rect 80697 995147 80763 995150
rect 92769 995147 92835 995150
rect 84469 994122 84535 994125
rect 97901 994122 97967 994125
rect 84469 994120 97967 994122
rect 84469 994064 84474 994120
rect 84530 994064 97906 994120
rect 97962 994064 97967 994120
rect 84469 994062 97967 994064
rect 84469 994059 84535 994062
rect 97901 994059 97967 994062
rect 80145 993850 80211 993853
rect 97349 993850 97415 993853
rect 80145 993848 97415 993850
rect 80145 993792 80150 993848
rect 80206 993792 97354 993848
rect 97410 993792 97415 993848
rect 80145 993790 97415 993792
rect 80145 993787 80211 993790
rect 97349 993787 97415 993790
rect 163999 993730 164059 995830
rect 187601 995754 187667 995757
rect 187734 995754 187740 995756
rect 187601 995752 187740 995754
rect 187601 995696 187606 995752
rect 187662 995696 187740 995752
rect 187601 995694 187740 995696
rect 187601 995691 187667 995694
rect 187734 995692 187740 995694
rect 187804 995692 187810 995756
rect 192477 995618 192543 995621
rect 207430 995618 207490 996132
rect 250437 996026 250503 996029
rect 240182 996024 250503 996026
rect 240182 995968 250442 996024
rect 250498 995968 250503 996024
rect 240182 995966 250503 995968
rect 240182 995890 240242 995966
rect 250437 995963 250503 995966
rect 250253 995890 250319 995893
rect 235766 995830 240242 995890
rect 240550 995888 250319 995890
rect 240550 995832 250258 995888
rect 250314 995832 250319 995888
rect 240550 995830 250319 995832
rect 235257 995754 235323 995757
rect 235766 995754 235826 995830
rect 235257 995752 235826 995754
rect 235257 995696 235262 995752
rect 235318 995696 235826 995752
rect 235257 995694 235826 995696
rect 235901 995754 235967 995757
rect 240550 995754 240610 995830
rect 250253 995827 250319 995830
rect 235901 995752 240610 995754
rect 235901 995696 235906 995752
rect 235962 995696 240610 995752
rect 235901 995694 240610 995696
rect 242065 995754 242131 995757
rect 250069 995754 250135 995757
rect 242065 995752 250135 995754
rect 242065 995696 242070 995752
rect 242126 995696 250074 995752
rect 250130 995696 250135 995752
rect 242065 995694 250135 995696
rect 235257 995691 235323 995694
rect 235901 995691 235967 995694
rect 242065 995691 242131 995694
rect 250069 995691 250135 995694
rect 192477 995616 207490 995618
rect 192477 995560 192482 995616
rect 192538 995560 207490 995616
rect 192477 995558 207490 995560
rect 240041 995618 240107 995621
rect 249701 995618 249767 995621
rect 240041 995616 249767 995618
rect 240041 995560 240046 995616
rect 240102 995560 249706 995616
rect 249762 995560 249767 995616
rect 240041 995558 249767 995560
rect 192477 995555 192543 995558
rect 240041 995555 240107 995558
rect 249701 995555 249767 995558
rect 236545 995482 236611 995485
rect 249885 995482 249951 995485
rect 236545 995480 249951 995482
rect 236545 995424 236550 995480
rect 236606 995424 249890 995480
rect 249946 995424 249951 995480
rect 236545 995422 249951 995424
rect 236545 995419 236611 995422
rect 249885 995419 249951 995422
rect 234383 995346 234449 995349
rect 246849 995346 246915 995349
rect 234383 995344 246915 995346
rect 234383 995288 234388 995344
rect 234444 995288 246854 995344
rect 246910 995288 246915 995344
rect 234383 995286 246915 995288
rect 234383 995283 234449 995286
rect 246849 995283 246915 995286
rect 232221 994122 232287 994125
rect 252461 994122 252527 994125
rect 232221 994120 252527 994122
rect 232221 994064 232226 994120
rect 232282 994064 252466 994120
rect 252522 994064 252527 994120
rect 232221 994062 252527 994064
rect 232221 994059 232287 994062
rect 252461 994059 252527 994062
rect 232865 993986 232931 993989
rect 259134 993986 259194 996132
rect 300761 995890 300827 995893
rect 303846 995890 303906 996132
rect 305134 995890 305194 996132
rect 305269 996104 305274 996160
rect 305330 996104 305532 996160
rect 306465 996160 306728 996162
rect 305269 996102 305532 996104
rect 305269 996099 305335 996102
rect 306330 995890 306390 996132
rect 306465 996104 306470 996160
rect 306526 996104 306728 996160
rect 306465 996102 306728 996104
rect 306925 996160 307188 996162
rect 306925 996104 306930 996160
rect 306986 996104 307188 996160
rect 306925 996102 307188 996104
rect 307293 996160 307556 996162
rect 307293 996104 307298 996160
rect 307354 996104 307556 996160
rect 307293 996102 307556 996104
rect 307753 996160 307924 996162
rect 307753 996104 307758 996160
rect 307814 996104 307924 996160
rect 309317 996160 309580 996162
rect 307753 996102 307924 996104
rect 306465 996099 306531 996102
rect 306925 996099 306991 996102
rect 307293 996099 307359 996102
rect 307753 996099 307819 996102
rect 292254 995830 300594 995890
rect 288065 995754 288131 995757
rect 292254 995754 292314 995830
rect 288065 995752 292314 995754
rect 288065 995696 288070 995752
rect 288126 995696 292314 995752
rect 288065 995694 292314 995696
rect 292481 995754 292547 995757
rect 300534 995754 300594 995830
rect 300761 995888 305194 995890
rect 300761 995832 300766 995888
rect 300822 995832 305194 995888
rect 300761 995830 305194 995832
rect 305318 995830 306390 995890
rect 300761 995827 300827 995830
rect 305318 995754 305378 995830
rect 292481 995752 300410 995754
rect 292481 995696 292486 995752
rect 292542 995696 300410 995752
rect 292481 995694 300410 995696
rect 300534 995694 305378 995754
rect 288065 995691 288131 995694
rect 292481 995691 292547 995694
rect 291101 995618 291167 995621
rect 300209 995618 300275 995621
rect 291101 995616 300275 995618
rect 291101 995560 291106 995616
rect 291162 995560 300214 995616
rect 300270 995560 300275 995616
rect 291101 995558 300275 995560
rect 300350 995618 300410 995694
rect 305269 995618 305335 995621
rect 300350 995616 305335 995618
rect 300350 995560 305274 995616
rect 305330 995560 305335 995616
rect 300350 995558 305335 995560
rect 291101 995555 291167 995558
rect 300209 995555 300275 995558
rect 305269 995555 305335 995558
rect 290549 995482 290615 995485
rect 297265 995482 297331 995485
rect 308722 995482 308782 996132
rect 290549 995480 295350 995482
rect 290549 995424 290554 995480
rect 290610 995424 295350 995480
rect 290549 995422 295350 995424
rect 290549 995419 290615 995422
rect 295290 995346 295350 995422
rect 297265 995480 308782 995482
rect 297265 995424 297270 995480
rect 297326 995424 308782 995480
rect 297265 995422 308782 995424
rect 297265 995419 297331 995422
rect 309182 995346 309242 996132
rect 309317 996104 309322 996160
rect 309378 996104 309580 996160
rect 309317 996102 309580 996104
rect 310145 996160 310408 996162
rect 310145 996104 310150 996160
rect 310206 996104 310408 996160
rect 310145 996102 310408 996104
rect 310605 996160 310868 996162
rect 310605 996104 310610 996160
rect 310666 996104 310868 996160
rect 310605 996102 310868 996104
rect 311604 996160 311867 996162
rect 311604 996104 311806 996160
rect 311862 996104 311867 996160
rect 311604 996102 311867 996104
rect 314088 996160 314351 996162
rect 314088 996104 314290 996160
rect 314346 996104 314351 996160
rect 314088 996102 314351 996104
rect 315284 996102 318550 996162
rect 309317 996099 309383 996102
rect 310145 996099 310211 996102
rect 310605 996099 310671 996102
rect 311801 996099 311867 996102
rect 314285 996099 314351 996102
rect 295290 995286 309242 995346
rect 232865 993984 259194 993986
rect 232865 993928 232870 993984
rect 232926 993928 259194 993984
rect 232865 993926 259194 993928
rect 232865 993923 232931 993926
rect 318490 993919 318550 996102
rect 318490 993859 319969 993919
rect 243261 993850 243327 993853
rect 316769 993850 316835 993853
rect 243261 993848 268540 993850
rect 243261 993792 243266 993848
rect 243322 993792 268540 993848
rect 243261 993790 268540 993792
rect 243261 993787 243327 993790
rect 268480 993733 268540 993790
rect 270945 993848 316835 993850
rect 270945 993792 316774 993848
rect 316830 993792 316835 993848
rect 270945 993790 316835 993792
rect 270945 993733 271005 993790
rect 316769 993787 316835 993790
rect 168373 993730 168439 993733
rect 163999 993728 168439 993730
rect 78305 993714 78371 993717
rect 104341 993714 104407 993717
rect 78305 993712 104407 993714
rect 78305 993656 78310 993712
rect 78366 993656 104346 993712
rect 104402 993656 104407 993712
rect 163999 993672 168378 993728
rect 168434 993672 168439 993728
rect 163999 993670 168439 993672
rect 168373 993667 168439 993670
rect 191833 993714 191899 993717
rect 248321 993714 248387 993717
rect 191833 993712 248387 993714
rect 78305 993654 104407 993656
rect 78305 993651 78371 993654
rect 104341 993651 104407 993654
rect 191833 993656 191838 993712
rect 191894 993656 248326 993712
rect 248382 993656 248387 993712
rect 268480 993673 271005 993733
rect 294505 993714 294571 993717
rect 294505 993712 319744 993714
rect 191833 993654 248387 993656
rect 191833 993651 191899 993654
rect 248321 993651 248387 993654
rect 294505 993656 294510 993712
rect 294566 993656 319744 993712
rect 294505 993654 319744 993656
rect 294505 993651 294571 993654
rect 319684 993376 319744 993654
rect 319909 993582 319969 993859
rect 366173 993714 366239 993717
rect 322820 993712 366239 993714
rect 322820 993656 366178 993712
rect 366234 993656 366239 993712
rect 322820 993654 366239 993656
rect 321461 993582 321527 993585
rect 319909 993580 321527 993582
rect 319909 993524 321466 993580
rect 321522 993524 321527 993580
rect 319909 993522 321527 993524
rect 321461 993519 321527 993522
rect 322820 993376 322880 993654
rect 366173 993651 366239 993654
rect 369053 993641 369113 997187
rect 372889 997248 400003 997250
rect 372889 997192 399942 997248
rect 399998 997192 400003 997248
rect 372889 997190 400003 997192
rect 372889 993641 372949 997190
rect 399937 997187 400003 997190
rect 439817 997250 439883 997253
rect 488901 997250 488967 997253
rect 439817 997248 488967 997250
rect 439817 997192 439822 997248
rect 439878 997192 488906 997248
rect 488962 997192 488967 997248
rect 439817 997190 488967 997192
rect 439817 997187 439883 997190
rect 488901 997187 488967 997190
rect 523861 996570 523927 996573
rect 523861 996568 528570 996570
rect 523861 996512 523866 996568
rect 523922 996512 528570 996568
rect 523861 996510 528570 996512
rect 523861 996507 523927 996510
rect 383091 996434 383157 996437
rect 524045 996434 524111 996437
rect 383091 996432 388178 996434
rect 383091 996376 383096 996432
rect 383152 996376 388178 996432
rect 383091 996374 388178 996376
rect 383091 996371 383157 996374
rect 388118 995757 388178 996374
rect 524045 996432 528018 996434
rect 524045 996376 524050 996432
rect 524106 996376 528018 996432
rect 524045 996374 528018 996376
rect 524045 996371 524111 996374
rect 527958 995757 528018 996374
rect 528510 995757 528570 996510
rect 388118 995752 388227 995757
rect 388118 995696 388166 995752
rect 388222 995696 388227 995752
rect 388118 995694 388227 995696
rect 388161 995691 388227 995694
rect 447317 995754 447383 995757
rect 481449 995754 481515 995757
rect 447317 995752 481515 995754
rect 447317 995696 447322 995752
rect 447378 995696 481454 995752
rect 481510 995696 481515 995752
rect 447317 995694 481515 995696
rect 447317 995691 447383 995694
rect 481449 995691 481515 995694
rect 520181 995754 520247 995757
rect 525425 995754 525491 995757
rect 520181 995752 525491 995754
rect 520181 995696 520186 995752
rect 520242 995696 525430 995752
rect 525486 995696 525491 995752
rect 520181 995694 525491 995696
rect 527958 995752 528067 995757
rect 527958 995696 528006 995752
rect 528062 995696 528067 995752
rect 527958 995694 528067 995696
rect 528510 995752 528619 995757
rect 528510 995696 528558 995752
rect 528614 995696 528619 995752
rect 528510 995694 528619 995696
rect 520181 995691 520247 995694
rect 525425 995691 525491 995694
rect 528001 995691 528067 995694
rect 528553 995691 528619 995694
rect 517605 995618 517671 995621
rect 526069 995618 526135 995621
rect 517605 995616 526135 995618
rect 517605 995560 517610 995616
rect 517666 995560 526074 995616
rect 526130 995560 526135 995616
rect 517605 995558 526135 995560
rect 517605 995555 517671 995558
rect 526069 995555 526135 995558
rect 520365 995482 520431 995485
rect 532141 995482 532207 995485
rect 520365 995480 532207 995482
rect 520365 995424 520370 995480
rect 520426 995424 532146 995480
rect 532202 995424 532207 995480
rect 520365 995422 532207 995424
rect 520365 995419 520431 995422
rect 532141 995419 532207 995422
rect 638539 995212 638605 995213
rect 638534 995210 638540 995212
rect 638448 995150 638540 995210
rect 638534 995148 638540 995150
rect 638604 995148 638610 995212
rect 638539 995147 638605 995148
rect 575565 994258 575631 994261
rect 634813 994258 634879 994261
rect 575565 994256 634879 994258
rect 575565 994200 575570 994256
rect 575626 994200 634818 994256
rect 634874 994200 634879 994256
rect 575565 994198 634879 994200
rect 575565 994195 575631 994198
rect 634813 994195 634879 994198
rect 571333 994122 571399 994125
rect 637021 994122 637087 994125
rect 571333 994120 637087 994122
rect 571333 994064 571338 994120
rect 571394 994064 637026 994120
rect 637082 994064 637087 994120
rect 571333 994062 637087 994064
rect 571333 994059 571399 994062
rect 637021 994059 637087 994062
rect 629661 993986 629727 993989
rect 568285 993984 629727 993986
rect 568285 993928 629666 993984
rect 629722 993928 629727 993984
rect 568285 993926 629727 993928
rect 378133 993850 378199 993853
rect 396993 993850 397059 993853
rect 378133 993848 397059 993850
rect 378133 993792 378138 993848
rect 378194 993792 396998 993848
rect 397054 993792 397059 993848
rect 378133 993790 397059 993792
rect 378133 993787 378199 993790
rect 396993 993787 397059 993790
rect 567009 993746 567075 993749
rect 568285 993746 568345 993926
rect 629661 993923 629727 993926
rect 569953 993850 570019 993853
rect 635181 993850 635247 993853
rect 569953 993848 635247 993850
rect 569953 993792 569958 993848
rect 570014 993792 635186 993848
rect 635242 993792 635247 993848
rect 569953 993790 635247 993792
rect 569953 993787 570019 993790
rect 635181 993787 635247 993790
rect 567009 993744 568345 993746
rect 375189 993714 375255 993717
rect 395153 993714 395219 993717
rect 375189 993712 395219 993714
rect 375189 993656 375194 993712
rect 375250 993656 395158 993712
rect 395214 993656 395219 993712
rect 375189 993654 395219 993656
rect 375189 993651 375255 993654
rect 395153 993651 395219 993654
rect 447133 993714 447199 993717
rect 478597 993714 478663 993717
rect 447133 993712 478663 993714
rect 447133 993656 447138 993712
rect 447194 993656 478602 993712
rect 478658 993656 478663 993712
rect 447133 993654 478663 993656
rect 447133 993651 447199 993654
rect 478597 993651 478663 993654
rect 517421 993714 517487 993717
rect 537385 993714 537451 993717
rect 517421 993712 537451 993714
rect 517421 993656 517426 993712
rect 517482 993656 537390 993712
rect 537446 993656 537451 993712
rect 517421 993654 537451 993656
rect 517421 993651 517487 993654
rect 537385 993651 537451 993654
rect 561765 993714 561831 993717
rect 561765 993712 566124 993714
rect 561765 993656 561770 993712
rect 561826 993656 566124 993712
rect 567009 993688 567014 993744
rect 567070 993688 568345 993744
rect 638861 993714 638927 993717
rect 567009 993686 568345 993688
rect 569216 993712 638927 993714
rect 567009 993683 567075 993686
rect 561765 993654 566124 993656
rect 561765 993651 561831 993654
rect 369053 993581 372949 993641
rect 566064 993438 566124 993654
rect 569216 993656 638866 993712
rect 638922 993656 638927 993712
rect 569216 993654 638927 993656
rect 569216 993438 569276 993654
rect 638861 993651 638927 993654
rect 566064 993378 569276 993438
rect 319684 993316 322880 993376
rect 638534 990524 638540 990588
rect 638604 990586 638610 990588
rect 641161 990586 641227 990589
rect 638604 990584 641227 990586
rect 638604 990528 641166 990584
rect 641222 990528 641227 990584
rect 638604 990526 641227 990528
rect 638604 990524 638610 990526
rect 641161 990523 641227 990526
rect 485313 989498 485379 989501
rect 511441 989498 511507 989501
rect 485313 989496 511507 989498
rect 485313 989440 485318 989496
rect 485374 989440 511446 989496
rect 511502 989440 511507 989496
rect 485313 989438 511507 989440
rect 485313 989435 485379 989438
rect 511441 989435 511507 989438
rect 564433 985962 564499 985965
rect 677166 985962 677172 985964
rect 564433 985960 677172 985962
rect 564433 985904 564438 985960
rect 564494 985904 677172 985960
rect 564433 985902 677172 985904
rect 564433 985899 564499 985902
rect 677166 985900 677172 985902
rect 677236 985900 677242 985964
rect 561029 985826 561095 985829
rect 561581 985826 561647 985829
rect 676982 985826 676988 985828
rect 561029 985824 676988 985826
rect 561029 985768 561034 985824
rect 561090 985768 561586 985824
rect 561642 985768 676988 985824
rect 561029 985766 676988 985768
rect 561029 985763 561095 985766
rect 561581 985763 561647 985766
rect 676982 985764 676988 985766
rect 677052 985764 677058 985828
rect 43662 985628 43668 985692
rect 43732 985690 43738 985692
rect 669129 985690 669195 985693
rect 43732 985688 669195 985690
rect 43732 985632 669134 985688
rect 669190 985632 669195 985688
rect 43732 985630 669195 985632
rect 43732 985628 43738 985630
rect 669129 985627 669195 985630
rect 44030 985492 44036 985556
rect 44100 985554 44106 985556
rect 670417 985554 670483 985557
rect 44100 985552 670483 985554
rect 44100 985496 670422 985552
rect 670478 985496 670483 985552
rect 44100 985494 670483 985496
rect 44100 985492 44106 985494
rect 670417 985491 670483 985494
rect 43478 985356 43484 985420
rect 43548 985418 43554 985420
rect 672533 985418 672599 985421
rect 43548 985416 672599 985418
rect 43548 985360 672538 985416
rect 672594 985360 672599 985416
rect 43548 985358 672599 985360
rect 43548 985356 43554 985358
rect 672533 985355 672599 985358
rect 43846 983044 43852 983108
rect 43916 983106 43922 983108
rect 669037 983106 669103 983109
rect 43916 983104 669103 983106
rect 43916 983048 669042 983104
rect 669098 983048 669103 983104
rect 43916 983046 669103 983048
rect 43916 983044 43922 983046
rect 669037 983043 669103 983046
rect 43294 982908 43300 982972
rect 43364 982970 43370 982972
rect 672625 982970 672691 982973
rect 43364 982968 672691 982970
rect 43364 982912 672630 982968
rect 672686 982912 672691 982968
rect 43364 982910 672691 982912
rect 43364 982908 43370 982910
rect 672625 982907 672691 982910
rect 58433 976034 58499 976037
rect 58433 976032 64492 976034
rect 58433 975976 58438 976032
rect 58494 975976 64492 976032
rect 58433 975974 64492 975976
rect 58433 975971 58499 975974
rect 655513 975898 655579 975901
rect 650164 975896 655579 975898
rect 650164 975840 655518 975896
rect 655574 975840 655579 975896
rect 650164 975838 655579 975840
rect 655513 975835 655579 975838
rect 41454 968764 41460 968828
rect 41524 968826 41530 968828
rect 41781 968826 41847 968829
rect 41524 968824 41847 968826
rect 41524 968768 41786 968824
rect 41842 968768 41847 968824
rect 41524 968766 41847 968768
rect 41524 968764 41530 968766
rect 41781 968763 41847 968766
rect 41638 965092 41644 965156
rect 41708 965154 41714 965156
rect 41781 965154 41847 965157
rect 41708 965152 41847 965154
rect 41708 965096 41786 965152
rect 41842 965096 41847 965152
rect 41708 965094 41847 965096
rect 41708 965092 41714 965094
rect 41781 965091 41847 965094
rect 41781 963388 41847 963389
rect 41781 963384 41828 963388
rect 41892 963386 41898 963388
rect 41781 963328 41786 963384
rect 41781 963324 41828 963328
rect 41892 963326 41938 963386
rect 41892 963324 41898 963326
rect 41781 963323 41847 963324
rect 57973 962978 58039 962981
rect 57973 962976 64492 962978
rect 57973 962920 57978 962976
rect 58034 962920 64492 962976
rect 57973 962918 64492 962920
rect 57973 962915 58039 962918
rect 655697 962570 655763 962573
rect 650164 962568 655763 962570
rect 650164 962512 655702 962568
rect 655758 962512 655763 962568
rect 650164 962510 655763 962512
rect 655697 962507 655763 962510
rect 58433 949922 58499 949925
rect 58433 949920 64492 949922
rect 58433 949864 58438 949920
rect 58494 949864 64492 949920
rect 58433 949862 64492 949864
rect 58433 949859 58499 949862
rect 35801 949514 35867 949517
rect 41822 949514 41828 949516
rect 35801 949512 41828 949514
rect 35801 949456 35806 949512
rect 35862 949456 41828 949512
rect 35801 949454 41828 949456
rect 35801 949451 35867 949454
rect 41822 949452 41828 949454
rect 41892 949452 41898 949516
rect 655789 949378 655855 949381
rect 650164 949376 655855 949378
rect 650164 949320 655794 949376
rect 655850 949320 655855 949376
rect 650164 949318 655855 949320
rect 655789 949315 655855 949318
rect 41505 943938 41571 943941
rect 41462 943936 41571 943938
rect 41462 943880 41510 943936
rect 41566 943880 41571 943936
rect 41462 943875 41571 943880
rect 41462 943500 41522 943875
rect 41781 943122 41847 943125
rect 41492 943120 41847 943122
rect 41492 943064 41786 943120
rect 41842 943064 41847 943120
rect 41492 943062 41847 943064
rect 41781 943059 41847 943062
rect 41781 942714 41847 942717
rect 41492 942712 41847 942714
rect 41492 942656 41786 942712
rect 41842 942656 41847 942712
rect 41492 942654 41847 942656
rect 41781 942651 41847 942654
rect 41873 942306 41939 942309
rect 41492 942304 41939 942306
rect 41492 942248 41878 942304
rect 41934 942248 41939 942304
rect 41492 942246 41939 942248
rect 41873 942243 41939 942246
rect 41965 941898 42031 941901
rect 41492 941896 42031 941898
rect 41492 941840 41970 941896
rect 42026 941840 42031 941896
rect 41492 941838 42031 941840
rect 41965 941835 42031 941838
rect 41781 941490 41847 941493
rect 41492 941488 41847 941490
rect 41492 941432 41786 941488
rect 41842 941432 41847 941488
rect 41492 941430 41847 941432
rect 41781 941427 41847 941430
rect 41873 941082 41939 941085
rect 41492 941080 41939 941082
rect 41492 941024 41878 941080
rect 41934 941024 41939 941080
rect 41492 941022 41939 941024
rect 41873 941019 41939 941022
rect 41492 940614 41752 940674
rect 41692 940541 41752 940614
rect 41689 940536 41755 940541
rect 41689 940480 41694 940536
rect 41750 940480 41755 940536
rect 41689 940475 41755 940480
rect 41965 940266 42031 940269
rect 41492 940264 42031 940266
rect 41492 940208 41970 940264
rect 42026 940208 42031 940264
rect 41492 940206 42031 940208
rect 41965 940203 42031 940206
rect 42977 939858 43043 939861
rect 41492 939856 43043 939858
rect 41492 939800 42982 939856
rect 43038 939800 43043 939856
rect 41492 939798 43043 939800
rect 42977 939795 43043 939798
rect 676262 939725 676322 939964
rect 676262 939720 676371 939725
rect 676262 939664 676310 939720
rect 676366 939664 676371 939720
rect 676262 939662 676371 939664
rect 676305 939659 676371 939662
rect 62297 939450 62363 939453
rect 41492 939448 62363 939450
rect 41492 939392 62302 939448
rect 62358 939392 62363 939448
rect 41492 939390 62363 939392
rect 62297 939387 62363 939390
rect 676121 939314 676187 939317
rect 676262 939314 676322 939556
rect 676121 939312 676322 939314
rect 676121 939256 676126 939312
rect 676182 939256 676322 939312
rect 676121 939254 676322 939256
rect 676121 939251 676187 939254
rect 42333 939042 42399 939045
rect 41492 939040 42399 939042
rect 41492 938984 42338 939040
rect 42394 938984 42399 939040
rect 41492 938982 42399 938984
rect 42333 938979 42399 938982
rect 676262 938909 676322 939148
rect 676213 938904 676322 938909
rect 676213 938848 676218 938904
rect 676274 938848 676322 938904
rect 676213 938846 676322 938848
rect 676213 938843 676279 938846
rect 675661 938770 675727 938773
rect 675661 938768 676292 938770
rect 675661 938712 675666 938768
rect 675722 938712 676292 938768
rect 675661 938710 676292 938712
rect 675661 938707 675727 938710
rect 42793 938634 42859 938637
rect 41492 938632 42859 938634
rect 41492 938576 42798 938632
rect 42854 938576 42859 938632
rect 41492 938574 42859 938576
rect 42793 938571 42859 938574
rect 41965 938498 42031 938501
rect 62481 938498 62547 938501
rect 41965 938496 62547 938498
rect 41965 938440 41970 938496
rect 42026 938440 62486 938496
rect 62542 938440 62547 938496
rect 41965 938438 62547 938440
rect 41965 938435 42031 938438
rect 62481 938435 62547 938438
rect 673862 938300 673868 938364
rect 673932 938362 673938 938364
rect 673932 938302 676292 938362
rect 673932 938300 673938 938302
rect 42241 938226 42307 938229
rect 41492 938224 42307 938226
rect 41492 938168 42246 938224
rect 42302 938168 42307 938224
rect 41492 938166 42307 938168
rect 42241 938163 42307 938166
rect 43161 937818 43227 937821
rect 41492 937816 43227 937818
rect 41492 937760 43166 937816
rect 43222 937760 43227 937816
rect 41492 937758 43227 937760
rect 43161 937755 43227 937758
rect 679022 937685 679082 937924
rect 678973 937680 679082 937685
rect 678973 937624 678978 937680
rect 679034 937624 679082 937680
rect 678973 937622 679082 937624
rect 678973 937619 679039 937622
rect 43069 937410 43135 937413
rect 41492 937408 43135 937410
rect 41492 937352 43074 937408
rect 43130 937352 43135 937408
rect 41492 937350 43135 937352
rect 43069 937347 43135 937350
rect 676814 937276 676874 937516
rect 676806 937212 676812 937276
rect 676876 937212 676882 937276
rect 674966 937076 674972 937140
rect 675036 937138 675042 937140
rect 675036 937078 676292 937138
rect 675036 937076 675042 937078
rect 41822 937002 41828 937004
rect 41492 936942 41828 937002
rect 41822 936940 41828 936942
rect 41892 936940 41898 937004
rect 58433 937002 58499 937005
rect 58433 937000 64492 937002
rect 58433 936944 58438 937000
rect 58494 936944 64492 937000
rect 58433 936942 64492 936944
rect 58433 936939 58499 936942
rect 41781 936594 41847 936597
rect 41492 936592 41847 936594
rect 41492 936536 41786 936592
rect 41842 936536 41847 936592
rect 41492 936534 41847 936536
rect 41781 936531 41847 936534
rect 676262 936461 676322 936700
rect 676213 936456 676322 936461
rect 676213 936400 676218 936456
rect 676274 936400 676322 936456
rect 676213 936398 676322 936400
rect 676213 936395 676279 936398
rect 674782 936260 674788 936324
rect 674852 936322 674858 936324
rect 674852 936262 676292 936322
rect 674852 936260 674858 936262
rect 43345 936186 43411 936189
rect 655605 936186 655671 936189
rect 41492 936184 43411 936186
rect 41492 936128 43350 936184
rect 43406 936128 43411 936184
rect 41492 936126 43411 936128
rect 650164 936184 655671 936186
rect 650164 936128 655610 936184
rect 655666 936128 655671 936184
rect 650164 936126 655671 936128
rect 43345 936123 43411 936126
rect 655605 936123 655671 936126
rect 676029 935914 676095 935917
rect 676029 935912 676292 935914
rect 676029 935856 676034 935912
rect 676090 935856 676292 935912
rect 676029 935854 676292 935856
rect 676029 935851 676095 935854
rect 43253 935778 43319 935781
rect 41492 935776 43319 935778
rect 41492 935720 43258 935776
rect 43314 935720 43319 935776
rect 41492 935718 43319 935720
rect 43253 935715 43319 935718
rect 675937 935506 676003 935509
rect 675937 935504 676292 935506
rect 675937 935448 675942 935504
rect 675998 935448 676292 935504
rect 675937 935446 676292 935448
rect 675937 935443 676003 935446
rect 42006 935370 42012 935372
rect 41492 935310 42012 935370
rect 42006 935308 42012 935310
rect 42076 935308 42082 935372
rect 676029 935098 676095 935101
rect 676029 935096 676292 935098
rect 676029 935040 676034 935096
rect 676090 935040 676292 935096
rect 676029 935038 676292 935040
rect 676029 935035 676095 935038
rect 35801 934962 35867 934965
rect 35788 934960 35867 934962
rect 35788 934904 35806 934960
rect 35862 934904 35867 934960
rect 35788 934902 35867 934904
rect 35801 934899 35867 934902
rect 675845 934690 675911 934693
rect 675845 934688 676292 934690
rect 675845 934632 675850 934688
rect 675906 934632 676292 934688
rect 675845 934630 676292 934632
rect 675845 934627 675911 934630
rect 35709 934554 35775 934557
rect 35709 934552 35788 934554
rect 35709 934496 35714 934552
rect 35770 934496 35788 934552
rect 35709 934494 35788 934496
rect 35709 934491 35775 934494
rect 675937 934282 676003 934285
rect 675937 934280 676292 934282
rect 675937 934224 675942 934280
rect 675998 934224 676292 934280
rect 675937 934222 676292 934224
rect 675937 934219 676003 934222
rect 35617 934146 35683 934149
rect 35604 934144 35683 934146
rect 35604 934088 35622 934144
rect 35678 934088 35683 934144
rect 35604 934086 35683 934088
rect 35617 934083 35683 934086
rect 676121 934010 676187 934013
rect 676121 934008 676322 934010
rect 676121 933952 676126 934008
rect 676182 933952 676322 934008
rect 676121 933950 676322 933952
rect 676121 933947 676187 933950
rect 676262 933844 676322 933950
rect 42885 933738 42951 933741
rect 41492 933736 42951 933738
rect 41492 933680 42890 933736
rect 42946 933680 42951 933736
rect 41492 933678 42951 933680
rect 42885 933675 42951 933678
rect 676029 933466 676095 933469
rect 676029 933464 676292 933466
rect 676029 933408 676034 933464
rect 676090 933408 676292 933464
rect 676029 933406 676292 933408
rect 676029 933403 676095 933406
rect 41781 933330 41847 933333
rect 41492 933328 41847 933330
rect 41492 933272 41786 933328
rect 41842 933272 41847 933328
rect 41492 933270 41847 933272
rect 41781 933267 41847 933270
rect 675753 933058 675819 933061
rect 675753 933056 676292 933058
rect 675753 933000 675758 933056
rect 675814 933000 676292 933056
rect 675753 932998 676292 933000
rect 675753 932995 675819 932998
rect 24902 932484 24962 932910
rect 676121 932786 676187 932789
rect 676121 932784 676322 932786
rect 676121 932728 676126 932784
rect 676182 932728 676322 932784
rect 676121 932726 676322 932728
rect 676121 932723 676187 932726
rect 676262 932620 676322 932726
rect 676121 932378 676187 932381
rect 676121 932376 676322 932378
rect 676121 932320 676126 932376
rect 676182 932320 676322 932376
rect 676121 932318 676322 932320
rect 676121 932315 676187 932318
rect 676262 932212 676322 932318
rect 41781 932106 41847 932109
rect 41492 932104 41847 932106
rect 41492 932048 41786 932104
rect 41842 932048 41847 932104
rect 41492 932046 41847 932048
rect 41781 932043 41847 932046
rect 676029 931834 676095 931837
rect 676029 931832 676292 931834
rect 676029 931776 676034 931832
rect 676090 931776 676292 931832
rect 676029 931774 676292 931776
rect 676029 931771 676095 931774
rect 676029 931426 676095 931429
rect 676029 931424 676292 931426
rect 676029 931368 676034 931424
rect 676090 931368 676292 931424
rect 676029 931366 676292 931368
rect 676029 931363 676095 931366
rect 675937 931018 676003 931021
rect 675937 931016 676292 931018
rect 675937 930960 675942 931016
rect 675998 930960 676292 931016
rect 675937 930958 676292 930960
rect 675937 930955 676003 930958
rect 676121 930746 676187 930749
rect 676121 930744 676322 930746
rect 676121 930688 676126 930744
rect 676182 930688 676322 930744
rect 676121 930686 676322 930688
rect 676121 930683 676187 930686
rect 676262 930580 676322 930686
rect 676029 930202 676095 930205
rect 676029 930200 676292 930202
rect 676029 930144 676034 930200
rect 676090 930144 676292 930200
rect 676029 930142 676292 930144
rect 676029 930139 676095 930142
rect 679022 929525 679082 929764
rect 678973 929520 679082 929525
rect 678973 929464 678978 929520
rect 679034 929464 679082 929520
rect 678973 929462 679082 929464
rect 678973 929459 679039 929462
rect 684542 928948 684602 929356
rect 678973 928706 679039 928709
rect 678973 928704 679082 928706
rect 678973 928648 678978 928704
rect 679034 928648 679082 928704
rect 678973 928643 679082 928648
rect 679022 928540 679082 928643
rect 43294 927148 43300 927212
rect 43364 927210 43370 927212
rect 43805 927210 43871 927213
rect 43364 927208 43871 927210
rect 43364 927152 43810 927208
rect 43866 927152 43871 927208
rect 43364 927150 43871 927152
rect 43364 927148 43370 927150
rect 43805 927147 43871 927150
rect 58433 923810 58499 923813
rect 58433 923808 64492 923810
rect 58433 923752 58438 923808
rect 58494 923752 64492 923808
rect 58433 923750 64492 923752
rect 58433 923747 58499 923750
rect 654869 922722 654935 922725
rect 650164 922720 654935 922722
rect 650164 922664 654874 922720
rect 654930 922664 654935 922720
rect 650164 922662 654935 922664
rect 654869 922659 654935 922662
rect 42793 922042 42859 922045
rect 43478 922042 43484 922044
rect 42793 922040 43484 922042
rect 42793 921984 42798 922040
rect 42854 921984 43484 922040
rect 42793 921982 43484 921984
rect 42793 921979 42859 921982
rect 43478 921980 43484 921982
rect 43548 921980 43554 922044
rect 59169 910754 59235 910757
rect 59169 910752 64492 910754
rect 59169 910696 59174 910752
rect 59230 910696 64492 910752
rect 59169 910694 64492 910696
rect 59169 910691 59235 910694
rect 654869 909530 654935 909533
rect 650164 909528 654935 909530
rect 650164 909472 654874 909528
rect 654930 909472 654935 909528
rect 650164 909470 654935 909472
rect 654869 909467 654935 909470
rect 58433 897834 58499 897837
rect 58433 897832 64492 897834
rect 58433 897776 58438 897832
rect 58494 897776 64492 897832
rect 58433 897774 64492 897776
rect 58433 897771 58499 897774
rect 654869 896202 654935 896205
rect 650164 896200 654935 896202
rect 650164 896144 654874 896200
rect 654930 896144 654935 896200
rect 650164 896142 654935 896144
rect 654869 896139 654935 896142
rect 58433 884778 58499 884781
rect 58433 884776 64492 884778
rect 58433 884720 58438 884776
rect 58494 884720 64492 884776
rect 58433 884718 64492 884720
rect 58433 884715 58499 884718
rect 655145 882874 655211 882877
rect 650164 882872 655211 882874
rect 650164 882816 655150 882872
rect 655206 882816 655211 882872
rect 650164 882814 655211 882816
rect 655145 882811 655211 882814
rect 675753 877298 675819 877301
rect 676070 877298 676076 877300
rect 675753 877296 676076 877298
rect 675753 877240 675758 877296
rect 675814 877240 676076 877296
rect 675753 877238 676076 877240
rect 675753 877235 675819 877238
rect 676070 877236 676076 877238
rect 676140 877236 676146 877300
rect 675661 876620 675727 876621
rect 675661 876616 675708 876620
rect 675772 876618 675778 876620
rect 675661 876560 675666 876616
rect 675661 876556 675708 876560
rect 675772 876558 675818 876618
rect 675772 876556 675778 876558
rect 675661 876555 675727 876556
rect 675477 875940 675543 875941
rect 675477 875936 675524 875940
rect 675588 875938 675594 875940
rect 675477 875880 675482 875936
rect 675477 875876 675524 875880
rect 675588 875878 675634 875938
rect 675588 875876 675594 875878
rect 675477 875875 675543 875876
rect 675385 874036 675451 874037
rect 675334 874034 675340 874036
rect 675294 873974 675340 874034
rect 675404 874032 675451 874036
rect 675446 873976 675451 874032
rect 675334 873972 675340 873974
rect 675404 873972 675451 873976
rect 675385 873971 675451 873972
rect 675753 872266 675819 872269
rect 675886 872266 675892 872268
rect 675753 872264 675892 872266
rect 675753 872208 675758 872264
rect 675814 872208 675892 872264
rect 675753 872206 675892 872208
rect 675753 872203 675819 872206
rect 675886 872204 675892 872206
rect 675956 872204 675962 872268
rect 58433 871722 58499 871725
rect 58433 871720 64492 871722
rect 58433 871664 58438 871720
rect 58494 871664 64492 871720
rect 58433 871662 64492 871664
rect 58433 871659 58499 871662
rect 656801 869682 656867 869685
rect 650164 869680 656867 869682
rect 650164 869624 656806 869680
rect 656862 869624 656867 869680
rect 650164 869622 656867 869624
rect 656801 869619 656867 869622
rect 58433 858666 58499 858669
rect 58433 858664 64492 858666
rect 58433 858608 58438 858664
rect 58494 858608 64492 858664
rect 58433 858606 64492 858608
rect 58433 858603 58499 858606
rect 654685 856354 654751 856357
rect 650164 856352 654751 856354
rect 650164 856296 654690 856352
rect 654746 856296 654751 856352
rect 650164 856294 654751 856296
rect 654685 856291 654751 856294
rect 58433 845610 58499 845613
rect 58433 845608 64492 845610
rect 58433 845552 58438 845608
rect 58494 845552 64492 845608
rect 58433 845550 64492 845552
rect 58433 845547 58499 845550
rect 655053 843026 655119 843029
rect 650164 843024 655119 843026
rect 650164 842968 655058 843024
rect 655114 842968 655119 843024
rect 650164 842966 655119 842968
rect 655053 842963 655119 842966
rect 57973 832554 58039 832557
rect 57973 832552 64492 832554
rect 57973 832496 57978 832552
rect 58034 832496 64492 832552
rect 57973 832494 64492 832496
rect 57973 832491 58039 832494
rect 655513 829834 655579 829837
rect 650164 829832 655579 829834
rect 650164 829776 655518 829832
rect 655574 829776 655579 829832
rect 650164 829774 655579 829776
rect 655513 829771 655579 829774
rect 59169 819498 59235 819501
rect 59169 819496 64492 819498
rect 59169 819440 59174 819496
rect 59230 819440 64492 819496
rect 59169 819438 64492 819440
rect 59169 819435 59235 819438
rect 41781 817730 41847 817733
rect 41492 817728 41847 817730
rect 41492 817672 41786 817728
rect 41842 817672 41847 817728
rect 41492 817670 41847 817672
rect 41781 817667 41847 817670
rect 41781 817322 41847 817325
rect 41492 817320 41847 817322
rect 41492 817264 41786 817320
rect 41842 817264 41847 817320
rect 41492 817262 41847 817264
rect 41781 817259 41847 817262
rect 53833 816914 53899 816917
rect 41492 816912 53899 816914
rect 41492 816856 53838 816912
rect 53894 816856 53899 816912
rect 41492 816854 53899 816856
rect 53833 816851 53899 816854
rect 41873 816506 41939 816509
rect 654133 816506 654199 816509
rect 41492 816504 41939 816506
rect 41492 816448 41878 816504
rect 41934 816448 41939 816504
rect 41492 816446 41939 816448
rect 650164 816504 654199 816506
rect 650164 816448 654138 816504
rect 654194 816448 654199 816504
rect 650164 816446 654199 816448
rect 41873 816443 41939 816446
rect 654133 816443 654199 816446
rect 42701 816098 42767 816101
rect 41492 816096 42767 816098
rect 41492 816040 42706 816096
rect 42762 816040 42767 816096
rect 41492 816038 42767 816040
rect 42701 816035 42767 816038
rect 41689 815824 41755 815829
rect 41689 815768 41694 815824
rect 41750 815768 41755 815824
rect 41689 815763 41755 815768
rect 41692 815690 41752 815763
rect 41492 815630 41752 815690
rect 43713 815282 43779 815285
rect 41492 815280 43779 815282
rect 41492 815224 43718 815280
rect 43774 815224 43779 815280
rect 41492 815222 43779 815224
rect 43713 815219 43779 815222
rect 42333 814874 42399 814877
rect 41492 814872 42399 814874
rect 41492 814816 42338 814872
rect 42394 814816 42399 814872
rect 41492 814814 42399 814816
rect 42333 814811 42399 814814
rect 41781 814466 41847 814469
rect 41492 814464 41847 814466
rect 41492 814408 41786 814464
rect 41842 814408 41847 814464
rect 41492 814406 41847 814408
rect 41781 814403 41847 814406
rect 41873 814196 41939 814197
rect 41822 814194 41828 814196
rect 41746 814134 41828 814194
rect 41892 814194 41939 814196
rect 62849 814194 62915 814197
rect 41892 814192 62915 814194
rect 41934 814136 62854 814192
rect 62910 814136 62915 814192
rect 41822 814132 41828 814134
rect 41892 814134 62915 814136
rect 41892 814132 41939 814134
rect 41873 814131 41939 814132
rect 62849 814131 62915 814134
rect 43345 814058 43411 814061
rect 41492 814056 43411 814058
rect 41492 814000 43350 814056
rect 43406 814000 43411 814056
rect 41492 813998 43411 814000
rect 43345 813995 43411 813998
rect 41781 813650 41847 813653
rect 41492 813648 41847 813650
rect 41492 813592 41786 813648
rect 41842 813592 41847 813648
rect 41492 813590 41847 813592
rect 41781 813587 41847 813590
rect 42977 813242 43043 813245
rect 41492 813240 43043 813242
rect 41492 813184 42982 813240
rect 43038 813184 43043 813240
rect 41492 813182 43043 813184
rect 42977 813179 43043 813182
rect 42885 812834 42951 812837
rect 41492 812832 42951 812834
rect 41492 812776 42890 812832
rect 42946 812776 42951 812832
rect 41492 812774 42951 812776
rect 42885 812771 42951 812774
rect 43437 812426 43503 812429
rect 41492 812424 43503 812426
rect 41492 812368 43442 812424
rect 43498 812368 43503 812424
rect 41492 812366 43503 812368
rect 43437 812363 43503 812366
rect 43529 812018 43595 812021
rect 41492 812016 43595 812018
rect 41492 811960 43534 812016
rect 43590 811960 43595 812016
rect 41492 811958 43595 811960
rect 43529 811955 43595 811958
rect 41781 811610 41847 811613
rect 41492 811608 41847 811610
rect 41492 811552 41786 811608
rect 41842 811552 41847 811608
rect 41492 811550 41847 811552
rect 41781 811547 41847 811550
rect 41873 811202 41939 811205
rect 41492 811200 41939 811202
rect 41492 811144 41878 811200
rect 41934 811144 41939 811200
rect 41492 811142 41939 811144
rect 41873 811139 41939 811142
rect 43897 810794 43963 810797
rect 41492 810792 43963 810794
rect 41492 810736 43902 810792
rect 43958 810736 43963 810792
rect 41492 810734 43963 810736
rect 43897 810731 43963 810734
rect 43161 810386 43227 810389
rect 41492 810384 43227 810386
rect 41492 810328 43166 810384
rect 43222 810328 43227 810384
rect 41492 810326 43227 810328
rect 43161 810323 43227 810326
rect 43989 809978 44055 809981
rect 41492 809976 44055 809978
rect 41492 809920 43994 809976
rect 44050 809920 44055 809976
rect 41492 809918 44055 809920
rect 43989 809915 44055 809918
rect 43069 809570 43135 809573
rect 41492 809568 43135 809570
rect 41492 809512 43074 809568
rect 43130 809512 43135 809568
rect 41492 809510 43135 809512
rect 43069 809507 43135 809510
rect 43253 809162 43319 809165
rect 41492 809160 43319 809162
rect 41492 809104 43258 809160
rect 43314 809104 43319 809160
rect 41492 809102 43319 809104
rect 43253 809099 43319 809102
rect 43621 808754 43687 808757
rect 41492 808752 43687 808754
rect 41492 808696 43626 808752
rect 43682 808696 43687 808752
rect 41492 808694 43687 808696
rect 43621 808691 43687 808694
rect 41781 808346 41847 808349
rect 41492 808344 41847 808346
rect 41492 808288 41786 808344
rect 41842 808288 41847 808344
rect 41492 808286 41847 808288
rect 41781 808283 41847 808286
rect 41781 807938 41847 807941
rect 41492 807936 41847 807938
rect 41492 807880 41786 807936
rect 41842 807880 41847 807936
rect 41492 807878 41847 807880
rect 41781 807875 41847 807878
rect 41965 807530 42031 807533
rect 41492 807528 42031 807530
rect 41492 807472 41970 807528
rect 42026 807472 42031 807528
rect 41492 807470 42031 807472
rect 41965 807467 42031 807470
rect 30422 806684 30482 807092
rect 58433 806578 58499 806581
rect 58433 806576 64492 806578
rect 58433 806520 58438 806576
rect 58494 806520 64492 806576
rect 58433 806518 64492 806520
rect 58433 806515 58499 806518
rect 41965 806306 42031 806309
rect 41492 806304 42031 806306
rect 41492 806248 41970 806304
rect 42026 806248 42031 806304
rect 41492 806246 42031 806248
rect 41965 806243 42031 806246
rect 656801 803314 656867 803317
rect 650164 803312 656867 803314
rect 650164 803256 656806 803312
rect 656862 803256 656867 803312
rect 650164 803254 656867 803256
rect 656801 803251 656867 803254
rect 674281 797738 674347 797741
rect 676254 797738 676260 797740
rect 674281 797736 676260 797738
rect 674281 797680 674286 797736
rect 674342 797680 676260 797736
rect 674281 797678 676260 797680
rect 674281 797675 674347 797678
rect 676254 797676 676260 797678
rect 676324 797676 676330 797740
rect 58065 793522 58131 793525
rect 58065 793520 64492 793522
rect 58065 793464 58070 793520
rect 58126 793464 64492 793520
rect 58065 793462 64492 793464
rect 58065 793459 58131 793462
rect 674189 792026 674255 792029
rect 676438 792026 676444 792028
rect 674189 792024 676444 792026
rect 674189 791968 674194 792024
rect 674250 791968 676444 792024
rect 674189 791966 676444 791968
rect 674189 791963 674255 791966
rect 676438 791964 676444 791966
rect 676508 791964 676514 792028
rect 655053 789986 655119 789989
rect 650164 789984 655119 789986
rect 650164 789928 655058 789984
rect 655114 789928 655119 789984
rect 650164 789926 655119 789928
rect 655053 789923 655119 789926
rect 674966 787748 674972 787812
rect 675036 787810 675042 787812
rect 675385 787810 675451 787813
rect 675036 787808 675451 787810
rect 675036 787752 675390 787808
rect 675446 787752 675451 787808
rect 675036 787750 675451 787752
rect 675036 787748 675042 787750
rect 675385 787747 675451 787750
rect 674598 787204 674604 787268
rect 674668 787266 674674 787268
rect 675385 787266 675451 787269
rect 674668 787264 675451 787266
rect 674668 787208 675390 787264
rect 675446 787208 675451 787264
rect 674668 787206 675451 787208
rect 674668 787204 674674 787206
rect 675385 787203 675451 787206
rect 674414 786796 674420 786860
rect 674484 786858 674490 786860
rect 675385 786858 675451 786861
rect 674484 786856 675451 786858
rect 674484 786800 675390 786856
rect 675446 786800 675451 786856
rect 674484 786798 675451 786800
rect 674484 786796 674490 786798
rect 675385 786795 675451 786798
rect 675150 784076 675156 784140
rect 675220 784138 675226 784140
rect 675385 784138 675451 784141
rect 675220 784136 675451 784138
rect 675220 784080 675390 784136
rect 675446 784080 675451 784136
rect 675220 784078 675451 784080
rect 675220 784076 675226 784078
rect 675385 784075 675451 784078
rect 674782 783804 674788 783868
rect 674852 783866 674858 783868
rect 675477 783866 675543 783869
rect 674852 783864 675543 783866
rect 674852 783808 675482 783864
rect 675538 783808 675543 783864
rect 674852 783806 675543 783808
rect 674852 783804 674858 783806
rect 675477 783803 675543 783806
rect 58433 780466 58499 780469
rect 58433 780464 64492 780466
rect 58433 780408 58438 780464
rect 58494 780408 64492 780464
rect 58433 780406 64492 780408
rect 58433 780403 58499 780406
rect 674230 777412 674236 777476
rect 674300 777474 674306 777476
rect 674373 777474 674439 777477
rect 674300 777472 674439 777474
rect 674300 777416 674378 777472
rect 674434 777416 674439 777472
rect 674300 777414 674439 777416
rect 674300 777412 674306 777414
rect 674373 777411 674439 777414
rect 655513 776658 655579 776661
rect 650164 776656 655579 776658
rect 650164 776600 655518 776656
rect 655574 776600 655579 776656
rect 650164 776598 655579 776600
rect 655513 776595 655579 776598
rect 41505 774754 41571 774757
rect 41462 774752 41571 774754
rect 41462 774696 41510 774752
rect 41566 774696 41571 774752
rect 41462 774691 41571 774696
rect 41462 774452 41522 774691
rect 41505 774346 41571 774349
rect 41462 774344 41571 774346
rect 41462 774288 41510 774344
rect 41566 774288 41571 774344
rect 41462 774283 41571 774288
rect 41462 774044 41522 774283
rect 41505 773938 41571 773941
rect 41462 773936 41571 773938
rect 41462 773880 41510 773936
rect 41566 773880 41571 773936
rect 41462 773875 41571 773880
rect 41462 773636 41522 773875
rect 674230 773332 674236 773396
rect 674300 773394 674306 773396
rect 675753 773394 675819 773397
rect 674300 773392 675819 773394
rect 674300 773336 675758 773392
rect 675814 773336 675819 773392
rect 674300 773334 675819 773336
rect 674300 773332 674306 773334
rect 675753 773331 675819 773334
rect 42057 773258 42123 773261
rect 41492 773256 42123 773258
rect 41492 773200 42062 773256
rect 42118 773200 42123 773256
rect 41492 773198 42123 773200
rect 42057 773195 42123 773198
rect 39982 773060 39988 773124
rect 40052 773060 40058 773124
rect 39990 772820 40050 773060
rect 676806 772652 676812 772716
rect 676876 772714 676882 772716
rect 679065 772714 679131 772717
rect 676876 772712 679131 772714
rect 676876 772656 679070 772712
rect 679126 772656 679131 772712
rect 676876 772654 679131 772656
rect 676876 772652 676882 772654
rect 679065 772651 679131 772654
rect 43345 772442 43411 772445
rect 41492 772440 43411 772442
rect 41492 772384 43350 772440
rect 43406 772384 43411 772440
rect 41492 772382 43411 772384
rect 43345 772379 43411 772382
rect 42149 772034 42215 772037
rect 41492 772032 42215 772034
rect 41492 771976 42154 772032
rect 42210 771976 42215 772032
rect 41492 771974 42215 771976
rect 42149 771971 42215 771974
rect 39990 771492 40050 771596
rect 39982 771428 39988 771492
rect 40052 771428 40058 771492
rect 43713 771218 43779 771221
rect 41492 771216 43779 771218
rect 41492 771188 43718 771216
rect 41462 771160 43718 771188
rect 43774 771160 43779 771216
rect 41462 771158 43779 771160
rect 41462 771084 41522 771158
rect 43713 771155 43779 771158
rect 41454 771020 41460 771084
rect 41524 771020 41530 771084
rect 44081 770810 44147 770813
rect 41492 770808 44147 770810
rect 41492 770752 44086 770808
rect 44142 770752 44147 770808
rect 41492 770750 44147 770752
rect 44081 770747 44147 770750
rect 42885 770402 42951 770405
rect 41492 770400 42951 770402
rect 41492 770344 42890 770400
rect 42946 770344 42951 770400
rect 41492 770342 42951 770344
rect 42885 770339 42951 770342
rect 43989 769994 44055 769997
rect 41492 769992 44055 769994
rect 41492 769936 43994 769992
rect 44050 769936 44055 769992
rect 41492 769934 44055 769936
rect 43989 769931 44055 769934
rect 42425 769586 42491 769589
rect 41492 769584 42491 769586
rect 41492 769528 42430 769584
rect 42486 769528 42491 769584
rect 41492 769526 42491 769528
rect 42425 769523 42491 769526
rect 43253 769178 43319 769181
rect 41492 769176 43319 769178
rect 41492 769120 43258 769176
rect 43314 769120 43319 769176
rect 41492 769118 43319 769120
rect 43253 769115 43319 769118
rect 43437 768770 43503 768773
rect 41492 768768 43503 768770
rect 41492 768712 43442 768768
rect 43498 768712 43503 768768
rect 41492 768710 43503 768712
rect 43437 768707 43503 768710
rect 43161 768362 43227 768365
rect 41492 768360 43227 768362
rect 41492 768304 43166 768360
rect 43222 768304 43227 768360
rect 41492 768302 43227 768304
rect 43161 768299 43227 768302
rect 41873 767954 41939 767957
rect 41492 767952 41939 767954
rect 41492 767896 41878 767952
rect 41934 767896 41939 767952
rect 41492 767894 41939 767896
rect 41873 767891 41939 767894
rect 43621 767546 43687 767549
rect 41492 767544 43687 767546
rect 41492 767488 43626 767544
rect 43682 767488 43687 767544
rect 41492 767486 43687 767488
rect 43621 767483 43687 767486
rect 58433 767410 58499 767413
rect 58433 767408 64492 767410
rect 58433 767352 58438 767408
rect 58494 767352 64492 767408
rect 58433 767350 64492 767352
rect 58433 767347 58499 767350
rect 42701 767138 42767 767141
rect 41492 767136 42767 767138
rect 41492 767080 42706 767136
rect 42762 767080 42767 767136
rect 41492 767078 42767 767080
rect 42701 767075 42767 767078
rect 41965 766730 42031 766733
rect 41492 766728 42031 766730
rect 41492 766672 41970 766728
rect 42026 766672 42031 766728
rect 41492 766670 42031 766672
rect 41965 766667 42031 766670
rect 43069 766322 43135 766325
rect 41492 766320 43135 766322
rect 41492 766264 43074 766320
rect 43130 766264 43135 766320
rect 41492 766262 43135 766264
rect 43069 766259 43135 766262
rect 43253 765914 43319 765917
rect 41492 765912 43319 765914
rect 41492 765856 43258 765912
rect 43314 765856 43319 765912
rect 41492 765854 43319 765856
rect 43253 765851 43319 765854
rect 43713 765506 43779 765509
rect 41492 765504 43779 765506
rect 41492 765448 43718 765504
rect 43774 765448 43779 765504
rect 41492 765446 43779 765448
rect 43713 765443 43779 765446
rect 43161 765098 43227 765101
rect 41492 765096 43227 765098
rect 41492 765040 43166 765096
rect 43222 765040 43227 765096
rect 41492 765038 43227 765040
rect 43161 765035 43227 765038
rect 42885 764690 42951 764693
rect 41492 764688 42951 764690
rect 41492 764632 42890 764688
rect 42946 764632 42951 764688
rect 41492 764630 42951 764632
rect 42885 764627 42951 764630
rect 41462 764149 41522 764252
rect 41462 764144 41571 764149
rect 41462 764088 41510 764144
rect 41566 764088 41571 764144
rect 41462 764086 41571 764088
rect 41505 764083 41571 764086
rect 30422 763436 30482 763844
rect 654777 763330 654843 763333
rect 650164 763328 654843 763330
rect 650164 763272 654782 763328
rect 654838 763272 654843 763328
rect 650164 763270 654843 763272
rect 654777 763267 654843 763270
rect 41462 762925 41522 763028
rect 41462 762920 41571 762925
rect 41462 762864 41510 762920
rect 41566 762864 41571 762920
rect 41462 762862 41571 762864
rect 41505 762859 41571 762862
rect 679022 761293 679082 761532
rect 678973 761288 679082 761293
rect 678973 761232 678978 761288
rect 679034 761232 679082 761288
rect 678973 761230 679082 761232
rect 678973 761227 679039 761230
rect 676262 760885 676322 761124
rect 676213 760880 676322 760885
rect 676213 760824 676218 760880
rect 676274 760824 676322 760880
rect 676213 760822 676322 760824
rect 676213 760819 676279 760822
rect 676121 760474 676187 760477
rect 676262 760474 676322 760716
rect 676121 760472 676322 760474
rect 676121 760416 676126 760472
rect 676182 760416 676322 760472
rect 676121 760414 676322 760416
rect 676121 760411 676187 760414
rect 673545 760338 673611 760341
rect 673862 760338 673868 760340
rect 673545 760336 673868 760338
rect 673545 760280 673550 760336
rect 673606 760280 673868 760336
rect 673545 760278 673868 760280
rect 673545 760275 673611 760278
rect 673862 760276 673868 760278
rect 673932 760338 673938 760340
rect 673932 760278 676292 760338
rect 673932 760276 673938 760278
rect 676262 759661 676322 759900
rect 676262 759656 676371 759661
rect 679065 759658 679131 759661
rect 676262 759600 676310 759656
rect 676366 759600 676371 759656
rect 676262 759598 676371 759600
rect 676305 759595 676371 759598
rect 679022 759656 679131 759658
rect 679022 759600 679070 759656
rect 679126 759600 679131 759656
rect 679022 759595 679131 759600
rect 679022 759492 679082 759595
rect 669773 759114 669839 759117
rect 673545 759114 673611 759117
rect 669773 759112 673611 759114
rect 669773 759056 669778 759112
rect 669834 759056 673550 759112
rect 673606 759056 673611 759112
rect 669773 759054 673611 759056
rect 669773 759051 669839 759054
rect 673545 759051 673611 759054
rect 676029 759114 676095 759117
rect 676029 759112 676292 759114
rect 676029 759056 676034 759112
rect 676090 759056 676292 759112
rect 676029 759054 676292 759056
rect 676029 759051 676095 759054
rect 679022 758437 679082 758676
rect 678973 758432 679082 758437
rect 678973 758376 678978 758432
rect 679034 758376 679082 758432
rect 678973 758374 679082 758376
rect 678973 758371 679039 758374
rect 676262 758029 676322 758268
rect 676262 758024 676371 758029
rect 676262 757968 676310 758024
rect 676366 757968 676371 758024
rect 676262 757966 676371 757968
rect 676305 757963 676371 757966
rect 43294 757692 43300 757756
rect 43364 757754 43370 757756
rect 43621 757754 43687 757757
rect 43364 757752 43687 757754
rect 43364 757696 43626 757752
rect 43682 757696 43687 757752
rect 43364 757694 43687 757696
rect 43364 757692 43370 757694
rect 43621 757691 43687 757694
rect 676121 757618 676187 757621
rect 676262 757618 676322 757860
rect 676121 757616 676322 757618
rect 676121 757560 676126 757616
rect 676182 757560 676322 757616
rect 676121 757558 676322 757560
rect 676121 757555 676187 757558
rect 676262 757213 676322 757452
rect 676213 757208 676322 757213
rect 676213 757152 676218 757208
rect 676274 757152 676322 757208
rect 676213 757150 676322 757152
rect 676213 757147 676279 757150
rect 41781 757076 41847 757077
rect 41781 757074 41828 757076
rect 41736 757072 41828 757074
rect 41736 757016 41786 757072
rect 41736 757014 41828 757016
rect 41781 757012 41828 757014
rect 41892 757012 41898 757076
rect 41965 757074 42031 757077
rect 42190 757074 42196 757076
rect 41965 757072 42196 757074
rect 41965 757016 41970 757072
rect 42026 757016 42196 757072
rect 41965 757014 42196 757016
rect 41781 757011 41847 757012
rect 41965 757011 42031 757014
rect 42190 757012 42196 757014
rect 42260 757012 42266 757076
rect 675518 757012 675524 757076
rect 675588 757074 675594 757076
rect 675588 757014 676292 757074
rect 675588 757012 675594 757014
rect 676029 756666 676095 756669
rect 676029 756664 676292 756666
rect 676029 756608 676034 756664
rect 676090 756608 676292 756664
rect 676029 756606 676292 756608
rect 676029 756603 676095 756606
rect 676070 756332 676076 756396
rect 676140 756394 676146 756396
rect 676140 756334 676322 756394
rect 676140 756332 676146 756334
rect 676262 756228 676322 756334
rect 675334 755788 675340 755852
rect 675404 755850 675410 755852
rect 675404 755790 676292 755850
rect 675404 755788 675410 755790
rect 676121 755578 676187 755581
rect 676121 755576 676322 755578
rect 676121 755520 676126 755576
rect 676182 755520 676322 755576
rect 676121 755518 676322 755520
rect 676121 755515 676187 755518
rect 676262 755412 676322 755518
rect 42190 755244 42196 755308
rect 42260 755306 42266 755308
rect 42609 755306 42675 755309
rect 42260 755304 42675 755306
rect 42260 755248 42614 755304
rect 42670 755248 42675 755304
rect 42260 755246 42675 755248
rect 42260 755244 42266 755246
rect 42609 755243 42675 755246
rect 676029 755034 676095 755037
rect 676029 755032 676292 755034
rect 676029 754976 676034 755032
rect 676090 754976 676292 755032
rect 676029 754974 676292 754976
rect 676029 754971 676095 754974
rect 675702 754564 675708 754628
rect 675772 754626 675778 754628
rect 675772 754566 676292 754626
rect 675772 754564 675778 754566
rect 58341 754354 58407 754357
rect 58341 754352 64492 754354
rect 58341 754296 58346 754352
rect 58402 754296 64492 754352
rect 58341 754294 64492 754296
rect 58341 754291 58407 754294
rect 675569 754218 675635 754221
rect 675569 754216 676292 754218
rect 675569 754160 675574 754216
rect 675630 754160 676292 754216
rect 675569 754158 676292 754160
rect 675569 754155 675635 754158
rect 41873 754084 41939 754085
rect 41822 754020 41828 754084
rect 41892 754082 41939 754084
rect 41892 754080 41984 754082
rect 41934 754024 41984 754080
rect 41892 754022 41984 754024
rect 41892 754020 41939 754022
rect 41873 754019 41939 754020
rect 675753 753810 675819 753813
rect 675753 753808 676292 753810
rect 675753 753752 675758 753808
rect 675814 753752 676292 753808
rect 675753 753750 676292 753752
rect 675753 753747 675819 753750
rect 676029 753402 676095 753405
rect 676029 753400 676292 753402
rect 676029 753344 676034 753400
rect 676090 753344 676292 753400
rect 676029 753342 676292 753344
rect 676029 753339 676095 753342
rect 43069 752994 43135 752997
rect 43294 752994 43300 752996
rect 43069 752992 43300 752994
rect 43069 752936 43074 752992
rect 43130 752936 43300 752992
rect 43069 752934 43300 752936
rect 43069 752931 43135 752934
rect 43294 752932 43300 752934
rect 43364 752932 43370 752996
rect 676029 752994 676095 752997
rect 676029 752992 676292 752994
rect 676029 752936 676034 752992
rect 676090 752936 676292 752992
rect 676029 752934 676292 752936
rect 676029 752931 676095 752934
rect 675886 752524 675892 752588
rect 675956 752586 675962 752588
rect 675956 752526 676292 752586
rect 675956 752524 675962 752526
rect 676438 752252 676444 752316
rect 676508 752252 676514 752316
rect 676446 752148 676506 752252
rect 676254 751844 676260 751908
rect 676324 751844 676330 751908
rect 676262 751740 676322 751844
rect 679022 751093 679082 751332
rect 678973 751088 679082 751093
rect 678973 751032 678978 751088
rect 679034 751032 679082 751088
rect 678973 751030 679082 751032
rect 678973 751027 679039 751030
rect 679022 750516 679082 750924
rect 678973 750274 679039 750277
rect 678973 750272 679082 750274
rect 678973 750216 678978 750272
rect 679034 750216 679082 750272
rect 678973 750211 679082 750216
rect 654869 750138 654935 750141
rect 650164 750136 654935 750138
rect 650164 750080 654874 750136
rect 654930 750080 654935 750136
rect 679022 750108 679082 750211
rect 650164 750078 654935 750080
rect 654869 750075 654935 750078
rect 675477 744154 675543 744157
rect 676622 744154 676628 744156
rect 675477 744152 676628 744154
rect 675477 744096 675482 744152
rect 675538 744096 676628 744152
rect 675477 744094 676628 744096
rect 675477 744091 675543 744094
rect 676622 744092 676628 744094
rect 676692 744092 676698 744156
rect 675661 744018 675727 744021
rect 676254 744018 676260 744020
rect 675661 744016 676260 744018
rect 675661 743960 675666 744016
rect 675722 743960 676260 744016
rect 675661 743958 676260 743960
rect 675661 743955 675727 743958
rect 676254 743956 676260 743958
rect 676324 743956 676330 744020
rect 675753 742930 675819 742933
rect 675886 742930 675892 742932
rect 675753 742928 675892 742930
rect 675753 742872 675758 742928
rect 675814 742872 675892 742928
rect 675753 742870 675892 742872
rect 675753 742867 675819 742870
rect 675886 742868 675892 742870
rect 675956 742868 675962 742932
rect 675753 742522 675819 742525
rect 676070 742522 676076 742524
rect 675753 742520 676076 742522
rect 675753 742464 675758 742520
rect 675814 742464 676076 742520
rect 675753 742462 676076 742464
rect 675753 742459 675819 742462
rect 676070 742460 676076 742462
rect 676140 742460 676146 742524
rect 674046 741644 674052 741708
rect 674116 741706 674122 741708
rect 675477 741706 675543 741709
rect 674116 741704 675543 741706
rect 674116 741648 675482 741704
rect 675538 741648 675543 741704
rect 674116 741646 675543 741648
rect 674116 741644 674122 741646
rect 675477 741643 675543 741646
rect 58433 741298 58499 741301
rect 58433 741296 64492 741298
rect 58433 741240 58438 741296
rect 58494 741240 64492 741296
rect 58433 741238 64492 741240
rect 58433 741235 58499 741238
rect 673862 739740 673868 739804
rect 673932 739802 673938 739804
rect 675385 739802 675451 739805
rect 673932 739800 675451 739802
rect 673932 739744 675390 739800
rect 675446 739744 675451 739800
rect 673932 739742 675451 739744
rect 673932 739740 673938 739742
rect 675385 739739 675451 739742
rect 673678 739060 673684 739124
rect 673748 739122 673754 739124
rect 675385 739122 675451 739125
rect 673748 739120 675451 739122
rect 673748 739064 675390 739120
rect 675446 739064 675451 739120
rect 673748 739062 675451 739064
rect 673748 739060 673754 739062
rect 675385 739059 675451 739062
rect 675661 738580 675727 738581
rect 675661 738576 675708 738580
rect 675772 738578 675778 738580
rect 675661 738520 675666 738576
rect 675661 738516 675708 738520
rect 675772 738518 675818 738578
rect 675772 738516 675778 738518
rect 675661 738515 675727 738516
rect 675753 738034 675819 738037
rect 676438 738034 676444 738036
rect 675753 738032 676444 738034
rect 675753 737976 675758 738032
rect 675814 737976 676444 738032
rect 675753 737974 676444 737976
rect 675753 737971 675819 737974
rect 676438 737972 676444 737974
rect 676508 737972 676514 738036
rect 654777 736810 654843 736813
rect 650164 736808 654843 736810
rect 650164 736752 654782 736808
rect 654838 736752 654843 736808
rect 650164 736750 654843 736752
rect 654777 736747 654843 736750
rect 51257 731370 51323 731373
rect 41492 731368 51323 731370
rect 41492 731312 51262 731368
rect 51318 731312 51323 731368
rect 41492 731310 51323 731312
rect 51257 731307 51323 731310
rect 39757 731098 39823 731101
rect 39982 731098 39988 731100
rect 39757 731096 39988 731098
rect 39757 731040 39762 731096
rect 39818 731040 39988 731096
rect 39757 731038 39988 731040
rect 39757 731035 39823 731038
rect 39982 731036 39988 731038
rect 40052 731036 40058 731100
rect 48589 730962 48655 730965
rect 41492 730960 48655 730962
rect 41492 730904 48594 730960
rect 48650 730904 48655 730960
rect 41492 730902 48655 730904
rect 48589 730899 48655 730902
rect 51073 730554 51139 730557
rect 41492 730552 51139 730554
rect 41492 730496 51078 730552
rect 51134 730496 51139 730552
rect 41492 730494 51139 730496
rect 51073 730491 51139 730494
rect 39757 730282 39823 730285
rect 63033 730282 63099 730285
rect 39757 730280 63099 730282
rect 39757 730224 39762 730280
rect 39818 730224 63038 730280
rect 63094 730224 63099 730280
rect 39757 730222 63099 730224
rect 39757 730219 39823 730222
rect 63033 730219 63099 730222
rect 42793 730146 42859 730149
rect 44173 730146 44239 730149
rect 41492 730144 44239 730146
rect 41492 730088 42798 730144
rect 42854 730088 44178 730144
rect 44234 730088 44239 730144
rect 41492 730086 44239 730088
rect 42793 730083 42859 730086
rect 44173 730083 44239 730086
rect 42977 729738 43043 729741
rect 41492 729736 43043 729738
rect 41492 729680 42982 729736
rect 43038 729680 43043 729736
rect 41492 729678 43043 729680
rect 42977 729675 43043 729678
rect 41505 729466 41571 729469
rect 41462 729464 41571 729466
rect 41462 729408 41510 729464
rect 41566 729408 41571 729464
rect 41462 729403 41571 729408
rect 41462 729300 41522 729403
rect 41781 728922 41847 728925
rect 41492 728920 41847 728922
rect 41492 728864 41786 728920
rect 41842 728864 41847 728920
rect 41492 728862 41847 728864
rect 41781 728859 41847 728862
rect 43621 728514 43687 728517
rect 41492 728512 43687 728514
rect 41492 728456 43626 728512
rect 43682 728456 43687 728512
rect 41492 728454 43687 728456
rect 43621 728451 43687 728454
rect 39757 728242 39823 728245
rect 58433 728242 58499 728245
rect 39757 728240 39866 728242
rect 39757 728184 39762 728240
rect 39818 728184 39866 728240
rect 39757 728179 39866 728184
rect 58433 728240 64492 728242
rect 58433 728184 58438 728240
rect 58494 728184 64492 728240
rect 58433 728182 64492 728184
rect 58433 728179 58499 728182
rect 39806 728076 39866 728179
rect 44265 727698 44331 727701
rect 41492 727696 44331 727698
rect 41492 727640 44270 727696
rect 44326 727640 44331 727696
rect 41492 727638 44331 727640
rect 44265 727635 44331 727638
rect 42517 727290 42583 727293
rect 41492 727288 42583 727290
rect 41492 727232 42522 727288
rect 42578 727232 42583 727288
rect 41492 727230 42583 727232
rect 42517 727227 42583 727230
rect 43529 726882 43595 726885
rect 41492 726880 43595 726882
rect 41492 726824 43534 726880
rect 43590 726824 43595 726880
rect 41492 726822 43595 726824
rect 43529 726819 43595 726822
rect 42885 726474 42951 726477
rect 41492 726472 42951 726474
rect 41492 726416 42890 726472
rect 42946 726416 42951 726472
rect 41492 726414 42951 726416
rect 42885 726411 42951 726414
rect 43253 726066 43319 726069
rect 41492 726064 43319 726066
rect 41492 726008 43258 726064
rect 43314 726008 43319 726064
rect 41492 726006 43319 726008
rect 43253 726003 43319 726006
rect 43437 725658 43503 725661
rect 41492 725656 43503 725658
rect 41492 725600 43442 725656
rect 43498 725600 43503 725656
rect 41492 725598 43503 725600
rect 43437 725595 43503 725598
rect 43345 725250 43411 725253
rect 41492 725248 43411 725250
rect 41492 725192 43350 725248
rect 43406 725192 43411 725248
rect 41492 725190 43411 725192
rect 43345 725187 43411 725190
rect 41873 724842 41939 724845
rect 41492 724840 41939 724842
rect 41492 724784 41878 724840
rect 41934 724784 41939 724840
rect 41492 724782 41939 724784
rect 41873 724779 41939 724782
rect 42977 724434 43043 724437
rect 41492 724432 43043 724434
rect 41492 724376 42982 724432
rect 43038 724376 43043 724432
rect 41492 724374 43043 724376
rect 42977 724371 43043 724374
rect 41278 723757 41338 723996
rect 41278 723752 41387 723757
rect 41278 723696 41326 723752
rect 41382 723696 41387 723752
rect 41278 723694 41387 723696
rect 41321 723691 41387 723694
rect 43069 723618 43135 723621
rect 41492 723616 43135 723618
rect 41492 723560 43074 723616
rect 43130 723560 43135 723616
rect 41492 723558 43135 723560
rect 43069 723555 43135 723558
rect 655513 723482 655579 723485
rect 650164 723480 655579 723482
rect 650164 723424 655518 723480
rect 655574 723424 655579 723480
rect 650164 723422 655579 723424
rect 655513 723419 655579 723422
rect 42793 723210 42859 723213
rect 41492 723208 42859 723210
rect 41492 723152 42798 723208
rect 42854 723152 42859 723208
rect 41492 723150 42859 723152
rect 42793 723147 42859 723150
rect 43897 722802 43963 722805
rect 41492 722800 43963 722802
rect 41492 722744 43902 722800
rect 43958 722744 43963 722800
rect 41492 722742 43963 722744
rect 43897 722739 43963 722742
rect 43989 722394 44055 722397
rect 41492 722392 44055 722394
rect 41492 722336 43994 722392
rect 44050 722336 44055 722392
rect 41492 722334 44055 722336
rect 43989 722331 44055 722334
rect 43805 721986 43871 721989
rect 41492 721984 43871 721986
rect 41492 721928 43810 721984
rect 43866 721928 43871 721984
rect 41492 721926 43871 721928
rect 43805 721923 43871 721926
rect 43161 721578 43227 721581
rect 41492 721576 43227 721578
rect 41492 721520 43166 721576
rect 43222 721520 43227 721576
rect 41492 721518 43227 721520
rect 43161 721515 43227 721518
rect 41462 720901 41522 721140
rect 41462 720896 41571 720901
rect 41462 720840 41510 720896
rect 41566 720840 41571 720896
rect 41462 720838 41571 720840
rect 41505 720835 41571 720838
rect 24902 720324 24962 720732
rect 41462 719677 41522 719916
rect 41462 719672 41571 719677
rect 41462 719616 41510 719672
rect 41566 719616 41571 719672
rect 41462 719614 41571 719616
rect 41505 719611 41571 719614
rect 676029 716546 676095 716549
rect 676029 716544 676292 716546
rect 676029 716488 676034 716544
rect 676090 716488 676292 716544
rect 676029 716486 676292 716488
rect 676029 716483 676095 716486
rect 675937 716138 676003 716141
rect 675937 716136 676292 716138
rect 675937 716080 675942 716136
rect 675998 716080 676292 716136
rect 675937 716078 676292 716080
rect 675937 716075 676003 716078
rect 675937 715730 676003 715733
rect 675937 715728 676292 715730
rect 675937 715672 675942 715728
rect 675998 715672 676292 715728
rect 675937 715670 676292 715672
rect 675937 715667 676003 715670
rect 58433 715322 58499 715325
rect 675937 715322 676003 715325
rect 58433 715320 64492 715322
rect 58433 715264 58438 715320
rect 58494 715264 64492 715320
rect 58433 715262 64492 715264
rect 675937 715320 676292 715322
rect 675937 715264 675942 715320
rect 675998 715264 676292 715320
rect 675937 715262 676292 715264
rect 58433 715259 58499 715262
rect 675937 715259 676003 715262
rect 676029 714914 676095 714917
rect 676029 714912 676292 714914
rect 676029 714856 676034 714912
rect 676090 714856 676292 714912
rect 676029 714854 676292 714856
rect 676029 714851 676095 714854
rect 678973 714506 679039 714509
rect 678973 714504 679052 714506
rect 678973 714448 678978 714504
rect 679034 714448 679052 714504
rect 678973 714446 679052 714448
rect 678973 714443 679039 714446
rect 676029 714098 676095 714101
rect 676029 714096 676292 714098
rect 676029 714040 676034 714096
rect 676090 714040 676292 714096
rect 676029 714038 676292 714040
rect 676029 714035 676095 714038
rect 676029 713690 676095 713693
rect 676029 713688 676292 713690
rect 676029 713632 676034 713688
rect 676090 713632 676292 713688
rect 676029 713630 676292 713632
rect 676029 713627 676095 713630
rect 676029 713282 676095 713285
rect 676029 713280 676292 713282
rect 676029 713224 676034 713280
rect 676090 713224 676292 713280
rect 676029 713222 676292 713224
rect 676029 713219 676095 713222
rect 676029 712874 676095 712877
rect 676029 712872 676292 712874
rect 676029 712816 676034 712872
rect 676090 712816 676292 712872
rect 676029 712814 676292 712816
rect 676029 712811 676095 712814
rect 676029 712466 676095 712469
rect 676029 712464 676292 712466
rect 676029 712408 676034 712464
rect 676090 712408 676292 712464
rect 676029 712406 676292 712408
rect 676029 712403 676095 712406
rect 674414 711996 674420 712060
rect 674484 712058 674490 712060
rect 674484 711998 676292 712058
rect 674484 711996 674490 711998
rect 676305 711890 676371 711891
rect 676254 711888 676260 711890
rect 676214 711828 676260 711888
rect 676324 711886 676371 711890
rect 676366 711830 676371 711886
rect 676254 711826 676260 711828
rect 676324 711826 676371 711830
rect 676305 711825 676371 711826
rect 676949 711890 677015 711891
rect 676949 711886 676996 711890
rect 677060 711888 677066 711890
rect 676949 711830 676954 711886
rect 676949 711826 676996 711830
rect 677060 711828 677106 711888
rect 677060 711826 677066 711828
rect 676949 711825 677015 711826
rect 675753 711650 675819 711653
rect 675753 711648 676292 711650
rect 675753 711592 675758 711648
rect 675814 711592 676292 711648
rect 675753 711590 676292 711592
rect 675753 711587 675819 711590
rect 674966 711180 674972 711244
rect 675036 711242 675042 711244
rect 675036 711182 676292 711242
rect 675036 711180 675042 711182
rect 675845 710834 675911 710837
rect 675845 710832 676292 710834
rect 675845 710776 675850 710832
rect 675906 710776 676292 710832
rect 675845 710774 676292 710776
rect 675845 710771 675911 710774
rect 675937 710426 676003 710429
rect 675937 710424 676292 710426
rect 675937 710368 675942 710424
rect 675998 710368 676292 710424
rect 675937 710366 676292 710368
rect 675937 710363 676003 710366
rect 655973 710290 656039 710293
rect 650164 710288 656039 710290
rect 650164 710232 655978 710288
rect 656034 710232 656039 710288
rect 650164 710230 656039 710232
rect 655973 710227 656039 710230
rect 676029 710018 676095 710021
rect 676029 710016 676292 710018
rect 676029 709960 676034 710016
rect 676090 709960 676292 710016
rect 676029 709958 676292 709960
rect 676029 709955 676095 709958
rect 674598 709548 674604 709612
rect 674668 709610 674674 709612
rect 674668 709550 676292 709610
rect 674668 709548 674674 709550
rect 675150 709140 675156 709204
rect 675220 709202 675226 709204
rect 675220 709142 676292 709202
rect 675220 709140 675226 709142
rect 674782 708732 674788 708796
rect 674852 708794 674858 708796
rect 674852 708734 676292 708794
rect 674852 708732 674858 708734
rect 676029 708386 676095 708389
rect 676029 708384 676292 708386
rect 676029 708328 676034 708384
rect 676090 708328 676292 708384
rect 676029 708326 676292 708328
rect 676029 708323 676095 708326
rect 676029 707978 676095 707981
rect 676029 707976 676292 707978
rect 676029 707920 676034 707976
rect 676090 707920 676292 707976
rect 676029 707918 676292 707920
rect 676029 707915 676095 707918
rect 676029 707570 676095 707573
rect 676029 707568 676292 707570
rect 676029 707512 676034 707568
rect 676090 707512 676292 707568
rect 676029 707510 676292 707512
rect 676029 707507 676095 707510
rect 676305 707162 676371 707165
rect 676292 707160 676371 707162
rect 676292 707104 676310 707160
rect 676366 707104 676371 707160
rect 676292 707102 676371 707104
rect 676305 707099 676371 707102
rect 676029 706754 676095 706757
rect 676029 706752 676292 706754
rect 676029 706696 676034 706752
rect 676090 706696 676292 706752
rect 676029 706694 676292 706696
rect 676029 706691 676095 706694
rect 676029 706346 676095 706349
rect 676029 706344 676292 706346
rect 676029 706288 676034 706344
rect 676090 706288 676292 706344
rect 676029 706286 676292 706288
rect 676029 706283 676095 706286
rect 684542 705500 684602 705908
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 58617 702266 58683 702269
rect 58617 702264 64492 702266
rect 58617 702208 58622 702264
rect 58678 702208 64492 702264
rect 58617 702206 64492 702208
rect 58617 702203 58683 702206
rect 673821 699818 673887 699821
rect 676806 699818 676812 699820
rect 673821 699816 676812 699818
rect 673821 699760 673826 699816
rect 673882 699760 676812 699816
rect 673821 699758 676812 699760
rect 673821 699755 673887 699758
rect 676806 699756 676812 699758
rect 676876 699756 676882 699820
rect 674005 699682 674071 699685
rect 676254 699682 676260 699684
rect 674005 699680 676260 699682
rect 674005 699624 674010 699680
rect 674066 699624 676260 699680
rect 674005 699622 676260 699624
rect 674005 699619 674071 699622
rect 676254 699620 676260 699622
rect 676324 699620 676330 699684
rect 673729 699546 673795 699549
rect 676990 699546 676996 699548
rect 673729 699544 676996 699546
rect 673729 699488 673734 699544
rect 673790 699488 676996 699544
rect 673729 699486 676996 699488
rect 673729 699483 673795 699486
rect 676990 699484 676996 699486
rect 677060 699484 677066 699548
rect 675477 698188 675543 698189
rect 675477 698184 675524 698188
rect 675588 698186 675594 698188
rect 675477 698128 675482 698184
rect 675477 698124 675524 698128
rect 675588 698126 675634 698186
rect 675588 698124 675594 698126
rect 675477 698123 675543 698124
rect 675385 697236 675451 697237
rect 675334 697234 675340 697236
rect 675294 697174 675340 697234
rect 675404 697232 675451 697236
rect 675446 697176 675451 697232
rect 675334 697172 675340 697174
rect 675404 697172 675451 697176
rect 675385 697171 675451 697172
rect 654685 696962 654751 696965
rect 650164 696960 654751 696962
rect 650164 696904 654690 696960
rect 654746 696904 654751 696960
rect 650164 696902 654751 696904
rect 654685 696899 654751 696902
rect 674230 696628 674236 696692
rect 674300 696690 674306 696692
rect 675385 696690 675451 696693
rect 674300 696688 675451 696690
rect 674300 696632 675390 696688
rect 675446 696632 675451 696688
rect 674300 696630 675451 696632
rect 674300 696628 674306 696630
rect 675385 696627 675451 696630
rect 674414 694996 674420 695060
rect 674484 695058 674490 695060
rect 675385 695058 675451 695061
rect 674484 695056 675451 695058
rect 674484 695000 675390 695056
rect 675446 695000 675451 695056
rect 674484 694998 675451 695000
rect 674484 694996 674490 694998
rect 675385 694995 675451 694998
rect 674598 694180 674604 694244
rect 674668 694242 674674 694244
rect 675477 694242 675543 694245
rect 674668 694240 675543 694242
rect 674668 694184 675482 694240
rect 675538 694184 675543 694240
rect 674668 694182 675543 694184
rect 674668 694180 674674 694182
rect 675477 694179 675543 694182
rect 673494 693636 673500 693700
rect 673564 693698 673570 693700
rect 675385 693698 675451 693701
rect 673564 693696 675451 693698
rect 673564 693640 675390 693696
rect 675446 693640 675451 693696
rect 673564 693638 675451 693640
rect 673564 693636 673570 693638
rect 675385 693635 675451 693638
rect 675753 693018 675819 693021
rect 677174 693018 677180 693020
rect 675753 693016 677180 693018
rect 675753 692960 675758 693016
rect 675814 692960 677180 693016
rect 675753 692958 677180 692960
rect 675753 692955 675819 692958
rect 677174 692956 677180 692958
rect 677244 692956 677250 693020
rect 675753 690162 675819 690165
rect 676622 690162 676628 690164
rect 675753 690160 676628 690162
rect 675753 690104 675758 690160
rect 675814 690104 676628 690160
rect 675753 690102 676628 690104
rect 675753 690099 675819 690102
rect 676622 690100 676628 690102
rect 676692 690100 676698 690164
rect 58433 689210 58499 689213
rect 58433 689208 64492 689210
rect 58433 689152 58438 689208
rect 58494 689152 64492 689208
rect 58433 689150 64492 689152
rect 58433 689147 58499 689150
rect 41505 688394 41571 688397
rect 41462 688392 41571 688394
rect 41462 688336 41510 688392
rect 41566 688336 41571 688392
rect 41462 688331 41571 688336
rect 41462 688092 41522 688331
rect 41781 687714 41847 687717
rect 41492 687712 41847 687714
rect 41492 687656 41786 687712
rect 41842 687656 41847 687712
rect 41492 687654 41847 687656
rect 41781 687651 41847 687654
rect 41689 687578 41755 687581
rect 41462 687576 41755 687578
rect 41462 687520 41694 687576
rect 41750 687520 41755 687576
rect 41462 687518 41755 687520
rect 41462 687276 41522 687518
rect 41689 687515 41755 687518
rect 41278 686764 41338 686868
rect 41270 686700 41276 686764
rect 41340 686700 41346 686764
rect 44173 686490 44239 686493
rect 41492 686488 44239 686490
rect 41492 686432 44178 686488
rect 44234 686432 44239 686488
rect 41492 686430 44239 686432
rect 44173 686427 44239 686430
rect 44357 686082 44423 686085
rect 41492 686080 44423 686082
rect 41492 686024 44362 686080
rect 44418 686024 44423 686080
rect 41492 686022 44423 686024
rect 44357 686019 44423 686022
rect 43161 685674 43227 685677
rect 41492 685672 43227 685674
rect 41492 685616 43166 685672
rect 43222 685616 43227 685672
rect 41492 685614 43227 685616
rect 43161 685611 43227 685614
rect 43345 685266 43411 685269
rect 44030 685266 44036 685268
rect 41492 685264 44036 685266
rect 41492 685208 43350 685264
rect 43406 685208 44036 685264
rect 41492 685206 44036 685208
rect 43345 685203 43411 685206
rect 44030 685204 44036 685206
rect 44100 685204 44106 685268
rect 42977 684858 43043 684861
rect 41492 684856 43043 684858
rect 41492 684800 42982 684856
rect 43038 684800 43043 684856
rect 41492 684798 43043 684800
rect 42977 684795 43043 684798
rect 42793 684450 42859 684453
rect 41492 684448 42859 684450
rect 41492 684392 42798 684448
rect 42854 684392 42859 684448
rect 41492 684390 42859 684392
rect 42793 684387 42859 684390
rect 39982 684252 39988 684316
rect 40052 684314 40058 684316
rect 41270 684314 41276 684316
rect 40052 684254 41276 684314
rect 40052 684252 40058 684254
rect 41270 684252 41276 684254
rect 41340 684314 41346 684316
rect 63125 684314 63191 684317
rect 41340 684312 63191 684314
rect 41340 684256 63130 684312
rect 63186 684256 63191 684312
rect 41340 684254 63191 684256
rect 41340 684252 41346 684254
rect 63125 684251 63191 684254
rect 44265 684042 44331 684045
rect 46473 684042 46539 684045
rect 41492 684040 46539 684042
rect 41492 683984 44270 684040
rect 44326 683984 46478 684040
rect 46534 683984 46539 684040
rect 41492 683982 46539 683984
rect 44265 683979 44331 683982
rect 46473 683979 46539 683982
rect 43621 683634 43687 683637
rect 654869 683634 654935 683637
rect 41492 683632 43687 683634
rect 41492 683576 43626 683632
rect 43682 683576 43687 683632
rect 41492 683574 43687 683576
rect 650164 683632 654935 683634
rect 650164 683576 654874 683632
rect 654930 683576 654935 683632
rect 650164 683574 654935 683576
rect 43621 683571 43687 683574
rect 654869 683571 654935 683574
rect 43897 683226 43963 683229
rect 41492 683224 43963 683226
rect 41492 683168 43902 683224
rect 43958 683168 43963 683224
rect 41492 683166 43963 683168
rect 43897 683163 43963 683166
rect 43069 682818 43135 682821
rect 41492 682816 43135 682818
rect 41492 682760 43074 682816
rect 43130 682760 43135 682816
rect 41492 682758 43135 682760
rect 43069 682755 43135 682758
rect 42977 682410 43043 682413
rect 41492 682408 43043 682410
rect 41492 682352 42982 682408
rect 43038 682352 43043 682408
rect 41492 682350 43043 682352
rect 42977 682347 43043 682350
rect 41462 681866 41522 681972
rect 41689 681866 41755 681869
rect 41462 681864 41755 681866
rect 41462 681808 41694 681864
rect 41750 681808 41755 681864
rect 41462 681806 41755 681808
rect 41689 681803 41755 681806
rect 41873 681594 41939 681597
rect 41492 681592 41939 681594
rect 41492 681536 41878 681592
rect 41934 681536 41939 681592
rect 41492 681534 41939 681536
rect 41873 681531 41939 681534
rect 43805 681186 43871 681189
rect 41492 681184 43871 681186
rect 41492 681128 43810 681184
rect 43866 681128 43871 681184
rect 41492 681126 43871 681128
rect 43805 681123 43871 681126
rect 43253 680778 43319 680781
rect 41492 680776 43319 680778
rect 41492 680720 43258 680776
rect 43314 680720 43319 680776
rect 41492 680718 43319 680720
rect 43253 680715 43319 680718
rect 43437 680370 43503 680373
rect 41492 680368 43503 680370
rect 41492 680312 43442 680368
rect 43498 680312 43503 680368
rect 41492 680310 43503 680312
rect 43437 680307 43503 680310
rect 43713 679962 43779 679965
rect 41492 679960 43779 679962
rect 41492 679904 43718 679960
rect 43774 679904 43779 679960
rect 41492 679902 43779 679904
rect 43713 679899 43779 679902
rect 43529 679554 43595 679557
rect 41492 679552 43595 679554
rect 41492 679496 43534 679552
rect 43590 679496 43595 679552
rect 41492 679494 43595 679496
rect 43529 679491 43595 679494
rect 43989 679146 44055 679149
rect 41492 679144 44055 679146
rect 41492 679088 43994 679144
rect 44050 679088 44055 679144
rect 41492 679086 44055 679088
rect 43989 679083 44055 679086
rect 41781 678738 41847 678741
rect 41492 678736 41847 678738
rect 41492 678680 41786 678736
rect 41842 678680 41847 678736
rect 41492 678678 41847 678680
rect 41781 678675 41847 678678
rect 41965 678330 42031 678333
rect 41492 678328 42031 678330
rect 41492 678272 41970 678328
rect 42026 678272 42031 678328
rect 41492 678270 42031 678272
rect 41965 678267 42031 678270
rect 41781 677922 41847 677925
rect 41492 677920 41847 677922
rect 41492 677864 41786 677920
rect 41842 677864 41847 677920
rect 41492 677862 41847 677864
rect 41781 677859 41847 677862
rect 30422 677076 30482 677484
rect 41781 676698 41847 676701
rect 41492 676696 41847 676698
rect 41492 676640 41786 676696
rect 41842 676640 41847 676696
rect 41492 676638 41847 676640
rect 41781 676635 41847 676638
rect 58433 676154 58499 676157
rect 58433 676152 64492 676154
rect 58433 676096 58438 676152
rect 58494 676096 64492 676152
rect 58433 676094 64492 676096
rect 58433 676091 58499 676094
rect 676213 671530 676279 671533
rect 676213 671528 676322 671530
rect 676213 671472 676218 671528
rect 676274 671472 676322 671528
rect 676213 671467 676322 671472
rect 676262 671364 676322 671467
rect 676029 670986 676095 670989
rect 676029 670984 676292 670986
rect 676029 670928 676034 670984
rect 676090 670928 676292 670984
rect 676029 670926 676292 670928
rect 676029 670923 676095 670926
rect 676029 670578 676095 670581
rect 676029 670576 676292 670578
rect 676029 670520 676034 670576
rect 676090 670520 676292 670576
rect 676029 670518 676292 670520
rect 676029 670515 676095 670518
rect 655513 670442 655579 670445
rect 650164 670440 655579 670442
rect 650164 670384 655518 670440
rect 655574 670384 655579 670440
rect 650164 670382 655579 670384
rect 655513 670379 655579 670382
rect 676213 670306 676279 670309
rect 676213 670304 676322 670306
rect 676213 670248 676218 670304
rect 676274 670248 676322 670304
rect 676213 670243 676322 670248
rect 676262 670140 676322 670243
rect 676029 669762 676095 669765
rect 676029 669760 676292 669762
rect 676029 669704 676034 669760
rect 676090 669704 676292 669760
rect 676029 669702 676292 669704
rect 676029 669699 676095 669702
rect 678973 669490 679039 669493
rect 678973 669488 679082 669490
rect 678973 669432 678978 669488
rect 679034 669432 679082 669488
rect 678973 669427 679082 669432
rect 679022 669324 679082 669427
rect 676029 668946 676095 668949
rect 676029 668944 676292 668946
rect 676029 668888 676034 668944
rect 676090 668888 676292 668944
rect 676029 668886 676292 668888
rect 676029 668883 676095 668886
rect 676213 668674 676279 668677
rect 676213 668672 676322 668674
rect 676213 668616 676218 668672
rect 676274 668616 676322 668672
rect 676213 668611 676322 668616
rect 676262 668508 676322 668611
rect 675937 668130 676003 668133
rect 675937 668128 676292 668130
rect 675937 668072 675942 668128
rect 675998 668072 676292 668128
rect 675937 668070 676292 668072
rect 675937 668067 676003 668070
rect 675937 667722 676003 667725
rect 675937 667720 676292 667722
rect 675937 667664 675942 667720
rect 675998 667664 676292 667720
rect 675937 667662 676292 667664
rect 675937 667659 676003 667662
rect 677366 667044 677426 667284
rect 677358 666980 677364 667044
rect 677428 666980 677434 667044
rect 674046 666844 674052 666908
rect 674116 666906 674122 666908
rect 674116 666846 676292 666906
rect 674116 666844 674122 666846
rect 676121 666634 676187 666637
rect 676121 666632 676322 666634
rect 676121 666576 676126 666632
rect 676182 666576 676322 666632
rect 676121 666574 676322 666576
rect 676121 666571 676187 666574
rect 676262 666468 676322 666574
rect 675886 666028 675892 666092
rect 675956 666090 675962 666092
rect 675956 666030 676292 666090
rect 675956 666028 675962 666030
rect 673862 665620 673868 665684
rect 673932 665682 673938 665684
rect 673932 665622 676292 665682
rect 673932 665620 673938 665622
rect 676029 665274 676095 665277
rect 676029 665272 676292 665274
rect 676029 665216 676034 665272
rect 676090 665216 676292 665272
rect 676029 665214 676292 665216
rect 676029 665211 676095 665214
rect 676029 664866 676095 664869
rect 676029 664864 676292 664866
rect 676029 664808 676034 664864
rect 676090 664808 676292 664864
rect 676029 664806 676292 664808
rect 676029 664803 676095 664806
rect 676070 664532 676076 664596
rect 676140 664594 676146 664596
rect 676140 664534 676322 664594
rect 676140 664532 676146 664534
rect 676262 664428 676322 664534
rect 673678 663988 673684 664052
rect 673748 664050 673754 664052
rect 673748 663990 676292 664050
rect 673748 663988 673754 663990
rect 675702 663580 675708 663644
rect 675772 663642 675778 663644
rect 675772 663582 676292 663642
rect 675772 663580 675778 663582
rect 676029 663234 676095 663237
rect 676029 663232 676292 663234
rect 676029 663176 676034 663232
rect 676090 663176 676292 663232
rect 676029 663174 676292 663176
rect 676029 663171 676095 663174
rect 58433 663098 58499 663101
rect 58433 663096 64492 663098
rect 58433 663040 58438 663096
rect 58494 663040 64492 663096
rect 58433 663038 64492 663040
rect 58433 663035 58499 663038
rect 676254 662900 676260 662964
rect 676324 662900 676330 662964
rect 676262 662796 676322 662900
rect 676438 662492 676444 662556
rect 676508 662492 676514 662556
rect 676446 662388 676506 662492
rect 676990 662084 676996 662148
rect 677060 662084 677066 662148
rect 676998 661980 677058 662084
rect 676806 661676 676812 661740
rect 676876 661676 676882 661740
rect 676814 661572 676874 661676
rect 679022 660925 679082 661164
rect 678973 660920 679082 660925
rect 678973 660864 678978 660920
rect 679034 660864 679082 660920
rect 678973 660862 679082 660864
rect 678973 660859 679039 660862
rect 684542 660348 684602 660756
rect 678973 660106 679039 660109
rect 678973 660104 679082 660106
rect 678973 660048 678978 660104
rect 679034 660048 679082 660104
rect 678973 660043 679082 660048
rect 679022 659940 679082 660043
rect 656157 657114 656223 657117
rect 650164 657112 656223 657114
rect 650164 657056 656162 657112
rect 656218 657056 656223 657112
rect 650164 657054 656223 657056
rect 656157 657051 656223 657054
rect 675150 652564 675156 652628
rect 675220 652626 675226 652628
rect 675385 652626 675451 652629
rect 675220 652624 675451 652626
rect 675220 652568 675390 652624
rect 675446 652568 675451 652624
rect 675220 652566 675451 652568
rect 675220 652564 675226 652566
rect 675385 652563 675451 652566
rect 674966 652156 674972 652220
rect 675036 652218 675042 652220
rect 675477 652218 675543 652221
rect 675036 652216 675543 652218
rect 675036 652160 675482 652216
rect 675538 652160 675543 652216
rect 675036 652158 675543 652160
rect 675036 652156 675042 652158
rect 675477 652155 675543 652158
rect 674782 651612 674788 651676
rect 674852 651674 674858 651676
rect 675385 651674 675451 651677
rect 674852 651672 675451 651674
rect 674852 651616 675390 651672
rect 675446 651616 675451 651672
rect 674852 651614 675451 651616
rect 674852 651612 674858 651614
rect 675385 651611 675451 651614
rect 59169 650042 59235 650045
rect 59169 650040 64492 650042
rect 59169 649984 59174 650040
rect 59230 649984 64492 650040
rect 59169 649982 64492 649984
rect 59169 649979 59235 649982
rect 675753 649226 675819 649229
rect 675886 649226 675892 649228
rect 675753 649224 675892 649226
rect 675753 649168 675758 649224
rect 675814 649168 675892 649224
rect 675753 649166 675892 649168
rect 675753 649163 675819 649166
rect 675886 649164 675892 649166
rect 675956 649164 675962 649228
rect 675661 648684 675727 648685
rect 675661 648680 675708 648684
rect 675772 648682 675778 648684
rect 675661 648624 675666 648680
rect 675661 648620 675708 648624
rect 675772 648622 675818 648682
rect 675772 648620 675778 648622
rect 675661 648619 675727 648620
rect 41505 645146 41571 645149
rect 41462 645144 41571 645146
rect 41462 645088 41510 645144
rect 41566 645088 41571 645144
rect 41462 645083 41571 645088
rect 41462 644912 41522 645083
rect 41781 644534 41847 644537
rect 41492 644532 41847 644534
rect 41492 644476 41786 644532
rect 41842 644476 41847 644532
rect 41492 644474 41847 644476
rect 41781 644471 41847 644474
rect 41505 644330 41571 644333
rect 41462 644328 41571 644330
rect 41462 644272 41510 644328
rect 41566 644272 41571 644328
rect 41462 644267 41571 644272
rect 41462 644096 41522 644267
rect 654869 643786 654935 643789
rect 650164 643784 654935 643786
rect 650164 643728 654874 643784
rect 654930 643728 654935 643784
rect 650164 643726 654935 643728
rect 654869 643723 654935 643726
rect 39982 643452 39988 643516
rect 40052 643452 40058 643516
rect 41462 643514 41522 643688
rect 43662 643514 43668 643516
rect 41462 643454 43668 643514
rect 43662 643452 43668 643454
rect 43732 643514 43738 643516
rect 44081 643514 44147 643517
rect 43732 643512 44147 643514
rect 43732 643456 44086 643512
rect 44142 643456 44147 643512
rect 43732 643454 44147 643456
rect 43732 643452 43738 643454
rect 39990 643280 40050 643452
rect 44081 643451 44147 643454
rect 43161 643106 43227 643109
rect 41462 643104 43227 643106
rect 41462 643048 43166 643104
rect 43222 643048 43227 643104
rect 41462 643046 43227 643048
rect 41462 642872 41522 643046
rect 43161 643043 43227 643046
rect 41462 642290 41522 642464
rect 44817 642290 44883 642293
rect 41462 642288 44883 642290
rect 41462 642232 44822 642288
rect 44878 642232 44883 642288
rect 41462 642230 44883 642232
rect 44817 642227 44883 642230
rect 41462 642018 41522 642056
rect 44357 642018 44423 642021
rect 41462 642016 44423 642018
rect 41462 641960 44362 642016
rect 44418 641960 44423 642016
rect 41462 641958 44423 641960
rect 44357 641955 44423 641958
rect 43345 641882 43411 641885
rect 41462 641880 43411 641882
rect 41462 641824 43350 641880
rect 43406 641824 43411 641880
rect 41462 641822 43411 641824
rect 41462 641648 41522 641822
rect 43345 641819 43411 641822
rect 41462 641202 41522 641240
rect 44633 641202 44699 641205
rect 41462 641200 44699 641202
rect 41462 641144 44638 641200
rect 44694 641144 44699 641200
rect 41462 641142 44699 641144
rect 44633 641139 44699 641142
rect 42793 641066 42859 641069
rect 41462 641064 42859 641066
rect 41462 641008 42798 641064
rect 42854 641008 42859 641064
rect 41462 641006 42859 641008
rect 41462 640832 41522 641006
rect 42793 641003 42859 641006
rect 41462 640386 41522 640424
rect 43345 640386 43411 640389
rect 41462 640384 43411 640386
rect 41462 640328 43350 640384
rect 43406 640328 43411 640384
rect 41462 640326 43411 640328
rect 43345 640323 43411 640326
rect 41462 639842 41522 640016
rect 43713 639842 43779 639845
rect 41462 639840 43779 639842
rect 41462 639784 43718 639840
rect 43774 639784 43779 639840
rect 41462 639782 43779 639784
rect 43713 639779 43779 639782
rect 41462 639434 41522 639608
rect 42793 639434 42859 639437
rect 41462 639432 42859 639434
rect 41462 639376 42798 639432
rect 42854 639376 42859 639432
rect 41462 639374 42859 639376
rect 42793 639371 42859 639374
rect 41462 639026 41522 639200
rect 43529 639026 43595 639029
rect 41462 639024 43595 639026
rect 41462 638968 43534 639024
rect 43590 638968 43595 639024
rect 41462 638966 43595 638968
rect 43529 638963 43595 638966
rect 41462 638618 41522 638792
rect 43897 638618 43963 638621
rect 41462 638616 43963 638618
rect 41462 638560 43902 638616
rect 43958 638560 43963 638616
rect 41462 638558 43963 638560
rect 43897 638555 43963 638558
rect 41781 638414 41847 638417
rect 41492 638412 41847 638414
rect 41492 638356 41786 638412
rect 41842 638356 41847 638412
rect 41492 638354 41847 638356
rect 41781 638351 41847 638354
rect 41462 637802 41522 637976
rect 42977 637802 43043 637805
rect 41462 637800 43043 637802
rect 41462 637744 42982 637800
rect 43038 637744 43043 637800
rect 41462 637742 43043 637744
rect 42977 637739 43043 637742
rect 42885 637666 42951 637669
rect 41462 637664 42951 637666
rect 41462 637608 42890 637664
rect 42946 637608 42951 637664
rect 41462 637606 42951 637608
rect 41462 637568 41522 637606
rect 42885 637603 42951 637606
rect 41462 636986 41522 637160
rect 58433 637122 58499 637125
rect 58433 637120 64492 637122
rect 58433 637064 58438 637120
rect 58494 637064 64492 637120
rect 58433 637062 64492 637064
rect 58433 637059 58499 637062
rect 43437 636986 43503 636989
rect 41462 636984 43503 636986
rect 41462 636928 43442 636984
rect 43498 636928 43503 636984
rect 41462 636926 43503 636928
rect 43437 636923 43503 636926
rect 41462 636578 41522 636752
rect 43069 636578 43135 636581
rect 41462 636576 43135 636578
rect 41462 636520 43074 636576
rect 43130 636520 43135 636576
rect 41462 636518 43135 636520
rect 43069 636515 43135 636518
rect 41462 636170 41522 636344
rect 43253 636170 43319 636173
rect 41462 636168 43319 636170
rect 41462 636112 43258 636168
rect 43314 636112 43319 636168
rect 41462 636110 43319 636112
rect 43253 636107 43319 636110
rect 41462 635762 41522 635936
rect 43805 635762 43871 635765
rect 41462 635760 43871 635762
rect 41462 635704 43810 635760
rect 43866 635704 43871 635760
rect 41462 635702 43871 635704
rect 43805 635699 43871 635702
rect 41462 635354 41522 635528
rect 43161 635354 43227 635357
rect 41462 635352 43227 635354
rect 41462 635296 43166 635352
rect 43222 635296 43227 635352
rect 41462 635294 43227 635296
rect 43161 635291 43227 635294
rect 30238 634949 30298 635120
rect 30238 634944 30347 634949
rect 30238 634888 30286 634944
rect 30342 634888 30347 634944
rect 30238 634886 30347 634888
rect 30281 634883 30347 634886
rect 41462 634541 41522 634712
rect 41462 634536 41571 634541
rect 41462 634480 41510 634536
rect 41566 634480 41571 634536
rect 41462 634478 41571 634480
rect 41505 634475 41571 634478
rect 30422 633896 30482 634304
rect 41462 633317 41522 633488
rect 41462 633312 41571 633317
rect 41462 633256 41510 633312
rect 41566 633256 41571 633312
rect 41462 633254 41571 633256
rect 41505 633251 41571 633254
rect 655053 630594 655119 630597
rect 650164 630592 655119 630594
rect 650164 630536 655058 630592
rect 655114 630536 655119 630592
rect 650164 630534 655119 630536
rect 655053 630531 655119 630534
rect 679022 626109 679082 626348
rect 678973 626104 679082 626109
rect 678973 626048 678978 626104
rect 679034 626048 679082 626104
rect 678973 626046 679082 626048
rect 678973 626043 679039 626046
rect 676262 625701 676322 625940
rect 676213 625696 676322 625701
rect 676213 625640 676218 625696
rect 676274 625640 676322 625696
rect 676213 625638 676322 625640
rect 676213 625635 676279 625638
rect 676262 625293 676322 625532
rect 676262 625288 676371 625293
rect 676262 625232 676310 625288
rect 676366 625232 676371 625288
rect 676262 625230 676371 625232
rect 676305 625227 676371 625230
rect 676029 625154 676095 625157
rect 676029 625152 676292 625154
rect 676029 625096 676034 625152
rect 676090 625096 676292 625152
rect 676029 625094 676292 625096
rect 676029 625091 676095 625094
rect 676121 624474 676187 624477
rect 676262 624474 676322 624716
rect 679065 624474 679131 624477
rect 676121 624472 676322 624474
rect 676121 624416 676126 624472
rect 676182 624416 676322 624472
rect 676121 624414 676322 624416
rect 679022 624472 679131 624474
rect 679022 624416 679070 624472
rect 679126 624416 679131 624472
rect 676121 624411 676187 624414
rect 679022 624411 679131 624416
rect 679022 624308 679082 624411
rect 58433 624066 58499 624069
rect 58433 624064 64492 624066
rect 58433 624008 58438 624064
rect 58494 624008 64492 624064
rect 58433 624006 64492 624008
rect 58433 624003 58499 624006
rect 676029 623930 676095 623933
rect 676029 623928 676292 623930
rect 676029 623872 676034 623928
rect 676090 623872 676292 623928
rect 676029 623870 676292 623872
rect 676029 623867 676095 623870
rect 679157 623658 679223 623661
rect 679022 623656 679223 623658
rect 679022 623600 679162 623656
rect 679218 623600 679223 623656
rect 679022 623598 679223 623600
rect 679022 623253 679082 623598
rect 679157 623595 679223 623598
rect 678973 623248 679082 623253
rect 678973 623192 678978 623248
rect 679034 623192 679082 623248
rect 678973 623190 679082 623192
rect 678973 623187 679039 623190
rect 673678 623052 673684 623116
rect 673748 623114 673754 623116
rect 673748 623054 676292 623114
rect 673748 623052 673754 623054
rect 677358 622780 677364 622844
rect 677428 622780 677434 622844
rect 677366 622706 677426 622780
rect 676292 622676 677426 622706
rect 676262 622646 677396 622676
rect 676262 622436 676322 622646
rect 676254 622372 676260 622436
rect 676324 622372 676330 622436
rect 676262 622029 676322 622268
rect 676213 622024 676322 622029
rect 676213 621968 676218 622024
rect 676274 621968 676322 622024
rect 676213 621966 676322 621968
rect 676213 621963 676279 621966
rect 674230 621828 674236 621892
rect 674300 621890 674306 621892
rect 674300 621830 676292 621890
rect 674300 621828 674306 621830
rect 670417 621618 670483 621621
rect 673678 621618 673684 621620
rect 670417 621616 673684 621618
rect 670417 621560 670422 621616
rect 670478 621560 673684 621616
rect 670417 621558 673684 621560
rect 670417 621555 670483 621558
rect 673678 621556 673684 621558
rect 673748 621556 673754 621620
rect 676029 621482 676095 621485
rect 676029 621480 676292 621482
rect 676029 621424 676034 621480
rect 676090 621424 676292 621480
rect 676029 621422 676292 621424
rect 676029 621419 676095 621422
rect 675518 621012 675524 621076
rect 675588 621074 675594 621076
rect 675588 621014 676292 621074
rect 675588 621012 675594 621014
rect 674414 620604 674420 620668
rect 674484 620666 674490 620668
rect 674484 620606 676292 620666
rect 674484 620604 674490 620606
rect 676121 620394 676187 620397
rect 676121 620392 676322 620394
rect 676121 620336 676126 620392
rect 676182 620336 676322 620392
rect 676121 620334 676322 620336
rect 676121 620331 676187 620334
rect 676262 620228 676322 620334
rect 676029 619850 676095 619853
rect 676029 619848 676292 619850
rect 676029 619792 676034 619848
rect 676090 619792 676292 619848
rect 676029 619790 676292 619792
rect 676029 619787 676095 619790
rect 670417 619578 670483 619581
rect 676070 619578 676076 619580
rect 670417 619576 676076 619578
rect 670417 619520 670422 619576
rect 670478 619520 676076 619576
rect 670417 619518 676076 619520
rect 670417 619515 670483 619518
rect 676070 619516 676076 619518
rect 676140 619516 676146 619580
rect 675334 619380 675340 619444
rect 675404 619442 675410 619444
rect 675404 619382 676292 619442
rect 675404 619380 675410 619382
rect 674598 618972 674604 619036
rect 674668 619034 674674 619036
rect 674668 618974 676292 619034
rect 674668 618972 674674 618974
rect 673494 618564 673500 618628
rect 673564 618626 673570 618628
rect 673564 618566 676292 618626
rect 673564 618564 673570 618566
rect 676029 618218 676095 618221
rect 676029 618216 676292 618218
rect 676029 618160 676034 618216
rect 676090 618160 676292 618216
rect 676029 618158 676292 618160
rect 676029 618155 676095 618158
rect 676213 617946 676279 617949
rect 676213 617944 676322 617946
rect 676213 617888 676218 617944
rect 676274 617888 676322 617944
rect 676213 617883 676322 617888
rect 676262 617780 676322 617883
rect 677174 617476 677180 617540
rect 677244 617476 677250 617540
rect 677182 617372 677242 617476
rect 654593 617266 654659 617269
rect 650164 617264 654659 617266
rect 650164 617208 654598 617264
rect 654654 617208 654659 617264
rect 650164 617206 654659 617208
rect 654593 617203 654659 617206
rect 676622 617068 676628 617132
rect 676692 617068 676698 617132
rect 676630 616964 676690 617068
rect 676213 616722 676279 616725
rect 676213 616720 676322 616722
rect 676213 616664 676218 616720
rect 676274 616664 676322 616720
rect 676213 616659 676322 616664
rect 676262 616556 676322 616659
rect 679022 615909 679082 616148
rect 678973 615904 679082 615909
rect 678973 615848 678978 615904
rect 679034 615848 679082 615904
rect 678973 615846 679082 615848
rect 678973 615843 679039 615846
rect 679022 615332 679082 615740
rect 678973 615090 679039 615093
rect 678973 615088 679082 615090
rect 678973 615032 678978 615088
rect 679034 615032 679082 615088
rect 678973 615027 679082 615032
rect 679022 614924 679082 615027
rect 58433 611010 58499 611013
rect 58433 611008 64492 611010
rect 58433 610952 58438 611008
rect 58494 610952 64492 611008
rect 58433 610950 64492 610952
rect 58433 610947 58499 610950
rect 674373 607746 674439 607749
rect 676438 607746 676444 607748
rect 674373 607744 676444 607746
rect 674373 607688 674378 607744
rect 674434 607688 676444 607744
rect 674373 607686 676444 607688
rect 674373 607683 674439 607686
rect 676438 607684 676444 607686
rect 676508 607684 676514 607748
rect 675477 607612 675543 607613
rect 675477 607608 675524 607612
rect 675588 607610 675594 607612
rect 675477 607552 675482 607608
rect 675477 607548 675524 607552
rect 675588 607550 675634 607610
rect 675588 607548 675594 607550
rect 675477 607547 675543 607548
rect 674741 607474 674807 607477
rect 676622 607474 676628 607476
rect 674741 607472 676628 607474
rect 674741 607416 674746 607472
rect 674802 607416 676628 607472
rect 674741 607414 676628 607416
rect 674741 607411 674807 607414
rect 676622 607412 676628 607414
rect 676692 607412 676698 607476
rect 675753 607338 675819 607341
rect 676070 607338 676076 607340
rect 675753 607336 676076 607338
rect 675753 607280 675758 607336
rect 675814 607280 676076 607336
rect 675753 607278 676076 607280
rect 675753 607275 675819 607278
rect 676070 607276 676076 607278
rect 676140 607276 676146 607340
rect 674414 606460 674420 606524
rect 674484 606522 674490 606524
rect 675385 606522 675451 606525
rect 674484 606520 675451 606522
rect 674484 606464 675390 606520
rect 675446 606464 675451 606520
rect 674484 606462 675451 606464
rect 674484 606460 674490 606462
rect 675385 606459 675451 606462
rect 674230 604692 674236 604756
rect 674300 604754 674306 604756
rect 675385 604754 675451 604757
rect 674300 604752 675451 604754
rect 674300 604696 675390 604752
rect 675446 604696 675451 604752
rect 674300 604694 675451 604696
rect 674300 604692 674306 604694
rect 675385 604691 675451 604694
rect 675385 604348 675451 604349
rect 675334 604346 675340 604348
rect 675294 604286 675340 604346
rect 675404 604344 675451 604348
rect 675446 604288 675451 604344
rect 675334 604284 675340 604286
rect 675404 604284 675451 604288
rect 675385 604283 675451 604284
rect 654317 603938 654383 603941
rect 650164 603936 654383 603938
rect 650164 603880 654322 603936
rect 654378 603880 654383 603936
rect 650164 603878 654383 603880
rect 654317 603875 654383 603878
rect 674598 603468 674604 603532
rect 674668 603530 674674 603532
rect 675477 603530 675543 603533
rect 674668 603528 675543 603530
rect 674668 603472 675482 603528
rect 675538 603472 675543 603528
rect 674668 603470 675543 603472
rect 674668 603468 674674 603470
rect 675477 603467 675543 603470
rect 675753 602986 675819 602989
rect 676254 602986 676260 602988
rect 675753 602984 676260 602986
rect 675753 602928 675758 602984
rect 675814 602928 676260 602984
rect 675753 602926 676260 602928
rect 675753 602923 675819 602926
rect 676254 602924 676260 602926
rect 676324 602924 676330 602988
rect 41505 601898 41571 601901
rect 41462 601896 41571 601898
rect 41462 601840 41510 601896
rect 41566 601840 41571 601896
rect 41462 601835 41571 601840
rect 41462 601732 41522 601835
rect 51073 601354 51139 601357
rect 41492 601352 51139 601354
rect 41492 601296 51078 601352
rect 51134 601296 51139 601352
rect 41492 601294 51139 601296
rect 51073 601291 51139 601294
rect 53833 600946 53899 600949
rect 41492 600944 53899 600946
rect 41492 600888 53838 600944
rect 53894 600888 53899 600944
rect 41492 600886 53899 600888
rect 53833 600883 53899 600886
rect 42425 600538 42491 600541
rect 41492 600536 42491 600538
rect 41492 600480 42430 600536
rect 42486 600480 42491 600536
rect 41492 600478 42491 600480
rect 42425 600475 42491 600478
rect 44173 600130 44239 600133
rect 41492 600128 44239 600130
rect 41492 600072 44178 600128
rect 44234 600072 44239 600128
rect 41492 600070 44239 600072
rect 44173 600067 44239 600070
rect 44817 599722 44883 599725
rect 41492 599720 44883 599722
rect 41492 599664 44822 599720
rect 44878 599664 44883 599720
rect 41492 599662 44883 599664
rect 44817 599659 44883 599662
rect 43437 599314 43503 599317
rect 41492 599312 43503 599314
rect 41492 599256 43442 599312
rect 43498 599256 43503 599312
rect 41492 599254 43503 599256
rect 43437 599251 43503 599254
rect 40174 598636 40234 598876
rect 40166 598572 40172 598636
rect 40236 598572 40242 598636
rect 44357 598498 44423 598501
rect 46565 598498 46631 598501
rect 41492 598496 46631 598498
rect 41492 598440 44362 598496
rect 44418 598440 46570 598496
rect 46626 598440 46631 598496
rect 41492 598438 46631 598440
rect 44357 598435 44423 598438
rect 46565 598435 46631 598438
rect 43846 598090 43852 598092
rect 41492 598030 43852 598090
rect 43846 598028 43852 598030
rect 43916 598090 43922 598092
rect 43989 598090 44055 598093
rect 43916 598088 44055 598090
rect 43916 598032 43994 598088
rect 44050 598032 44055 598088
rect 43916 598030 44055 598032
rect 43916 598028 43922 598030
rect 43989 598027 44055 598030
rect 59169 597954 59235 597957
rect 59169 597952 64492 597954
rect 59169 597896 59174 597952
rect 59230 597896 64492 597952
rect 59169 597894 64492 597896
rect 59169 597891 59235 597894
rect 44633 597682 44699 597685
rect 46749 597682 46815 597685
rect 41492 597680 46815 597682
rect 41492 597624 44638 597680
rect 44694 597624 46754 597680
rect 46810 597624 46815 597680
rect 41492 597622 46815 597624
rect 44633 597619 44699 597622
rect 46749 597619 46815 597622
rect 43253 597274 43319 597277
rect 41492 597272 43319 597274
rect 41492 597216 43258 597272
rect 43314 597216 43319 597272
rect 41492 597214 43319 597216
rect 43253 597211 43319 597214
rect 42885 596866 42951 596869
rect 41492 596864 42951 596866
rect 41492 596808 42890 596864
rect 42946 596808 42951 596864
rect 41492 596806 42951 596808
rect 42885 596803 42951 596806
rect 43069 596458 43135 596461
rect 41492 596456 43135 596458
rect 41492 596400 43074 596456
rect 43130 596400 43135 596456
rect 41492 596398 43135 596400
rect 43069 596395 43135 596398
rect 40166 596124 40172 596188
rect 40236 596186 40242 596188
rect 62573 596186 62639 596189
rect 40236 596184 62639 596186
rect 40236 596128 62578 596184
rect 62634 596128 62639 596184
rect 40236 596126 62639 596128
rect 40236 596124 40242 596126
rect 62573 596123 62639 596126
rect 43805 596050 43871 596053
rect 41492 596048 43871 596050
rect 41492 595992 43810 596048
rect 43866 595992 43871 596048
rect 41492 595990 43871 595992
rect 43805 595987 43871 595990
rect 43345 595642 43411 595645
rect 41492 595640 43411 595642
rect 41492 595584 43350 595640
rect 43406 595584 43411 595640
rect 41492 595582 43411 595584
rect 43345 595579 43411 595582
rect 41873 595234 41939 595237
rect 41492 595232 41939 595234
rect 41492 595176 41878 595232
rect 41934 595176 41939 595232
rect 41492 595174 41939 595176
rect 41873 595171 41939 595174
rect 42977 594826 43043 594829
rect 41492 594824 43043 594826
rect 41492 594768 42982 594824
rect 43038 594768 43043 594824
rect 41492 594766 43043 594768
rect 42977 594763 43043 594766
rect 41094 594149 41154 594388
rect 41094 594144 41203 594149
rect 41094 594088 41142 594144
rect 41198 594088 41203 594144
rect 41094 594086 41203 594088
rect 41137 594083 41203 594086
rect 43161 594010 43227 594013
rect 41492 594008 43227 594010
rect 41492 593952 43166 594008
rect 43222 593952 43227 594008
rect 41492 593950 43227 593952
rect 43161 593947 43227 593950
rect 42793 593602 42859 593605
rect 41492 593600 42859 593602
rect 41492 593544 42798 593600
rect 42854 593544 42859 593600
rect 41492 593542 42859 593544
rect 42793 593539 42859 593542
rect 43713 593194 43779 593197
rect 41492 593192 43779 593194
rect 41492 593136 43718 593192
rect 43774 593136 43779 593192
rect 41492 593134 43779 593136
rect 43713 593131 43779 593134
rect 43897 592786 43963 592789
rect 41492 592784 43963 592786
rect 41492 592728 43902 592784
rect 43958 592728 43963 592784
rect 41492 592726 43963 592728
rect 43897 592723 43963 592726
rect 43621 592378 43687 592381
rect 41492 592376 43687 592378
rect 41492 592320 43626 592376
rect 43682 592320 43687 592376
rect 41492 592318 43687 592320
rect 43621 592315 43687 592318
rect 43529 591970 43595 591973
rect 41492 591968 43595 591970
rect 41492 591912 43534 591968
rect 43590 591912 43595 591968
rect 41492 591910 43595 591912
rect 43529 591907 43595 591910
rect 41462 591293 41522 591532
rect 41462 591288 41571 591293
rect 41462 591232 41510 591288
rect 41566 591232 41571 591288
rect 41462 591230 41571 591232
rect 41505 591227 41571 591230
rect 30422 590716 30482 591124
rect 656801 590746 656867 590749
rect 650164 590744 656867 590746
rect 650164 590688 656806 590744
rect 656862 590688 656867 590744
rect 650164 590686 656867 590688
rect 656801 590683 656867 590686
rect 41462 590069 41522 590308
rect 41462 590064 41571 590069
rect 41462 590008 41510 590064
rect 41566 590008 41571 590064
rect 41462 590006 41571 590008
rect 41505 590003 41571 590006
rect 58433 584898 58499 584901
rect 58433 584896 64492 584898
rect 58433 584840 58438 584896
rect 58494 584840 64492 584896
rect 58433 584838 64492 584840
rect 58433 584835 58499 584838
rect 676262 580957 676322 581060
rect 676262 580952 676371 580957
rect 676262 580896 676310 580952
rect 676366 580896 676371 580952
rect 676262 580894 676371 580896
rect 676305 580891 676371 580894
rect 676121 580546 676187 580549
rect 676262 580546 676322 580652
rect 676121 580544 676322 580546
rect 676121 580488 676126 580544
rect 676182 580488 676322 580544
rect 676121 580486 676322 580488
rect 676121 580483 676187 580486
rect 676262 580141 676322 580244
rect 676213 580136 676322 580141
rect 676213 580080 676218 580136
rect 676274 580080 676322 580136
rect 676213 580078 676322 580080
rect 676213 580075 676279 580078
rect 676029 579866 676095 579869
rect 676029 579864 676292 579866
rect 676029 579808 676034 579864
rect 676090 579808 676292 579864
rect 676029 579806 676292 579808
rect 676029 579803 676095 579806
rect 676262 579325 676322 579428
rect 676213 579320 676322 579325
rect 676213 579264 676218 579320
rect 676274 579264 676322 579320
rect 676213 579262 676322 579264
rect 678973 579322 679039 579325
rect 678973 579320 679082 579322
rect 678973 579264 678978 579320
rect 679034 579264 679082 579320
rect 676213 579259 676279 579262
rect 678973 579259 679082 579264
rect 679022 579020 679082 579259
rect 676262 578509 676322 578612
rect 676213 578504 676322 578509
rect 676213 578448 676218 578504
rect 676274 578448 676322 578504
rect 676213 578446 676322 578448
rect 676213 578443 676279 578446
rect 674046 578172 674052 578236
rect 674116 578234 674122 578236
rect 674116 578174 676292 578234
rect 674116 578172 674122 578174
rect 676262 577693 676322 577796
rect 676213 577688 676322 577693
rect 676213 577632 676218 577688
rect 676274 577632 676322 577688
rect 676213 577630 676322 577632
rect 676213 577627 676279 577630
rect 655053 577418 655119 577421
rect 650164 577416 655119 577418
rect 650164 577360 655058 577416
rect 655114 577360 655119 577416
rect 650164 577358 655119 577360
rect 655053 577355 655119 577358
rect 676262 577285 676322 577388
rect 676213 577280 676322 577285
rect 676213 577224 676218 577280
rect 676274 577224 676322 577280
rect 676213 577222 676322 577224
rect 676213 577219 676279 577222
rect 676029 577010 676095 577013
rect 676029 577008 676292 577010
rect 676029 576952 676034 577008
rect 676090 576952 676292 577008
rect 676029 576950 676292 576952
rect 676029 576947 676095 576950
rect 674782 576540 674788 576604
rect 674852 576602 674858 576604
rect 674852 576542 676292 576602
rect 674852 576540 674858 576542
rect 675937 576194 676003 576197
rect 675937 576192 676292 576194
rect 675937 576136 675942 576192
rect 675998 576136 676292 576192
rect 675937 576134 676292 576136
rect 675937 576131 676003 576134
rect 675150 575724 675156 575788
rect 675220 575786 675226 575788
rect 675220 575726 676292 575786
rect 675220 575724 675226 575726
rect 676121 575650 676187 575653
rect 676121 575648 676322 575650
rect 676121 575592 676126 575648
rect 676182 575592 676322 575648
rect 676121 575590 676322 575592
rect 676121 575587 676187 575590
rect 676262 575348 676322 575590
rect 675937 574970 676003 574973
rect 675937 574968 676292 574970
rect 675937 574912 675942 574968
rect 675998 574912 676292 574968
rect 675937 574910 676292 574912
rect 675937 574907 676003 574910
rect 676029 574562 676095 574565
rect 676029 574560 676292 574562
rect 676029 574504 676034 574560
rect 676090 574504 676292 574560
rect 676029 574502 676292 574504
rect 676029 574499 676095 574502
rect 674966 574092 674972 574156
rect 675036 574154 675042 574156
rect 675036 574094 676292 574154
rect 675036 574092 675042 574094
rect 675886 573684 675892 573748
rect 675956 573746 675962 573748
rect 675956 573686 676292 573746
rect 675956 573684 675962 573686
rect 675702 573276 675708 573340
rect 675772 573338 675778 573340
rect 675772 573278 676292 573338
rect 675772 573276 675778 573278
rect 676029 572930 676095 572933
rect 676029 572928 676292 572930
rect 676029 572872 676034 572928
rect 676090 572872 676292 572928
rect 676029 572870 676292 572872
rect 676029 572867 676095 572870
rect 676029 572522 676095 572525
rect 676029 572520 676292 572522
rect 676029 572464 676034 572520
rect 676090 572464 676292 572520
rect 676029 572462 676292 572464
rect 676029 572459 676095 572462
rect 675661 572114 675727 572117
rect 675661 572112 676292 572114
rect 675661 572056 675666 572112
rect 675722 572056 676292 572112
rect 675661 572054 676292 572056
rect 675661 572051 675727 572054
rect 676622 571916 676628 571980
rect 676692 571916 676698 571980
rect 58433 571842 58499 571845
rect 58433 571840 64492 571842
rect 58433 571784 58438 571840
rect 58494 571784 64492 571840
rect 58433 571782 64492 571784
rect 58433 571779 58499 571782
rect 676630 571676 676690 571916
rect 676438 571508 676444 571572
rect 676508 571508 676514 571572
rect 676446 571268 676506 571508
rect 679022 570757 679082 570860
rect 678973 570752 679082 570757
rect 678973 570696 678978 570752
rect 679034 570696 679082 570752
rect 678973 570694 679082 570696
rect 678973 570691 679039 570694
rect 684542 570044 684602 570452
rect 678973 569938 679039 569941
rect 678973 569936 679082 569938
rect 678973 569880 678978 569936
rect 679034 569880 679082 569936
rect 678973 569875 679082 569880
rect 679022 569636 679082 569875
rect 674649 564498 674715 564501
rect 676806 564498 676812 564500
rect 674649 564496 676812 564498
rect 674649 564440 674654 564496
rect 674710 564440 676812 564496
rect 674649 564438 676812 564440
rect 674649 564435 674715 564438
rect 676806 564436 676812 564438
rect 676876 564436 676882 564500
rect 654317 564090 654383 564093
rect 650164 564088 654383 564090
rect 650164 564032 654322 564088
rect 654378 564032 654383 564088
rect 650164 564030 654383 564032
rect 654317 564027 654383 564030
rect 675753 562460 675819 562461
rect 675702 562458 675708 562460
rect 675662 562398 675708 562458
rect 675772 562456 675819 562460
rect 675814 562400 675819 562456
rect 675702 562396 675708 562398
rect 675772 562396 675819 562400
rect 675753 562395 675819 562396
rect 675753 562050 675819 562053
rect 675886 562050 675892 562052
rect 675753 562048 675892 562050
rect 675753 561992 675758 562048
rect 675814 561992 675892 562048
rect 675753 561990 675892 561992
rect 675753 561987 675819 561990
rect 675886 561988 675892 561990
rect 675956 561988 675962 562052
rect 674966 561172 674972 561236
rect 675036 561234 675042 561236
rect 675477 561234 675543 561237
rect 675036 561232 675543 561234
rect 675036 561176 675482 561232
rect 675538 561176 675543 561232
rect 675036 561174 675543 561176
rect 675036 561172 675042 561174
rect 675477 561171 675543 561174
rect 41505 558786 41571 558789
rect 41462 558784 41571 558786
rect 41462 558728 41510 558784
rect 41566 558728 41571 558784
rect 41462 558723 41571 558728
rect 58341 558786 58407 558789
rect 58341 558784 64492 558786
rect 58341 558728 58346 558784
rect 58402 558728 64492 558784
rect 58341 558726 64492 558728
rect 58341 558723 58407 558726
rect 675150 558724 675156 558788
rect 675220 558786 675226 558788
rect 675385 558786 675451 558789
rect 675220 558784 675451 558786
rect 675220 558728 675390 558784
rect 675446 558728 675451 558784
rect 675220 558726 675451 558728
rect 675220 558724 675226 558726
rect 675385 558723 675451 558726
rect 41462 558484 41522 558723
rect 41505 558378 41571 558381
rect 41462 558376 41571 558378
rect 41462 558320 41510 558376
rect 41566 558320 41571 558376
rect 41462 558315 41571 558320
rect 675753 558378 675819 558381
rect 676622 558378 676628 558380
rect 675753 558376 676628 558378
rect 675753 558320 675758 558376
rect 675814 558320 676628 558376
rect 675753 558318 676628 558320
rect 675753 558315 675819 558318
rect 676622 558316 676628 558318
rect 676692 558316 676698 558380
rect 41462 558076 41522 558315
rect 41413 557970 41479 557973
rect 41413 557968 41522 557970
rect 41413 557912 41418 557968
rect 41474 557912 41522 557968
rect 41413 557907 41522 557912
rect 41462 557668 41522 557907
rect 675753 557562 675819 557565
rect 676438 557562 676444 557564
rect 675753 557560 676444 557562
rect 675753 557504 675758 557560
rect 675814 557504 676444 557560
rect 675753 557502 676444 557504
rect 675753 557499 675819 557502
rect 676438 557500 676444 557502
rect 676508 557500 676514 557564
rect 43846 557290 43852 557292
rect 41492 557230 43852 557290
rect 43846 557228 43852 557230
rect 43916 557228 43922 557292
rect 42793 556882 42859 556885
rect 41492 556880 42859 556882
rect 41492 556824 42798 556880
rect 42854 556824 42859 556880
rect 41492 556822 42859 556824
rect 42793 556819 42859 556822
rect 43437 556474 43503 556477
rect 41492 556472 43503 556474
rect 41492 556416 43442 556472
rect 43498 556416 43503 556472
rect 41492 556414 43503 556416
rect 43437 556411 43503 556414
rect 43662 556066 43668 556068
rect 41492 556006 43668 556066
rect 43662 556004 43668 556006
rect 43732 556004 43738 556068
rect 39990 555524 40050 555628
rect 39982 555460 39988 555524
rect 40052 555460 40058 555524
rect 40166 555460 40172 555524
rect 40236 555460 40242 555524
rect 40174 555220 40234 555460
rect 41822 554842 41828 554844
rect 41492 554782 41828 554842
rect 41822 554780 41828 554782
rect 41892 554780 41898 554844
rect 43253 554434 43319 554437
rect 41492 554432 43319 554434
rect 41492 554376 43258 554432
rect 43314 554376 43319 554432
rect 41492 554374 43319 554376
rect 43253 554371 43319 554374
rect 43805 554026 43871 554029
rect 41492 554024 43871 554026
rect 41492 553968 43810 554024
rect 43866 553968 43871 554024
rect 41492 553966 43871 553968
rect 43805 553963 43871 553966
rect 42701 553618 42767 553621
rect 41492 553616 42767 553618
rect 41492 553560 42706 553616
rect 42762 553560 42767 553616
rect 41492 553558 42767 553560
rect 42701 553555 42767 553558
rect 43161 553210 43227 553213
rect 41492 553208 43227 553210
rect 41492 553152 43166 553208
rect 43222 553152 43227 553208
rect 41492 553150 43227 553152
rect 43161 553147 43227 553150
rect 43345 552802 43411 552805
rect 41492 552800 43411 552802
rect 41492 552744 43350 552800
rect 43406 552744 43411 552800
rect 41492 552742 43411 552744
rect 43345 552739 43411 552742
rect 43621 552394 43687 552397
rect 41492 552392 43687 552394
rect 41492 552336 43626 552392
rect 43682 552336 43687 552392
rect 41492 552334 43687 552336
rect 43621 552331 43687 552334
rect 41781 551986 41847 551989
rect 41492 551984 41847 551986
rect 41492 551928 41786 551984
rect 41842 551928 41847 551984
rect 41492 551926 41847 551928
rect 41781 551923 41847 551926
rect 43437 551578 43503 551581
rect 41492 551576 43503 551578
rect 41492 551520 43442 551576
rect 43498 551520 43503 551576
rect 41492 551518 43503 551520
rect 43437 551515 43503 551518
rect 43069 551170 43135 551173
rect 41492 551168 43135 551170
rect 41492 551112 43074 551168
rect 43130 551112 43135 551168
rect 41492 551110 43135 551112
rect 43069 551107 43135 551110
rect 654685 550898 654751 550901
rect 650164 550896 654751 550898
rect 650164 550840 654690 550896
rect 654746 550840 654751 550896
rect 650164 550838 654751 550840
rect 654685 550835 654751 550838
rect 43989 550762 44055 550765
rect 41492 550760 44055 550762
rect 41492 550704 43994 550760
rect 44050 550704 44055 550760
rect 41492 550702 44055 550704
rect 43989 550699 44055 550702
rect 42977 550354 43043 550357
rect 41492 550352 43043 550354
rect 41492 550296 42982 550352
rect 43038 550296 43043 550352
rect 41492 550294 43043 550296
rect 42977 550291 43043 550294
rect 43253 549946 43319 549949
rect 41492 549944 43319 549946
rect 41492 549888 43258 549944
rect 43314 549888 43319 549944
rect 41492 549886 43319 549888
rect 43253 549883 43319 549886
rect 43897 549538 43963 549541
rect 41492 549536 43963 549538
rect 41492 549480 43902 549536
rect 43958 549480 43963 549536
rect 41492 549478 43963 549480
rect 43897 549475 43963 549478
rect 41462 548997 41522 549100
rect 41462 548992 41571 548997
rect 41462 548936 41510 548992
rect 41566 548936 41571 548992
rect 41462 548934 41571 548936
rect 41505 548931 41571 548934
rect 41462 548589 41522 548692
rect 41462 548584 41571 548589
rect 41462 548528 41510 548584
rect 41566 548528 41571 548584
rect 41462 548526 41571 548528
rect 41505 548523 41571 548526
rect 41462 548178 41522 548284
rect 41597 548178 41663 548181
rect 41462 548176 41663 548178
rect 41462 548120 41602 548176
rect 41658 548120 41663 548176
rect 41462 548118 41663 548120
rect 41597 548115 41663 548118
rect 30422 547468 30482 547876
rect 41462 546954 41522 547060
rect 41597 546954 41663 546957
rect 41462 546952 41663 546954
rect 41462 546896 41602 546952
rect 41658 546896 41663 546952
rect 41462 546894 41663 546896
rect 41597 546891 41663 546894
rect 58341 545866 58407 545869
rect 58341 545864 64492 545866
rect 58341 545808 58346 545864
rect 58402 545808 64492 545864
rect 58341 545806 64492 545808
rect 58341 545803 58407 545806
rect 41454 540908 41460 540972
rect 41524 540970 41530 540972
rect 42885 540970 42951 540973
rect 41524 540968 42951 540970
rect 41524 540912 42890 540968
rect 42946 540912 42951 540968
rect 41524 540910 42951 540912
rect 41524 540908 41530 540910
rect 42885 540907 42951 540910
rect 41822 540772 41828 540836
rect 41892 540834 41898 540836
rect 44081 540834 44147 540837
rect 41892 540832 44147 540834
rect 41892 540776 44086 540832
rect 44142 540776 44147 540832
rect 41892 540774 44147 540776
rect 41892 540772 41898 540774
rect 44081 540771 44147 540774
rect 654869 537570 654935 537573
rect 650164 537568 654935 537570
rect 650164 537512 654874 537568
rect 654930 537512 654935 537568
rect 650164 537510 654935 537512
rect 654869 537507 654935 537510
rect 676262 535941 676322 536112
rect 676213 535936 676322 535941
rect 676213 535880 676218 535936
rect 676274 535880 676322 535936
rect 676213 535878 676322 535880
rect 676213 535875 676279 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 679022 535125 679082 535296
rect 678973 535120 679082 535125
rect 678973 535064 678978 535120
rect 679034 535064 679082 535120
rect 678973 535062 679082 535064
rect 678973 535059 679039 535062
rect 676029 534918 676095 534921
rect 676029 534916 676292 534918
rect 676029 534860 676034 534916
rect 676090 534860 676292 534916
rect 676029 534858 676292 534860
rect 676029 534855 676095 534858
rect 676121 534306 676187 534309
rect 676262 534306 676322 534480
rect 679065 534306 679131 534309
rect 676121 534304 676322 534306
rect 676121 534248 676126 534304
rect 676182 534248 676322 534304
rect 676121 534246 676322 534248
rect 679022 534304 679131 534306
rect 679022 534248 679070 534304
rect 679126 534248 679131 534304
rect 676121 534243 676187 534246
rect 679022 534243 679131 534248
rect 679022 534072 679082 534243
rect 679022 533493 679082 533664
rect 679022 533488 679131 533493
rect 679022 533432 679070 533488
rect 679126 533432 679131 533488
rect 679022 533430 679131 533432
rect 679065 533427 679131 533430
rect 676029 533286 676095 533289
rect 676029 533284 676292 533286
rect 676029 533228 676034 533284
rect 676090 533228 676292 533284
rect 676029 533226 676292 533228
rect 676029 533223 676095 533226
rect 675937 532878 676003 532881
rect 675937 532876 676292 532878
rect 675937 532820 675942 532876
rect 675998 532820 676292 532876
rect 675937 532818 676292 532820
rect 675937 532815 676003 532818
rect 59261 532810 59327 532813
rect 59261 532808 64492 532810
rect 59261 532752 59266 532808
rect 59322 532752 64492 532808
rect 59261 532750 64492 532752
rect 59261 532747 59327 532750
rect 676213 532674 676279 532677
rect 676213 532672 676322 532674
rect 676213 532616 676218 532672
rect 676274 532616 676322 532672
rect 676213 532611 676322 532616
rect 676262 532440 676322 532611
rect 676121 531858 676187 531861
rect 676262 531858 676322 532032
rect 676121 531856 676322 531858
rect 676121 531800 676126 531856
rect 676182 531800 676322 531856
rect 676121 531798 676322 531800
rect 676121 531795 676187 531798
rect 674414 531660 674420 531724
rect 674484 531722 674490 531724
rect 674484 531662 676322 531722
rect 674484 531660 674490 531662
rect 676262 531624 676322 531662
rect 676029 531246 676095 531249
rect 676029 531244 676292 531246
rect 676029 531188 676034 531244
rect 676090 531188 676292 531244
rect 676029 531186 676292 531188
rect 676029 531183 676095 531186
rect 675518 530980 675524 531044
rect 675588 531042 675594 531044
rect 675588 530982 676322 531042
rect 675588 530980 675594 530982
rect 676262 530808 676322 530982
rect 674230 530572 674236 530636
rect 674300 530634 674306 530636
rect 674300 530574 676322 530634
rect 674300 530572 674306 530574
rect 676262 530400 676322 530574
rect 676029 530022 676095 530025
rect 676029 530020 676292 530022
rect 676029 529964 676034 530020
rect 676090 529964 676292 530020
rect 676029 529962 676292 529964
rect 676029 529959 676095 529962
rect 676029 529614 676095 529617
rect 676029 529612 676292 529614
rect 676029 529556 676034 529612
rect 676090 529556 676292 529612
rect 676029 529554 676292 529556
rect 676029 529551 676095 529554
rect 676070 529348 676076 529412
rect 676140 529410 676146 529412
rect 676140 529350 676322 529410
rect 676140 529348 676146 529350
rect 676262 529176 676322 529350
rect 675334 528940 675340 529004
rect 675404 529002 675410 529004
rect 675404 528942 676322 529002
rect 675404 528940 675410 528942
rect 676262 528768 676322 528942
rect 674598 528532 674604 528596
rect 674668 528594 674674 528596
rect 674668 528534 676322 528594
rect 674668 528532 674674 528534
rect 676262 528360 676322 528534
rect 676029 527982 676095 527985
rect 676029 527980 676292 527982
rect 676029 527924 676034 527980
rect 676090 527924 676292 527980
rect 676029 527922 676292 527924
rect 676029 527919 676095 527922
rect 676029 527574 676095 527577
rect 676029 527572 676292 527574
rect 676029 527516 676034 527572
rect 676090 527516 676292 527572
rect 676029 527514 676292 527516
rect 676029 527511 676095 527514
rect 676254 527308 676260 527372
rect 676324 527308 676330 527372
rect 676262 527136 676322 527308
rect 676806 526900 676812 526964
rect 676876 526900 676882 526964
rect 676814 526728 676874 526900
rect 676029 526350 676095 526353
rect 676029 526348 676292 526350
rect 676029 526292 676034 526348
rect 676090 526292 676292 526348
rect 676029 526290 676292 526292
rect 676029 526287 676095 526290
rect 679022 525741 679082 525912
rect 678973 525736 679082 525741
rect 678973 525680 678978 525736
rect 679034 525680 679082 525736
rect 678973 525678 679082 525680
rect 678973 525675 679039 525678
rect 684542 525096 684602 525504
rect 678973 524922 679039 524925
rect 678973 524920 679082 524922
rect 678973 524864 678978 524920
rect 679034 524864 679082 524920
rect 678973 524859 679082 524864
rect 679022 524688 679082 524859
rect 654133 524242 654199 524245
rect 650164 524240 654199 524242
rect 650164 524184 654138 524240
rect 654194 524184 654199 524240
rect 650164 524182 654199 524184
rect 654133 524179 654199 524182
rect 58433 519754 58499 519757
rect 58433 519752 64492 519754
rect 58433 519696 58438 519752
rect 58494 519696 64492 519752
rect 58433 519694 64492 519696
rect 58433 519691 58499 519694
rect 654869 511050 654935 511053
rect 650164 511048 654935 511050
rect 650164 510992 654874 511048
rect 654930 510992 654935 511048
rect 650164 510990 654935 510992
rect 654869 510987 654935 510990
rect 58433 506698 58499 506701
rect 58433 506696 64492 506698
rect 58433 506640 58438 506696
rect 58494 506640 64492 506696
rect 58433 506638 64492 506640
rect 58433 506635 58499 506638
rect 656801 497722 656867 497725
rect 650164 497720 656867 497722
rect 650164 497664 656806 497720
rect 656862 497664 656867 497720
rect 650164 497662 656867 497664
rect 656801 497659 656867 497662
rect 57973 493642 58039 493645
rect 57973 493640 64492 493642
rect 57973 493584 57978 493640
rect 58034 493584 64492 493640
rect 57973 493582 64492 493584
rect 57973 493579 58039 493582
rect 676438 492356 676444 492420
rect 676508 492418 676514 492420
rect 676806 492418 676812 492420
rect 676508 492358 676812 492418
rect 676508 492356 676514 492358
rect 676806 492356 676812 492358
rect 676876 492356 676882 492420
rect 676029 492146 676095 492149
rect 676029 492144 676292 492146
rect 676029 492088 676034 492144
rect 676090 492088 676292 492144
rect 676029 492086 676292 492088
rect 676029 492083 676095 492086
rect 675937 491738 676003 491741
rect 675937 491736 676292 491738
rect 675937 491680 675942 491736
rect 675998 491680 676292 491736
rect 675937 491678 676292 491680
rect 675937 491675 676003 491678
rect 676029 491330 676095 491333
rect 676029 491328 676292 491330
rect 676029 491272 676034 491328
rect 676090 491272 676292 491328
rect 676029 491270 676292 491272
rect 676029 491267 676095 491270
rect 676029 490922 676095 490925
rect 676029 490920 676292 490922
rect 676029 490864 676034 490920
rect 676090 490864 676292 490920
rect 676029 490862 676292 490864
rect 676029 490859 676095 490862
rect 675937 490514 676003 490517
rect 675937 490512 676292 490514
rect 675937 490456 675942 490512
rect 675998 490456 676292 490512
rect 675937 490454 676292 490456
rect 675937 490451 676003 490454
rect 676029 490106 676095 490109
rect 676029 490104 676292 490106
rect 676029 490048 676034 490104
rect 676090 490048 676292 490104
rect 676029 490046 676292 490048
rect 676029 490043 676095 490046
rect 676029 489698 676095 489701
rect 676029 489696 676292 489698
rect 676029 489640 676034 489696
rect 676090 489640 676292 489696
rect 676029 489638 676292 489640
rect 676029 489635 676095 489638
rect 673678 489228 673684 489292
rect 673748 489290 673754 489292
rect 675845 489290 675911 489293
rect 673748 489288 676292 489290
rect 673748 489232 675850 489288
rect 675906 489232 676292 489288
rect 673748 489230 676292 489232
rect 673748 489228 673754 489230
rect 675845 489227 675911 489230
rect 675845 488882 675911 488885
rect 675845 488880 676292 488882
rect 675845 488824 675850 488880
rect 675906 488824 676292 488880
rect 675845 488822 676292 488824
rect 675845 488819 675911 488822
rect 675569 488474 675635 488477
rect 675569 488472 676292 488474
rect 675569 488416 675574 488472
rect 675630 488416 676292 488472
rect 675569 488414 676292 488416
rect 675569 488411 675635 488414
rect 675937 488066 676003 488069
rect 675937 488064 676292 488066
rect 675937 488008 675942 488064
rect 675998 488008 676292 488064
rect 675937 488006 676292 488008
rect 675937 488003 676003 488006
rect 674966 487596 674972 487660
rect 675036 487658 675042 487660
rect 675036 487598 676292 487658
rect 675036 487596 675042 487598
rect 676029 487250 676095 487253
rect 676029 487248 676292 487250
rect 676029 487192 676034 487248
rect 676090 487192 676292 487248
rect 676029 487190 676292 487192
rect 676029 487187 676095 487190
rect 675702 486780 675708 486844
rect 675772 486842 675778 486844
rect 675772 486782 676292 486842
rect 675772 486780 675778 486782
rect 675661 486434 675727 486437
rect 675661 486432 676292 486434
rect 675661 486376 675666 486432
rect 675722 486376 676292 486432
rect 675661 486374 676292 486376
rect 675661 486371 675727 486374
rect 676029 486026 676095 486029
rect 676029 486024 676292 486026
rect 676029 485968 676034 486024
rect 676090 485968 676292 486024
rect 676029 485966 676292 485968
rect 676029 485963 676095 485966
rect 676029 485618 676095 485621
rect 676029 485616 676292 485618
rect 676029 485560 676034 485616
rect 676090 485560 676292 485616
rect 676029 485558 676292 485560
rect 676029 485555 676095 485558
rect 675886 485148 675892 485212
rect 675956 485210 675962 485212
rect 675956 485150 676292 485210
rect 675956 485148 675962 485150
rect 675150 484740 675156 484804
rect 675220 484802 675226 484804
rect 675220 484742 676292 484802
rect 675220 484740 675226 484742
rect 676070 484468 676076 484532
rect 676140 484468 676146 484532
rect 654869 484394 654935 484397
rect 650164 484392 654935 484394
rect 650164 484336 654874 484392
rect 654930 484336 654935 484392
rect 650164 484334 654935 484336
rect 676078 484394 676138 484468
rect 676078 484334 676292 484394
rect 654869 484331 654935 484334
rect 676029 483986 676095 483989
rect 676029 483984 676292 483986
rect 676029 483928 676034 483984
rect 676090 483928 676292 483984
rect 676029 483926 676292 483928
rect 676029 483923 676095 483926
rect 674005 483578 674071 483581
rect 674005 483576 676292 483578
rect 674005 483520 674010 483576
rect 674066 483520 676292 483576
rect 674005 483518 676292 483520
rect 674005 483515 674071 483518
rect 676814 483002 676874 483140
rect 676806 482938 676812 483002
rect 676876 482938 676882 483002
rect 675661 482762 675727 482765
rect 675661 482760 676292 482762
rect 675661 482704 675666 482760
rect 675722 482704 676292 482760
rect 675661 482702 676292 482704
rect 675661 482699 675727 482702
rect 676029 482354 676095 482357
rect 676029 482352 676292 482354
rect 676029 482296 676034 482352
rect 676090 482296 676292 482352
rect 676029 482294 676292 482296
rect 676029 482291 676095 482294
rect 676029 481946 676095 481949
rect 676029 481944 676292 481946
rect 676029 481888 676034 481944
rect 676090 481888 676292 481944
rect 676029 481886 676292 481888
rect 676029 481883 676095 481886
rect 684542 481100 684602 481508
rect 676029 480722 676095 480725
rect 676029 480720 676292 480722
rect 676029 480664 676034 480720
rect 676090 480664 676292 480720
rect 676029 480662 676292 480664
rect 676029 480659 676095 480662
rect 58433 480586 58499 480589
rect 58433 480584 64492 480586
rect 58433 480528 58438 480584
rect 58494 480528 64492 480584
rect 58433 480526 64492 480528
rect 58433 480523 58499 480526
rect 654869 471202 654935 471205
rect 650164 471200 654935 471202
rect 650164 471144 654874 471200
rect 654930 471144 654935 471200
rect 650164 471142 654935 471144
rect 654869 471139 654935 471142
rect 58709 467530 58775 467533
rect 58709 467528 64492 467530
rect 58709 467472 58714 467528
rect 58770 467472 64492 467528
rect 58709 467470 64492 467472
rect 58709 467467 58775 467470
rect 43846 460124 43852 460188
rect 43916 460124 43922 460188
rect 43854 459916 43914 460124
rect 43846 459852 43852 459916
rect 43916 459852 43922 459916
rect 654225 457874 654291 457877
rect 650164 457872 654291 457874
rect 650164 457816 654230 457872
rect 654286 457816 654291 457872
rect 650164 457814 654291 457816
rect 654225 457811 654291 457814
rect 43662 455908 43668 455972
rect 43732 455970 43738 455972
rect 44030 455970 44036 455972
rect 43732 455910 44036 455970
rect 43732 455908 43738 455910
rect 44030 455908 44036 455910
rect 44100 455908 44106 455972
rect 59169 454610 59235 454613
rect 59169 454608 64492 454610
rect 59169 454552 59174 454608
rect 59230 454552 64492 454608
rect 59169 454550 64492 454552
rect 59169 454547 59235 454550
rect 42885 450802 42951 450805
rect 43662 450802 43668 450804
rect 42885 450800 43668 450802
rect 42885 450744 42890 450800
rect 42946 450744 43668 450800
rect 42885 450742 43668 450744
rect 42885 450739 42951 450742
rect 43662 450740 43668 450742
rect 43732 450740 43738 450804
rect 43662 445844 43668 445908
rect 43732 445906 43738 445908
rect 44214 445906 44220 445908
rect 43732 445846 44220 445906
rect 43732 445844 43738 445846
rect 44214 445844 44220 445846
rect 44284 445844 44290 445908
rect 654409 444546 654475 444549
rect 650164 444544 654475 444546
rect 650164 444488 654414 444544
rect 654470 444488 654475 444544
rect 650164 444486 654475 444488
rect 654409 444483 654475 444486
rect 58433 441554 58499 441557
rect 58433 441552 64492 441554
rect 58433 441496 58438 441552
rect 58494 441496 64492 441552
rect 58433 441494 64492 441496
rect 58433 441491 58499 441494
rect 654685 431354 654751 431357
rect 650164 431352 654751 431354
rect 650164 431296 654690 431352
rect 654746 431296 654751 431352
rect 650164 431294 654751 431296
rect 654685 431291 654751 431294
rect 41781 430946 41847 430949
rect 41492 430944 41847 430946
rect 41492 430888 41786 430944
rect 41842 430888 41847 430944
rect 41492 430886 41847 430888
rect 41781 430883 41847 430886
rect 43069 430674 43135 430677
rect 43662 430674 43668 430676
rect 43069 430672 43668 430674
rect 43069 430616 43074 430672
rect 43130 430616 43668 430672
rect 43069 430614 43668 430616
rect 43069 430611 43135 430614
rect 43662 430612 43668 430614
rect 43732 430674 43738 430676
rect 62573 430674 62639 430677
rect 43732 430672 62639 430674
rect 43732 430616 62578 430672
rect 62634 430616 62639 430672
rect 43732 430614 62639 430616
rect 43732 430612 43738 430614
rect 62573 430611 62639 430614
rect 51257 430538 51323 430541
rect 41492 430536 51323 430538
rect 41492 430480 51262 430536
rect 51318 430480 51323 430536
rect 41492 430478 51323 430480
rect 51257 430475 51323 430478
rect 53833 430130 53899 430133
rect 41492 430128 53899 430130
rect 41492 430072 53838 430128
rect 53894 430072 53899 430128
rect 41492 430070 53899 430072
rect 53833 430067 53899 430070
rect 43621 429722 43687 429725
rect 41492 429720 43687 429722
rect 41492 429664 43626 429720
rect 43682 429664 43687 429720
rect 41492 429662 43687 429664
rect 43621 429659 43687 429662
rect 43069 429314 43135 429317
rect 41492 429312 43135 429314
rect 41492 429256 43074 429312
rect 43130 429256 43135 429312
rect 41492 429254 43135 429256
rect 43069 429251 43135 429254
rect 43846 428906 43852 428908
rect 41492 428846 43852 428906
rect 43846 428844 43852 428846
rect 43916 428844 43922 428908
rect 43805 428498 43871 428501
rect 41492 428496 43871 428498
rect 41492 428440 43810 428496
rect 43866 428440 43871 428496
rect 41492 428438 43871 428440
rect 43805 428435 43871 428438
rect 58249 428498 58315 428501
rect 58249 428496 64492 428498
rect 58249 428440 58254 428496
rect 58310 428440 64492 428496
rect 58249 428438 64492 428440
rect 58249 428435 58315 428438
rect 39982 427858 39988 427922
rect 40052 427858 40058 427922
rect 39990 427682 40050 427858
rect 40358 427854 40418 428060
rect 62941 427954 63007 427957
rect 41692 427952 63007 427954
rect 41692 427920 62946 427952
rect 41278 427896 62946 427920
rect 63002 427896 63007 427952
rect 41278 427894 63007 427896
rect 41278 427860 41752 427894
rect 62941 427891 63007 427894
rect 40350 427790 40356 427854
rect 40420 427790 40426 427854
rect 41278 427682 41338 427860
rect 39990 427652 41338 427682
rect 40020 427622 41308 427652
rect 40028 427274 40034 427276
rect 40020 427214 40034 427274
rect 40028 427212 40034 427214
rect 40098 427212 40104 427276
rect 41781 426866 41847 426869
rect 41492 426864 41847 426866
rect 41492 426808 41786 426864
rect 41842 426808 41847 426864
rect 41492 426806 41847 426808
rect 41781 426803 41847 426806
rect 42885 426458 42951 426461
rect 41492 426456 42951 426458
rect 41492 426400 42890 426456
rect 42946 426400 42951 426456
rect 41492 426398 42951 426400
rect 42885 426395 42951 426398
rect 42793 426050 42859 426053
rect 41492 426048 42859 426050
rect 41492 425992 42798 426048
rect 42854 425992 42859 426048
rect 41492 425990 42859 425992
rect 42793 425987 42859 425990
rect 43253 425642 43319 425645
rect 41492 425640 43319 425642
rect 41492 425584 43258 425640
rect 43314 425584 43319 425640
rect 41492 425582 43319 425584
rect 43253 425579 43319 425582
rect 43345 425234 43411 425237
rect 41492 425232 43411 425234
rect 41492 425176 43350 425232
rect 43406 425176 43411 425232
rect 41492 425174 43411 425176
rect 43345 425171 43411 425174
rect 43437 424826 43503 424829
rect 41492 424824 43503 424826
rect 41492 424768 43442 424824
rect 43498 424768 43503 424824
rect 41492 424766 43503 424768
rect 43437 424763 43503 424766
rect 42333 424418 42399 424421
rect 41492 424416 42399 424418
rect 41492 424360 42338 424416
rect 42394 424360 42399 424416
rect 41492 424358 42399 424360
rect 42333 424355 42399 424358
rect 43897 424010 43963 424013
rect 41492 424008 43963 424010
rect 41492 423952 43902 424008
rect 43958 423952 43963 424008
rect 41492 423950 43963 423952
rect 43897 423947 43963 423950
rect 43713 423602 43779 423605
rect 41492 423600 43779 423602
rect 41492 423544 43718 423600
rect 43774 423544 43779 423600
rect 41492 423542 43779 423544
rect 43713 423539 43779 423542
rect 43529 423194 43595 423197
rect 41492 423192 43595 423194
rect 41492 423136 43534 423192
rect 43590 423136 43595 423192
rect 41492 423134 43595 423136
rect 43529 423131 43595 423134
rect 42977 422786 43043 422789
rect 41492 422784 43043 422786
rect 41492 422728 42982 422784
rect 43038 422728 43043 422784
rect 41492 422726 43043 422728
rect 42977 422723 43043 422726
rect 43161 422378 43227 422381
rect 41492 422376 43227 422378
rect 41492 422320 43166 422376
rect 43222 422320 43227 422376
rect 41492 422318 43227 422320
rect 43161 422315 43227 422318
rect 43989 421970 44055 421973
rect 41492 421968 44055 421970
rect 41492 421912 43994 421968
rect 44050 421912 44055 421968
rect 41492 421910 44055 421912
rect 43989 421907 44055 421910
rect 41873 421562 41939 421565
rect 41492 421560 41939 421562
rect 41492 421504 41878 421560
rect 41934 421504 41939 421560
rect 41492 421502 41939 421504
rect 41873 421499 41939 421502
rect 42517 421154 42583 421157
rect 41492 421152 42583 421154
rect 41492 421096 42522 421152
rect 42578 421096 42583 421152
rect 41492 421094 42583 421096
rect 42517 421091 42583 421094
rect 41781 420746 41847 420749
rect 41492 420744 41847 420746
rect 41492 420688 41786 420744
rect 41842 420688 41847 420744
rect 41492 420686 41847 420688
rect 41781 420683 41847 420686
rect 30422 419900 30482 420308
rect 41781 419522 41847 419525
rect 41492 419520 41847 419522
rect 41492 419464 41786 419520
rect 41842 419464 41847 419520
rect 41492 419462 41847 419464
rect 41781 419459 41847 419462
rect 655053 418026 655119 418029
rect 650164 418024 655119 418026
rect 650164 417968 655058 418024
rect 655114 417968 655119 418024
rect 650164 417966 655119 417968
rect 655053 417963 655119 417966
rect 58433 415442 58499 415445
rect 58433 415440 64492 415442
rect 58433 415384 58438 415440
rect 58494 415384 64492 415440
rect 58433 415382 64492 415384
rect 58433 415379 58499 415382
rect 43621 411498 43687 411501
rect 42934 411496 43687 411498
rect 42934 411440 43626 411496
rect 43682 411440 43687 411496
rect 42934 411438 43687 411440
rect 42793 411270 42859 411273
rect 42934 411270 42994 411438
rect 43621 411435 43687 411438
rect 42793 411268 42994 411270
rect 42793 411212 42798 411268
rect 42854 411212 42994 411268
rect 42793 411210 42994 411212
rect 42793 411207 42859 411210
rect 654869 404698 654935 404701
rect 650164 404696 654935 404698
rect 650164 404640 654874 404696
rect 654930 404640 654935 404696
rect 650164 404638 654935 404640
rect 654869 404635 654935 404638
rect 676262 403749 676322 403852
rect 676213 403744 676322 403749
rect 676213 403688 676218 403744
rect 676274 403688 676322 403744
rect 676213 403686 676322 403688
rect 676213 403683 676279 403686
rect 676262 403341 676322 403444
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 676213 403275 676279 403278
rect 675937 403066 676003 403069
rect 675937 403064 676292 403066
rect 675937 403008 675942 403064
rect 675998 403008 676292 403064
rect 675937 403006 676292 403008
rect 675937 403003 676003 403006
rect 676121 402930 676187 402933
rect 676121 402928 676322 402930
rect 676121 402872 676126 402928
rect 676182 402872 676322 402928
rect 676121 402870 676322 402872
rect 676121 402867 676187 402870
rect 676262 402628 676322 402870
rect 58433 402386 58499 402389
rect 58433 402384 64492 402386
rect 58433 402328 58438 402384
rect 58494 402328 64492 402384
rect 58433 402326 64492 402328
rect 58433 402323 58499 402326
rect 675753 402250 675819 402253
rect 675753 402248 676292 402250
rect 675753 402192 675758 402248
rect 675814 402192 676292 402248
rect 675753 402190 676292 402192
rect 675753 402187 675819 402190
rect 675845 401842 675911 401845
rect 675845 401840 676292 401842
rect 675845 401784 675850 401840
rect 675906 401784 676292 401840
rect 675845 401782 676292 401784
rect 675845 401779 675911 401782
rect 675661 401434 675727 401437
rect 675661 401432 676292 401434
rect 675661 401376 675666 401432
rect 675722 401376 676292 401432
rect 675661 401374 676292 401376
rect 675661 401371 675727 401374
rect 673678 400964 673684 401028
rect 673748 401026 673754 401028
rect 675569 401026 675635 401029
rect 673748 401024 676292 401026
rect 673748 400968 675574 401024
rect 675630 400968 676292 401024
rect 673748 400966 676292 400968
rect 673748 400964 673754 400966
rect 675569 400963 675635 400966
rect 676121 400482 676187 400485
rect 676262 400482 676322 400588
rect 676121 400480 676322 400482
rect 676121 400424 676126 400480
rect 676182 400424 676322 400480
rect 676121 400422 676322 400424
rect 676121 400419 676187 400422
rect 673862 400148 673868 400212
rect 673932 400210 673938 400212
rect 676029 400210 676095 400213
rect 673932 400208 676292 400210
rect 673932 400152 676034 400208
rect 676090 400152 676292 400208
rect 673932 400150 676292 400152
rect 673932 400148 673938 400150
rect 676029 400147 676095 400150
rect 676029 399802 676095 399805
rect 676029 399800 676292 399802
rect 676029 399744 676034 399800
rect 676090 399744 676292 399800
rect 676029 399742 676292 399744
rect 676029 399739 676095 399742
rect 676029 399394 676095 399397
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 676121 398850 676187 398853
rect 676262 398850 676322 398956
rect 676121 398848 676322 398850
rect 676121 398792 676126 398848
rect 676182 398792 676322 398848
rect 676121 398790 676322 398792
rect 676121 398787 676187 398790
rect 675845 398578 675911 398581
rect 675845 398576 676292 398578
rect 675845 398520 675850 398576
rect 675906 398520 676292 398576
rect 675845 398518 676292 398520
rect 675845 398515 675911 398518
rect 676029 398170 676095 398173
rect 676029 398168 676292 398170
rect 676029 398112 676034 398168
rect 676090 398112 676292 398168
rect 676029 398110 676292 398112
rect 676029 398107 676095 398110
rect 675937 397762 676003 397765
rect 675937 397760 676292 397762
rect 675937 397704 675942 397760
rect 675998 397704 676292 397760
rect 675937 397702 676292 397704
rect 675937 397699 676003 397702
rect 676029 397354 676095 397357
rect 676029 397352 676292 397354
rect 676029 397296 676034 397352
rect 676090 397296 676292 397352
rect 676029 397294 676292 397296
rect 676029 397291 676095 397294
rect 675293 396946 675359 396949
rect 675293 396944 676292 396946
rect 675293 396888 675298 396944
rect 675354 396888 676292 396944
rect 675293 396886 676292 396888
rect 675293 396883 675359 396886
rect 676029 396538 676095 396541
rect 676029 396536 676292 396538
rect 676029 396480 676034 396536
rect 676090 396480 676292 396536
rect 676029 396478 676292 396480
rect 676029 396475 676095 396478
rect 676121 395994 676187 395997
rect 676262 395994 676322 396100
rect 676121 395992 676322 395994
rect 676121 395936 676126 395992
rect 676182 395936 676322 395992
rect 676121 395934 676322 395936
rect 676121 395931 676187 395934
rect 675937 395722 676003 395725
rect 675937 395720 676292 395722
rect 675937 395664 675942 395720
rect 675998 395664 676292 395720
rect 675937 395662 676292 395664
rect 675937 395659 676003 395662
rect 675937 395314 676003 395317
rect 675937 395312 676292 395314
rect 675937 395256 675942 395312
rect 675998 395256 676292 395312
rect 675937 395254 676292 395256
rect 675937 395251 676003 395254
rect 676029 394906 676095 394909
rect 676029 394904 676292 394906
rect 676029 394848 676034 394904
rect 676090 394848 676292 394904
rect 676029 394846 676292 394848
rect 676029 394843 676095 394846
rect 676029 394498 676095 394501
rect 676029 394496 676292 394498
rect 676029 394440 676034 394496
rect 676090 394440 676292 394496
rect 676029 394438 676292 394440
rect 676029 394435 676095 394438
rect 676121 393954 676187 393957
rect 676262 393954 676322 394060
rect 676121 393952 676322 393954
rect 676121 393896 676126 393952
rect 676182 393896 676322 393952
rect 676121 393894 676322 393896
rect 676121 393891 676187 393894
rect 679022 393549 679082 393652
rect 679022 393544 679131 393549
rect 679022 393488 679070 393544
rect 679126 393488 679131 393544
rect 679022 393486 679131 393488
rect 679065 393483 679131 393486
rect 684542 392836 684602 393244
rect 679065 392730 679131 392733
rect 679022 392728 679131 392730
rect 679022 392672 679070 392728
rect 679126 392672 679131 392728
rect 679022 392667 679131 392672
rect 679022 392428 679082 392667
rect 654317 391506 654383 391509
rect 650164 391504 654383 391506
rect 650164 391448 654322 391504
rect 654378 391448 654383 391504
rect 650164 391446 654383 391448
rect 654317 391443 654383 391446
rect 57973 389330 58039 389333
rect 57973 389328 64492 389330
rect 57973 389272 57978 389328
rect 58034 389272 64492 389328
rect 57973 389270 64492 389272
rect 57973 389267 58039 389270
rect 40166 388996 40172 389060
rect 40236 389058 40242 389060
rect 41137 389058 41203 389061
rect 40236 389056 41203 389058
rect 40236 389000 41142 389056
rect 41198 389000 41203 389056
rect 40236 388998 41203 389000
rect 40236 388996 40242 388998
rect 41137 388995 41203 388998
rect 41505 387970 41571 387973
rect 41462 387968 41571 387970
rect 41462 387912 41510 387968
rect 41566 387912 41571 387968
rect 41462 387907 41571 387912
rect 41462 387668 41522 387907
rect 41505 387562 41571 387565
rect 41462 387560 41571 387562
rect 41462 387504 41510 387560
rect 41566 387504 41571 387560
rect 41462 387499 41571 387504
rect 41462 387260 41522 387499
rect 41505 387154 41571 387157
rect 41462 387152 41571 387154
rect 41462 387096 41510 387152
rect 41566 387096 41571 387152
rect 41462 387091 41571 387096
rect 41462 386852 41522 387091
rect 41137 386746 41203 386749
rect 63217 386746 63283 386749
rect 41137 386744 63283 386746
rect 41137 386688 41142 386744
rect 41198 386688 63222 386744
rect 63278 386688 63283 386744
rect 41137 386686 63283 386688
rect 41137 386683 41203 386686
rect 63217 386683 63283 386686
rect 41462 386338 41522 386444
rect 42926 386338 42932 386340
rect 41462 386278 42932 386338
rect 42926 386276 42932 386278
rect 42996 386338 43002 386340
rect 62113 386338 62179 386341
rect 42996 386336 62179 386338
rect 42996 386280 62118 386336
rect 62174 386280 62179 386336
rect 42996 386278 62179 386280
rect 42996 386276 43002 386278
rect 62113 386275 62179 386278
rect 42793 386066 42859 386069
rect 41492 386064 42859 386066
rect 41492 386008 42798 386064
rect 42854 386008 42859 386064
rect 41492 386006 42859 386008
rect 42793 386003 42859 386006
rect 43805 385658 43871 385661
rect 41492 385656 43871 385658
rect 41492 385600 43810 385656
rect 43866 385600 43871 385656
rect 41492 385598 43871 385600
rect 43805 385595 43871 385598
rect 43529 385250 43595 385253
rect 41492 385248 43595 385250
rect 41492 385192 43534 385248
rect 43590 385192 43595 385248
rect 41492 385190 43595 385192
rect 43529 385187 43595 385190
rect 41137 384706 41203 384709
rect 41278 384708 41338 384812
rect 41094 384704 41203 384706
rect 41094 384648 41142 384704
rect 41198 384648 41203 384704
rect 41094 384643 41203 384648
rect 41270 384644 41276 384708
rect 41340 384644 41346 384708
rect 41094 384404 41154 384643
rect 42742 384026 42748 384028
rect 41492 383966 42748 384026
rect 42742 383964 42748 383966
rect 42812 383964 42818 384028
rect 39982 383828 39988 383892
rect 40052 383890 40058 383892
rect 40052 383830 40234 383890
rect 40052 383828 40058 383830
rect 40174 383618 40234 383830
rect 63309 383754 63375 383757
rect 41830 383752 63375 383754
rect 41830 383696 63314 383752
rect 63370 383696 63375 383752
rect 41830 383694 63375 383696
rect 41830 383618 41890 383694
rect 63309 383691 63375 383694
rect 40174 383588 41890 383618
rect 40204 383558 41890 383588
rect 42742 383420 42748 383484
rect 42812 383482 42818 383484
rect 62205 383482 62271 383485
rect 42812 383480 62271 383482
rect 42812 383424 62210 383480
rect 62266 383424 62271 383480
rect 42812 383422 62271 383424
rect 42812 383420 42818 383422
rect 62205 383419 62271 383422
rect 43345 383210 43411 383213
rect 41492 383208 43411 383210
rect 41492 383152 43350 383208
rect 43406 383152 43411 383208
rect 41492 383150 43411 383152
rect 43345 383147 43411 383150
rect 39982 383012 39988 383076
rect 40052 383074 40058 383076
rect 41270 383074 41276 383076
rect 40052 383014 41276 383074
rect 40052 383012 40058 383014
rect 41270 383012 41276 383014
rect 41340 383074 41346 383076
rect 62021 383074 62087 383077
rect 41340 383072 62087 383074
rect 41340 383016 62026 383072
rect 62082 383016 62087 383072
rect 41340 383014 62087 383016
rect 41340 383012 41346 383014
rect 62021 383011 62087 383014
rect 42793 382802 42859 382805
rect 41492 382800 42859 382802
rect 41492 382744 42798 382800
rect 42854 382744 42859 382800
rect 41492 382742 42859 382744
rect 42793 382739 42859 382742
rect 41462 382260 41522 382364
rect 41454 382196 41460 382260
rect 41524 382196 41530 382260
rect 42977 381986 43043 381989
rect 41492 381984 43043 381986
rect 41492 381928 42982 381984
rect 43038 381928 43043 381984
rect 41492 381926 43043 381928
rect 42977 381923 43043 381926
rect 43897 381578 43963 381581
rect 41492 381576 43963 381578
rect 41492 381520 43902 381576
rect 43958 381520 43963 381576
rect 41492 381518 43963 381520
rect 43897 381515 43963 381518
rect 42333 381170 42399 381173
rect 41492 381168 42399 381170
rect 41492 381112 42338 381168
rect 42394 381112 42399 381168
rect 41492 381110 42399 381112
rect 42333 381107 42399 381110
rect 43437 380762 43503 380765
rect 41492 380760 43503 380762
rect 41492 380704 43442 380760
rect 43498 380704 43503 380760
rect 41492 380702 43503 380704
rect 43437 380699 43503 380702
rect 43621 380354 43687 380357
rect 41492 380352 43687 380354
rect 41492 380296 43626 380352
rect 43682 380296 43687 380352
rect 41492 380294 43687 380296
rect 43621 380291 43687 380294
rect 43713 379946 43779 379949
rect 41492 379944 43779 379946
rect 41492 379888 43718 379944
rect 43774 379888 43779 379944
rect 41492 379886 43779 379888
rect 43713 379883 43779 379886
rect 42885 379538 42951 379541
rect 41492 379536 42951 379538
rect 41492 379480 42890 379536
rect 42946 379480 42951 379536
rect 41492 379478 42951 379480
rect 42885 379475 42951 379478
rect 43161 379130 43227 379133
rect 41492 379128 43227 379130
rect 41492 379072 43166 379128
rect 43222 379072 43227 379128
rect 41492 379070 43227 379072
rect 43161 379067 43227 379070
rect 43253 378722 43319 378725
rect 41492 378720 43319 378722
rect 41492 378664 43258 378720
rect 43314 378664 43319 378720
rect 41492 378662 43319 378664
rect 43253 378659 43319 378662
rect 43069 378314 43135 378317
rect 41492 378312 43135 378314
rect 41492 378256 43074 378312
rect 43130 378256 43135 378312
rect 41492 378254 43135 378256
rect 43069 378251 43135 378254
rect 656801 378178 656867 378181
rect 650164 378176 656867 378178
rect 650164 378120 656806 378176
rect 656862 378120 656867 378176
rect 650164 378118 656867 378120
rect 656801 378115 656867 378118
rect 41462 377773 41522 377876
rect 41462 377768 41571 377773
rect 41462 377712 41510 377768
rect 41566 377712 41571 377768
rect 41462 377710 41571 377712
rect 41505 377707 41571 377710
rect 41462 377362 41522 377468
rect 41597 377362 41663 377365
rect 41462 377360 41663 377362
rect 41462 377304 41602 377360
rect 41658 377304 41663 377360
rect 41462 377302 41663 377304
rect 41597 377299 41663 377302
rect 30422 376652 30482 377060
rect 58433 376274 58499 376277
rect 58433 376272 64492 376274
rect 41462 376138 41522 376244
rect 58433 376216 58438 376272
rect 58494 376216 64492 376272
rect 58433 376214 64492 376216
rect 58433 376211 58499 376214
rect 41597 376138 41663 376141
rect 41462 376136 41663 376138
rect 41462 376080 41602 376136
rect 41658 376080 41663 376136
rect 41462 376078 41663 376080
rect 41597 376075 41663 376078
rect 656801 364850 656867 364853
rect 650164 364848 656867 364850
rect 650164 364792 656806 364848
rect 656862 364792 656867 364848
rect 650164 364790 656867 364792
rect 656801 364787 656867 364790
rect 58433 363354 58499 363357
rect 58433 363352 64492 363354
rect 58433 363296 58438 363352
rect 58494 363296 64492 363352
rect 58433 363294 64492 363296
rect 58433 363291 58499 363294
rect 675845 358730 675911 358733
rect 675845 358728 676292 358730
rect 675845 358672 675850 358728
rect 675906 358672 676292 358728
rect 675845 358670 676292 358672
rect 675845 358667 675911 358670
rect 675937 358322 676003 358325
rect 675937 358320 676292 358322
rect 675937 358264 675942 358320
rect 675998 358264 676292 358320
rect 675937 358262 676292 358264
rect 675937 358259 676003 358262
rect 676029 357914 676095 357917
rect 676029 357912 676292 357914
rect 676029 357856 676034 357912
rect 676090 357856 676292 357912
rect 676029 357854 676292 357856
rect 676029 357851 676095 357854
rect 674046 357444 674052 357508
rect 674116 357506 674122 357508
rect 675753 357506 675819 357509
rect 674116 357504 676292 357506
rect 674116 357448 675758 357504
rect 675814 357448 676292 357504
rect 674116 357446 676292 357448
rect 674116 357444 674122 357446
rect 675753 357443 675819 357446
rect 675753 357098 675819 357101
rect 675753 357096 676292 357098
rect 675753 357040 675758 357096
rect 675814 357040 676292 357096
rect 675753 357038 676292 357040
rect 675753 357035 675819 357038
rect 675661 356690 675727 356693
rect 675661 356688 676292 356690
rect 675661 356632 675666 356688
rect 675722 356632 676292 356688
rect 675661 356630 676292 356632
rect 675661 356627 675727 356630
rect 676029 356282 676095 356285
rect 676029 356280 676292 356282
rect 676029 356224 676034 356280
rect 676090 356224 676292 356280
rect 676029 356222 676292 356224
rect 676029 356219 676095 356222
rect 674230 355812 674236 355876
rect 674300 355874 674306 355876
rect 675293 355874 675359 355877
rect 674300 355872 676292 355874
rect 674300 355816 675298 355872
rect 675354 355816 676292 355872
rect 674300 355814 676292 355816
rect 674300 355812 674306 355814
rect 675293 355811 675359 355814
rect 41454 355676 41460 355740
rect 41524 355738 41530 355740
rect 41781 355738 41847 355741
rect 41524 355736 41847 355738
rect 41524 355680 41786 355736
rect 41842 355680 41847 355736
rect 41524 355678 41847 355680
rect 41524 355676 41530 355678
rect 41781 355675 41847 355678
rect 676029 355466 676095 355469
rect 676029 355464 676292 355466
rect 676029 355408 676034 355464
rect 676090 355408 676292 355464
rect 676029 355406 676292 355408
rect 676029 355403 676095 355406
rect 674414 354996 674420 355060
rect 674484 355058 674490 355060
rect 674741 355058 674807 355061
rect 674484 355056 676292 355058
rect 674484 355000 674746 355056
rect 674802 355000 676292 355056
rect 674484 354998 676292 355000
rect 674484 354996 674490 354998
rect 674741 354995 674807 354998
rect 676029 354650 676095 354653
rect 676029 354648 676292 354650
rect 676029 354592 676034 354648
rect 676090 354592 676292 354648
rect 676029 354590 676292 354592
rect 676029 354587 676095 354590
rect 676029 354242 676095 354245
rect 676029 354240 676292 354242
rect 676029 354184 676034 354240
rect 676090 354184 676292 354240
rect 676029 354182 676292 354184
rect 676029 354179 676095 354182
rect 676078 353774 676292 353834
rect 676078 353700 676138 353774
rect 676070 353636 676076 353700
rect 676140 353636 676146 353700
rect 676029 353426 676095 353429
rect 676029 353424 676292 353426
rect 676029 353368 676034 353424
rect 676090 353368 676292 353424
rect 676029 353366 676292 353368
rect 676029 353363 676095 353366
rect 676029 353018 676095 353021
rect 676029 353016 676292 353018
rect 676029 352960 676034 353016
rect 676090 352960 676292 353016
rect 676029 352958 676292 352960
rect 676029 352955 676095 352958
rect 675937 352610 676003 352613
rect 675937 352608 676292 352610
rect 675937 352552 675942 352608
rect 675998 352552 676292 352608
rect 675937 352550 676292 352552
rect 675937 352547 676003 352550
rect 675886 352140 675892 352204
rect 675956 352202 675962 352204
rect 675956 352142 676292 352202
rect 675956 352140 675962 352142
rect 33041 351930 33107 351933
rect 42926 351930 42932 351932
rect 33041 351928 42932 351930
rect 33041 351872 33046 351928
rect 33102 351872 42932 351928
rect 33041 351870 42932 351872
rect 33041 351867 33107 351870
rect 42926 351868 42932 351870
rect 42996 351868 43002 351932
rect 675293 351794 675359 351797
rect 675293 351792 676292 351794
rect 675293 351736 675298 351792
rect 675354 351736 676292 351792
rect 675293 351734 676292 351736
rect 675293 351731 675359 351734
rect 654869 351658 654935 351661
rect 650164 351656 654935 351658
rect 650164 351600 654874 351656
rect 654930 351600 654935 351656
rect 650164 351598 654935 351600
rect 654869 351595 654935 351598
rect 676029 351386 676095 351389
rect 676029 351384 676292 351386
rect 676029 351328 676034 351384
rect 676090 351328 676292 351384
rect 676029 351326 676292 351328
rect 676029 351323 676095 351326
rect 675937 350978 676003 350981
rect 675937 350976 676292 350978
rect 675937 350920 675942 350976
rect 675998 350920 676292 350976
rect 675937 350918 676292 350920
rect 675937 350915 676003 350918
rect 675702 350508 675708 350572
rect 675772 350570 675778 350572
rect 675772 350510 676292 350570
rect 675772 350508 675778 350510
rect 58433 350298 58499 350301
rect 58433 350296 64492 350298
rect 58433 350240 58438 350296
rect 58494 350240 64492 350296
rect 58433 350238 64492 350240
rect 58433 350235 58499 350238
rect 676029 350162 676095 350165
rect 676029 350160 676292 350162
rect 676029 350104 676034 350160
rect 676090 350104 676292 350160
rect 676029 350102 676292 350104
rect 676029 350099 676095 350102
rect 676029 349754 676095 349757
rect 676029 349752 676292 349754
rect 676029 349696 676034 349752
rect 676090 349696 676292 349752
rect 676029 349694 676292 349696
rect 676029 349691 676095 349694
rect 675937 349346 676003 349349
rect 675937 349344 676292 349346
rect 675937 349288 675942 349344
rect 675998 349288 676292 349344
rect 675937 349286 676292 349288
rect 675937 349283 676003 349286
rect 675937 348938 676003 348941
rect 675937 348936 676292 348938
rect 675937 348880 675942 348936
rect 675998 348880 676292 348936
rect 675937 348878 676292 348880
rect 675937 348875 676003 348878
rect 676078 348470 676292 348530
rect 676078 347309 676138 348470
rect 679022 347684 679082 348092
rect 676029 347306 676138 347309
rect 675948 347304 676292 347306
rect 675948 347248 676034 347304
rect 676090 347248 676292 347304
rect 675948 347246 676292 347248
rect 676029 347243 676095 347246
rect 41781 344586 41847 344589
rect 41492 344584 41847 344586
rect 41492 344528 41786 344584
rect 41842 344528 41847 344584
rect 41492 344526 41847 344528
rect 41781 344523 41847 344526
rect 41597 344314 41663 344317
rect 41462 344312 41663 344314
rect 41462 344256 41602 344312
rect 41658 344256 41663 344312
rect 41462 344254 41663 344256
rect 41462 344148 41522 344254
rect 41597 344251 41663 344254
rect 41597 343906 41663 343909
rect 41462 343904 41663 343906
rect 41462 343848 41602 343904
rect 41658 343848 41663 343904
rect 41462 343846 41663 343848
rect 41462 343740 41522 343846
rect 41597 343843 41663 343846
rect 41781 343362 41847 343365
rect 41492 343360 41847 343362
rect 41492 343304 41786 343360
rect 41842 343304 41847 343360
rect 41492 343302 41847 343304
rect 41781 343299 41847 343302
rect 33041 343090 33107 343093
rect 32998 343088 33107 343090
rect 32998 343032 33046 343088
rect 33102 343032 33107 343088
rect 32998 343027 33107 343032
rect 32998 342924 33058 343027
rect 41505 342682 41571 342685
rect 41462 342680 41571 342682
rect 41462 342624 41510 342680
rect 41566 342624 41571 342680
rect 41462 342619 41571 342624
rect 41462 342516 41522 342619
rect 43253 342138 43319 342141
rect 41492 342136 43319 342138
rect 41492 342080 43258 342136
rect 43314 342080 43319 342136
rect 41492 342078 43319 342080
rect 43253 342075 43319 342078
rect 44265 341730 44331 341733
rect 41492 341728 44331 341730
rect 41492 341672 44270 341728
rect 44326 341672 44331 341728
rect 41492 341670 44331 341672
rect 44265 341667 44331 341670
rect 39982 341396 39988 341460
rect 40052 341396 40058 341460
rect 39990 341292 40050 341396
rect 44357 340914 44423 340917
rect 41492 340912 44423 340914
rect 41492 340856 44362 340912
rect 44418 340856 44423 340912
rect 41492 340854 44423 340856
rect 44357 340851 44423 340854
rect 42742 340506 42748 340508
rect 41492 340446 42748 340506
rect 42742 340444 42748 340446
rect 42812 340444 42818 340508
rect 41822 340098 41828 340100
rect 41492 340038 41828 340098
rect 41822 340036 41828 340038
rect 41892 340036 41898 340100
rect 44265 339962 44331 339965
rect 46197 339962 46263 339965
rect 44265 339960 46263 339962
rect 44265 339904 44270 339960
rect 44326 339904 46202 339960
rect 46258 339904 46263 339960
rect 44265 339902 46263 339904
rect 44265 339899 44331 339902
rect 46197 339899 46263 339902
rect 32673 339826 32739 339829
rect 32630 339824 32739 339826
rect 32630 339768 32678 339824
rect 32734 339768 32739 339824
rect 32630 339763 32739 339768
rect 32630 339660 32690 339763
rect 44357 339554 44423 339557
rect 46381 339554 46447 339557
rect 44357 339552 46447 339554
rect 44357 339496 44362 339552
rect 44418 339496 46386 339552
rect 46442 339496 46447 339552
rect 44357 339494 46447 339496
rect 44357 339491 44423 339494
rect 46381 339491 46447 339494
rect 42558 339282 42564 339284
rect 41492 339222 42564 339282
rect 42558 339220 42564 339222
rect 42628 339220 42634 339284
rect 42006 338874 42012 338876
rect 41492 338814 42012 338874
rect 42006 338812 42012 338814
rect 42076 338812 42082 338876
rect 32814 338197 32874 338436
rect 655053 338330 655119 338333
rect 650164 338328 655119 338330
rect 650164 338272 655058 338328
rect 655114 338272 655119 338328
rect 650164 338270 655119 338272
rect 655053 338267 655119 338270
rect 32765 338192 32874 338197
rect 32765 338136 32770 338192
rect 32826 338136 32874 338192
rect 32765 338134 32874 338136
rect 32765 338131 32831 338134
rect 32998 337789 33058 338028
rect 32998 337784 33107 337789
rect 32998 337728 33046 337784
rect 33102 337728 33107 337784
rect 32998 337726 33107 337728
rect 33041 337723 33107 337726
rect 41462 337378 41522 337620
rect 41638 337378 41644 337380
rect 41462 337318 41644 337378
rect 41638 337316 41644 337318
rect 41708 337316 41714 337380
rect 42190 337242 42196 337244
rect 41492 337182 42196 337242
rect 42190 337180 42196 337182
rect 42260 337180 42266 337244
rect 58433 337242 58499 337245
rect 58433 337240 64492 337242
rect 58433 337184 58438 337240
rect 58494 337184 64492 337240
rect 58433 337182 64492 337184
rect 58433 337179 58499 337182
rect 42374 336834 42380 336836
rect 41492 336774 42380 336834
rect 42374 336772 42380 336774
rect 42444 336772 42450 336836
rect 32814 336157 32874 336396
rect 32814 336152 32923 336157
rect 32814 336096 32862 336152
rect 32918 336096 32923 336152
rect 32814 336094 32923 336096
rect 32857 336091 32923 336094
rect 32998 335749 33058 335988
rect 32949 335744 33058 335749
rect 32949 335688 32954 335744
rect 33010 335688 33058 335744
rect 32949 335686 33058 335688
rect 32949 335683 33015 335686
rect 43069 335610 43135 335613
rect 41492 335608 43135 335610
rect 41492 335552 43074 335608
rect 43130 335552 43135 335608
rect 41492 335550 43135 335552
rect 43069 335547 43135 335550
rect 42977 335202 43043 335205
rect 41492 335200 43043 335202
rect 41492 335144 42982 335200
rect 43038 335144 43043 335200
rect 41492 335142 43043 335144
rect 42977 335139 43043 335142
rect 43161 334794 43227 334797
rect 41492 334792 43227 334794
rect 41492 334736 43166 334792
rect 43222 334736 43227 334792
rect 41492 334734 43227 334736
rect 43161 334731 43227 334734
rect 41462 334117 41522 334356
rect 41462 334112 41571 334117
rect 41462 334056 41510 334112
rect 41566 334056 41571 334112
rect 41462 334054 41571 334056
rect 41505 334051 41571 334054
rect 30422 333540 30482 333948
rect 41462 332893 41522 333132
rect 41462 332888 41571 332893
rect 41462 332832 41510 332888
rect 41566 332832 41571 332888
rect 41462 332830 41571 332832
rect 41505 332827 41571 332830
rect 675661 330580 675727 330581
rect 675661 330576 675708 330580
rect 675772 330578 675778 330580
rect 675661 330520 675666 330576
rect 675661 330516 675708 330520
rect 675772 330518 675818 330578
rect 675772 330516 675778 330518
rect 675661 330515 675727 330516
rect 32765 329762 32831 329765
rect 41454 329762 41460 329764
rect 32765 329760 41460 329762
rect 32765 329704 32770 329760
rect 32826 329704 41460 329760
rect 32765 329702 41460 329704
rect 32765 329699 32831 329702
rect 41454 329700 41460 329702
rect 41524 329700 41530 329764
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 675753 326906 675819 326909
rect 675886 326906 675892 326908
rect 675753 326904 675892 326906
rect 675753 326848 675758 326904
rect 675814 326848 675892 326904
rect 675753 326846 675892 326848
rect 675753 326843 675819 326846
rect 675886 326844 675892 326846
rect 675956 326844 675962 326908
rect 654869 325002 654935 325005
rect 650164 325000 654935 325002
rect 650164 324944 654874 325000
rect 654930 324944 654935 325000
rect 650164 324942 654935 324944
rect 654869 324939 654935 324942
rect 58157 324186 58223 324189
rect 58157 324184 64492 324186
rect 58157 324128 58162 324184
rect 58218 324128 64492 324184
rect 58157 324126 64492 324128
rect 58157 324123 58223 324126
rect 41454 319908 41460 319972
rect 41524 319970 41530 319972
rect 41781 319970 41847 319973
rect 41524 319968 41847 319970
rect 41524 319912 41786 319968
rect 41842 319912 41847 319968
rect 41524 319910 41847 319912
rect 41524 319908 41530 319910
rect 41781 319907 41847 319910
rect 42149 316978 42215 316981
rect 42374 316978 42380 316980
rect 42149 316976 42380 316978
rect 42149 316920 42154 316976
rect 42210 316920 42380 316976
rect 42149 316918 42380 316920
rect 42149 316915 42215 316918
rect 42374 316916 42380 316918
rect 42444 316916 42450 316980
rect 42149 316300 42215 316301
rect 42149 316298 42196 316300
rect 42104 316296 42196 316298
rect 42104 316240 42154 316296
rect 42104 316238 42196 316240
rect 42149 316236 42196 316238
rect 42260 316236 42266 316300
rect 42149 316235 42215 316236
rect 41965 315620 42031 315621
rect 41965 315616 42012 315620
rect 42076 315618 42082 315620
rect 41965 315560 41970 315616
rect 41965 315556 42012 315560
rect 42076 315558 42122 315618
rect 42076 315556 42082 315558
rect 41965 315555 42031 315556
rect 41873 313852 41939 313853
rect 41822 313850 41828 313852
rect 41782 313790 41828 313850
rect 41892 313848 41939 313852
rect 41934 313792 41939 313848
rect 41822 313788 41828 313790
rect 41892 313788 41939 313792
rect 41873 313787 41939 313788
rect 676029 313714 676095 313717
rect 676029 313712 676292 313714
rect 676029 313656 676034 313712
rect 676090 313656 676292 313712
rect 676029 313654 676292 313656
rect 676029 313651 676095 313654
rect 676262 313173 676322 313276
rect 676213 313168 676322 313173
rect 676213 313112 676218 313168
rect 676274 313112 676322 313168
rect 676213 313110 676322 313112
rect 676213 313107 676279 313110
rect 41638 312972 41644 313036
rect 41708 313034 41714 313036
rect 41781 313034 41847 313037
rect 41708 313032 41847 313034
rect 41708 312976 41786 313032
rect 41842 312976 41847 313032
rect 41708 312974 41847 312976
rect 41708 312972 41714 312974
rect 41781 312971 41847 312974
rect 676029 312898 676095 312901
rect 676029 312896 676292 312898
rect 676029 312840 676034 312896
rect 676090 312840 676292 312896
rect 676029 312838 676292 312840
rect 676029 312835 676095 312838
rect 676029 312490 676095 312493
rect 676029 312488 676292 312490
rect 676029 312432 676034 312488
rect 676090 312432 676292 312488
rect 676029 312430 676292 312432
rect 676029 312427 676095 312430
rect 42149 312354 42215 312357
rect 42558 312354 42564 312356
rect 42149 312352 42564 312354
rect 42149 312296 42154 312352
rect 42210 312296 42564 312352
rect 42149 312294 42564 312296
rect 42149 312291 42215 312294
rect 42558 312292 42564 312294
rect 42628 312292 42634 312356
rect 676029 312082 676095 312085
rect 676029 312080 676292 312082
rect 676029 312024 676034 312080
rect 676090 312024 676292 312080
rect 676029 312022 676292 312024
rect 676029 312019 676095 312022
rect 654133 311810 654199 311813
rect 650164 311808 654199 311810
rect 650164 311752 654138 311808
rect 654194 311752 654199 311808
rect 650164 311750 654199 311752
rect 654133 311747 654199 311750
rect 676029 311674 676095 311677
rect 676029 311672 676292 311674
rect 676029 311616 676034 311672
rect 676090 311616 676292 311672
rect 676029 311614 676292 311616
rect 676029 311611 676095 311614
rect 676029 311266 676095 311269
rect 676029 311264 676292 311266
rect 676029 311208 676034 311264
rect 676090 311208 676292 311264
rect 676029 311206 676292 311208
rect 676029 311203 676095 311206
rect 59261 311130 59327 311133
rect 59261 311128 64492 311130
rect 59261 311072 59266 311128
rect 59322 311072 64492 311128
rect 59261 311070 64492 311072
rect 59261 311067 59327 311070
rect 676029 310858 676095 310861
rect 676029 310856 676292 310858
rect 676029 310800 676034 310856
rect 676090 310800 676292 310856
rect 676029 310798 676292 310800
rect 676029 310795 676095 310798
rect 676029 310450 676095 310453
rect 676029 310448 676292 310450
rect 676029 310392 676034 310448
rect 676090 310392 676292 310448
rect 676029 310390 676292 310392
rect 676029 310387 676095 310390
rect 676029 310042 676095 310045
rect 676029 310040 676292 310042
rect 676029 309984 676034 310040
rect 676090 309984 676292 310040
rect 676029 309982 676292 309984
rect 676029 309979 676095 309982
rect 676029 309634 676095 309637
rect 676029 309632 676292 309634
rect 676029 309576 676034 309632
rect 676090 309576 676292 309632
rect 676029 309574 676292 309576
rect 676029 309571 676095 309574
rect 676029 309226 676095 309229
rect 676029 309224 676292 309226
rect 676029 309168 676034 309224
rect 676090 309168 676292 309224
rect 676029 309166 676292 309168
rect 676029 309163 676095 309166
rect 676029 308818 676095 308821
rect 676029 308816 676292 308818
rect 676029 308760 676034 308816
rect 676090 308760 676292 308816
rect 676029 308758 676292 308760
rect 676029 308755 676095 308758
rect 675753 308410 675819 308413
rect 675753 308408 676292 308410
rect 675753 308352 675758 308408
rect 675814 308352 676292 308408
rect 675753 308350 676292 308352
rect 675753 308347 675819 308350
rect 676029 308002 676095 308005
rect 676029 308000 676292 308002
rect 676029 307944 676034 308000
rect 676090 307944 676292 308000
rect 676029 307942 676292 307944
rect 676029 307939 676095 307942
rect 676121 307458 676187 307461
rect 676262 307458 676322 307564
rect 676121 307456 676322 307458
rect 676121 307400 676126 307456
rect 676182 307400 676322 307456
rect 676121 307398 676322 307400
rect 676121 307395 676187 307398
rect 675937 307186 676003 307189
rect 675937 307184 676292 307186
rect 675937 307128 675942 307184
rect 675998 307128 676292 307184
rect 675937 307126 676292 307128
rect 675937 307123 676003 307126
rect 675477 306778 675543 306781
rect 675477 306776 676292 306778
rect 675477 306720 675482 306776
rect 675538 306720 676292 306776
rect 675477 306718 676292 306720
rect 675477 306715 675543 306718
rect 676029 306370 676095 306373
rect 676029 306368 676292 306370
rect 676029 306312 676034 306368
rect 676090 306312 676292 306368
rect 676029 306310 676292 306312
rect 676029 306307 676095 306310
rect 675886 305900 675892 305964
rect 675956 305962 675962 305964
rect 675956 305902 676292 305962
rect 675956 305900 675962 305902
rect 676121 305418 676187 305421
rect 676262 305418 676322 305524
rect 676121 305416 676322 305418
rect 676121 305360 676126 305416
rect 676182 305360 676322 305416
rect 676121 305358 676322 305360
rect 676121 305355 676187 305358
rect 676121 305010 676187 305013
rect 676262 305010 676322 305116
rect 676121 305008 676322 305010
rect 676121 304952 676126 305008
rect 676182 304952 676322 305008
rect 676121 304950 676322 304952
rect 676121 304947 676187 304950
rect 676121 304602 676187 304605
rect 676262 304602 676322 304708
rect 676121 304600 676322 304602
rect 676121 304544 676126 304600
rect 676182 304544 676322 304600
rect 676121 304542 676322 304544
rect 676121 304539 676187 304542
rect 675937 304330 676003 304333
rect 675937 304328 676292 304330
rect 675937 304272 675942 304328
rect 675998 304272 676292 304328
rect 675937 304270 676292 304272
rect 675937 304267 676003 304270
rect 675845 303922 675911 303925
rect 675845 303920 676292 303922
rect 675845 303864 675850 303920
rect 675906 303864 676292 303920
rect 675845 303862 676292 303864
rect 675845 303859 675911 303862
rect 679022 303381 679082 303484
rect 678973 303376 679082 303381
rect 678973 303320 678978 303376
rect 679034 303320 679082 303376
rect 678973 303318 679082 303320
rect 678973 303315 679039 303318
rect 684542 302668 684602 303076
rect 678973 302562 679039 302565
rect 678973 302560 679082 302562
rect 678973 302504 678978 302560
rect 679034 302504 679082 302560
rect 678973 302499 679082 302504
rect 679022 302260 679082 302499
rect 41505 301610 41571 301613
rect 41462 301608 41571 301610
rect 41462 301552 41510 301608
rect 41566 301552 41571 301608
rect 41462 301547 41571 301552
rect 41462 301308 41522 301547
rect 41781 300930 41847 300933
rect 41492 300928 41847 300930
rect 41492 300872 41786 300928
rect 41842 300872 41847 300928
rect 41492 300870 41847 300872
rect 41781 300867 41847 300870
rect 53833 300522 53899 300525
rect 41492 300520 53899 300522
rect 41492 300464 53838 300520
rect 53894 300464 53899 300520
rect 41492 300462 53899 300464
rect 53833 300459 53899 300462
rect 42374 300114 42380 300116
rect 41492 300054 42380 300114
rect 42374 300052 42380 300054
rect 42444 300114 42450 300116
rect 48313 300114 48379 300117
rect 42444 300112 48379 300114
rect 42444 300056 48318 300112
rect 48374 300056 48379 300112
rect 42444 300054 48379 300056
rect 42444 300052 42450 300054
rect 48313 300051 48379 300054
rect 44173 299706 44239 299709
rect 41492 299704 44239 299706
rect 41492 299648 44178 299704
rect 44234 299648 44239 299704
rect 41492 299646 44239 299648
rect 44173 299643 44239 299646
rect 43069 299298 43135 299301
rect 41492 299296 43135 299298
rect 41492 299240 43074 299296
rect 43130 299240 43135 299296
rect 41492 299238 43135 299240
rect 43069 299235 43135 299238
rect 43437 298890 43503 298893
rect 41492 298888 43503 298890
rect 41492 298832 43442 298888
rect 43498 298832 43503 298888
rect 41492 298830 43503 298832
rect 43437 298827 43503 298830
rect 41822 298482 41828 298484
rect 41492 298422 41828 298482
rect 41822 298420 41828 298422
rect 41892 298482 41898 298484
rect 46105 298482 46171 298485
rect 655605 298482 655671 298485
rect 41892 298480 46171 298482
rect 41892 298424 46110 298480
rect 46166 298424 46171 298480
rect 41892 298422 46171 298424
rect 650164 298480 655671 298482
rect 650164 298424 655610 298480
rect 655666 298424 655671 298480
rect 650164 298422 655671 298424
rect 41892 298420 41898 298422
rect 46105 298419 46171 298422
rect 655605 298419 655671 298422
rect 59353 298210 59419 298213
rect 59353 298208 64492 298210
rect 59353 298152 59358 298208
rect 59414 298152 64492 298208
rect 59353 298150 64492 298152
rect 59353 298147 59419 298150
rect 44265 298074 44331 298077
rect 41492 298072 44331 298074
rect 41492 298016 44270 298072
rect 44326 298016 44331 298072
rect 41492 298014 44331 298016
rect 44265 298011 44331 298014
rect 42190 297666 42196 297668
rect 41492 297606 42196 297666
rect 42190 297604 42196 297606
rect 42260 297666 42266 297668
rect 48221 297666 48287 297669
rect 42260 297664 48287 297666
rect 42260 297608 48226 297664
rect 48282 297608 48287 297664
rect 42260 297606 48287 297608
rect 42260 297604 42266 297606
rect 48221 297603 48287 297606
rect 44357 297258 44423 297261
rect 41492 297256 44423 297258
rect 41492 297200 44362 297256
rect 44418 297200 44423 297256
rect 41492 297198 44423 297200
rect 44357 297195 44423 297198
rect 32581 296850 32647 296853
rect 32581 296848 32660 296850
rect 32581 296792 32586 296848
rect 32642 296792 32660 296848
rect 32581 296790 32660 296792
rect 32581 296787 32647 296790
rect 32673 296442 32739 296445
rect 32660 296440 32739 296442
rect 32660 296384 32678 296440
rect 32734 296384 32739 296440
rect 32660 296382 32739 296384
rect 32673 296379 32739 296382
rect 32949 296034 33015 296037
rect 32949 296032 33028 296034
rect 32949 295976 32954 296032
rect 33010 295976 33028 296032
rect 32949 295974 33028 295976
rect 32949 295971 33015 295974
rect 42006 295626 42012 295628
rect 41492 295566 42012 295626
rect 42006 295564 42012 295566
rect 42076 295564 42082 295628
rect 41822 295292 41828 295356
rect 41892 295354 41898 295356
rect 42190 295354 42196 295356
rect 41892 295294 42196 295354
rect 41892 295292 41898 295294
rect 42190 295292 42196 295294
rect 42260 295292 42266 295356
rect 32857 295218 32923 295221
rect 32844 295216 32923 295218
rect 32844 295160 32862 295216
rect 32918 295160 32923 295216
rect 32844 295158 32923 295160
rect 32857 295155 32923 295158
rect 41873 294810 41939 294813
rect 41492 294808 41939 294810
rect 41492 294752 41878 294808
rect 41934 294752 41939 294808
rect 41492 294750 41939 294752
rect 41873 294747 41939 294750
rect 33041 294402 33107 294405
rect 33028 294400 33107 294402
rect 33028 294344 33046 294400
rect 33102 294344 33107 294400
rect 33028 294342 33107 294344
rect 33041 294339 33107 294342
rect 41781 293994 41847 293997
rect 41492 293992 41847 293994
rect 41492 293936 41786 293992
rect 41842 293936 41847 293992
rect 41492 293934 41847 293936
rect 41781 293931 41847 293934
rect 42425 293586 42491 293589
rect 41492 293584 42491 293586
rect 41492 293528 42430 293584
rect 42486 293528 42491 293584
rect 41492 293526 42491 293528
rect 42425 293523 42491 293526
rect 43069 293178 43135 293181
rect 41492 293176 43135 293178
rect 41492 293120 43074 293176
rect 43130 293120 43135 293176
rect 41492 293118 43135 293120
rect 43069 293115 43135 293118
rect 43253 292770 43319 292773
rect 41492 292768 43319 292770
rect 41492 292712 43258 292768
rect 43314 292712 43319 292768
rect 41492 292710 43319 292712
rect 43253 292707 43319 292710
rect 32765 292362 32831 292365
rect 32765 292360 32844 292362
rect 32765 292304 32770 292360
rect 32826 292304 32844 292360
rect 32765 292302 32844 292304
rect 32765 292299 32831 292302
rect 41781 291954 41847 291957
rect 41492 291952 41847 291954
rect 41492 291896 41786 291952
rect 41842 291896 41847 291952
rect 41492 291894 41847 291896
rect 41781 291891 41847 291894
rect 675753 291682 675819 291685
rect 675886 291682 675892 291684
rect 675753 291680 675892 291682
rect 675753 291624 675758 291680
rect 675814 291624 675892 291680
rect 675753 291622 675892 291624
rect 675753 291619 675819 291622
rect 675886 291620 675892 291622
rect 675956 291620 675962 291684
rect 41781 291546 41847 291549
rect 41492 291544 41847 291546
rect 41492 291488 41786 291544
rect 41842 291488 41847 291544
rect 41492 291486 41847 291488
rect 41781 291483 41847 291486
rect 46381 291138 46447 291141
rect 41492 291136 46447 291138
rect 41492 291080 46386 291136
rect 46442 291080 46447 291136
rect 41492 291078 46447 291080
rect 46381 291075 46447 291078
rect 46105 290730 46171 290733
rect 41492 290728 46171 290730
rect 41492 290672 46110 290728
rect 46166 290672 46171 290728
rect 41492 290670 46171 290672
rect 46105 290667 46171 290670
rect 45369 289914 45435 289917
rect 41492 289912 45435 289914
rect 41492 289856 45374 289912
rect 45430 289856 45435 289912
rect 41492 289854 45435 289856
rect 45369 289851 45435 289854
rect 41638 289172 41644 289236
rect 41708 289234 41714 289236
rect 42374 289234 42380 289236
rect 41708 289174 42380 289234
rect 41708 289172 41714 289174
rect 42374 289172 42380 289174
rect 42444 289172 42450 289236
rect 33041 285970 33107 285973
rect 42374 285970 42380 285972
rect 33041 285968 42380 285970
rect 33041 285912 33046 285968
rect 33102 285912 42380 285968
rect 33041 285910 42380 285912
rect 33041 285907 33107 285910
rect 42374 285908 42380 285910
rect 42444 285908 42450 285972
rect 32949 285834 33015 285837
rect 42190 285834 42196 285836
rect 32949 285832 42196 285834
rect 32949 285776 32954 285832
rect 33010 285776 42196 285832
rect 32949 285774 42196 285776
rect 32949 285771 33015 285774
rect 42190 285772 42196 285774
rect 42260 285772 42266 285836
rect 32581 285698 32647 285701
rect 42558 285698 42564 285700
rect 32581 285696 42564 285698
rect 32581 285640 32586 285696
rect 32642 285640 42564 285696
rect 32581 285638 42564 285640
rect 32581 285635 32647 285638
rect 42558 285636 42564 285638
rect 42628 285636 42634 285700
rect 655329 285290 655395 285293
rect 650164 285288 655395 285290
rect 650164 285232 655334 285288
rect 655390 285232 655395 285288
rect 650164 285230 655395 285232
rect 655329 285227 655395 285230
rect 59445 285154 59511 285157
rect 59445 285152 64492 285154
rect 59445 285096 59450 285152
rect 59506 285096 64492 285152
rect 59445 285094 64492 285096
rect 59445 285091 59511 285094
rect 673678 279690 673684 279692
rect 670928 279630 673684 279690
rect 44030 278428 44036 278492
rect 44100 278490 44106 278492
rect 670928 278490 670988 279630
rect 673678 279628 673684 279630
rect 673748 279628 673754 279692
rect 674046 279554 674052 279556
rect 44100 278430 670988 278490
rect 671064 279494 674052 279554
rect 44100 278428 44106 278430
rect 62297 278354 62363 278357
rect 671064 278354 671124 279494
rect 674046 279492 674052 279494
rect 674116 279492 674122 279556
rect 674414 279418 674420 279420
rect 62297 278352 671124 278354
rect 62297 278296 62302 278352
rect 62358 278296 671124 278352
rect 62297 278294 671124 278296
rect 671200 279358 674420 279418
rect 62297 278291 62363 278294
rect 62665 278218 62731 278221
rect 671200 278218 671260 279358
rect 674414 279356 674420 279358
rect 674484 279356 674490 279420
rect 674230 279282 674236 279284
rect 62665 278216 671260 278218
rect 62665 278160 62670 278216
rect 62726 278160 671260 278216
rect 62665 278158 671260 278160
rect 671336 279222 674236 279282
rect 62665 278155 62731 278158
rect 62481 278082 62547 278085
rect 671336 278082 671396 279222
rect 674230 279220 674236 279222
rect 674300 279220 674306 279284
rect 673862 279146 673868 279148
rect 62481 278080 671396 278082
rect 62481 278024 62486 278080
rect 62542 278024 671396 278080
rect 62481 278022 671396 278024
rect 671472 279086 673868 279146
rect 62481 278019 62547 278022
rect 62849 277946 62915 277949
rect 671472 277946 671532 279086
rect 673862 279084 673868 279086
rect 673932 279084 673938 279148
rect 673494 279010 673500 279012
rect 62849 277944 671532 277946
rect 62849 277888 62854 277944
rect 62910 277888 671532 277944
rect 62849 277886 671532 277888
rect 671608 278950 673500 279010
rect 62849 277883 62915 277886
rect 63033 277810 63099 277813
rect 671608 277810 671668 278950
rect 673494 278948 673500 278950
rect 673564 278948 673570 279012
rect 63033 277808 671668 277810
rect 63033 277752 63038 277808
rect 63094 277752 671668 277808
rect 63033 277750 671668 277752
rect 63033 277747 63099 277750
rect 388253 275906 388319 275909
rect 586053 275906 586119 275909
rect 388253 275904 586119 275906
rect 388253 275848 388258 275904
rect 388314 275848 586058 275904
rect 586114 275848 586119 275904
rect 388253 275846 586119 275848
rect 388253 275843 388319 275846
rect 586053 275843 586119 275846
rect 391289 275770 391355 275773
rect 593137 275770 593203 275773
rect 391289 275768 593203 275770
rect 391289 275712 391294 275768
rect 391350 275712 593142 275768
rect 593198 275712 593203 275768
rect 391289 275710 593203 275712
rect 391289 275707 391355 275710
rect 593137 275707 593203 275710
rect 393589 275634 393655 275637
rect 600221 275634 600287 275637
rect 393589 275632 600287 275634
rect 393589 275576 393594 275632
rect 393650 275576 600226 275632
rect 600282 275576 600287 275632
rect 393589 275574 600287 275576
rect 393589 275571 393655 275574
rect 600221 275571 600287 275574
rect 396257 275498 396323 275501
rect 607305 275498 607371 275501
rect 396257 275496 607371 275498
rect 396257 275440 396262 275496
rect 396318 275440 607310 275496
rect 607366 275440 607371 275496
rect 396257 275438 607371 275440
rect 396257 275435 396323 275438
rect 607305 275435 607371 275438
rect 398925 275362 398991 275365
rect 614389 275362 614455 275365
rect 398925 275360 614455 275362
rect 398925 275304 398930 275360
rect 398986 275304 614394 275360
rect 614450 275304 614455 275360
rect 398925 275302 614455 275304
rect 398925 275299 398991 275302
rect 614389 275299 614455 275302
rect 401685 275226 401751 275229
rect 621473 275226 621539 275229
rect 401685 275224 621539 275226
rect 401685 275168 401690 275224
rect 401746 275168 621478 275224
rect 621534 275168 621539 275224
rect 401685 275166 621539 275168
rect 401685 275163 401751 275166
rect 621473 275163 621539 275166
rect 404261 275090 404327 275093
rect 628557 275090 628623 275093
rect 404261 275088 628623 275090
rect 404261 275032 404266 275088
rect 404322 275032 628562 275088
rect 628618 275032 628623 275088
rect 404261 275030 628623 275032
rect 404261 275027 404327 275030
rect 628557 275027 628623 275030
rect 402697 274954 402763 274957
rect 623865 274954 623931 274957
rect 402697 274952 623931 274954
rect 402697 274896 402702 274952
rect 402758 274896 623870 274952
rect 623926 274896 623931 274952
rect 402697 274894 623931 274896
rect 402697 274891 402763 274894
rect 623865 274891 623931 274894
rect 405457 274818 405523 274821
rect 630949 274818 631015 274821
rect 405457 274816 631015 274818
rect 405457 274760 405462 274816
rect 405518 274760 630954 274816
rect 631010 274760 631015 274816
rect 405457 274758 631015 274760
rect 405457 274755 405523 274758
rect 630949 274755 631015 274758
rect 406929 274682 406995 274685
rect 635641 274682 635707 274685
rect 406929 274680 635707 274682
rect 406929 274624 406934 274680
rect 406990 274624 635646 274680
rect 635702 274624 635707 274680
rect 406929 274622 635707 274624
rect 406929 274619 406995 274622
rect 635641 274619 635707 274622
rect 408217 274546 408283 274549
rect 638033 274546 638099 274549
rect 408217 274544 638099 274546
rect 408217 274488 408222 274544
rect 408278 274488 638038 274544
rect 638094 274488 638099 274544
rect 408217 274486 638099 274488
rect 408217 274483 408283 274486
rect 638033 274483 638099 274486
rect 111977 273186 112043 273189
rect 209221 273186 209287 273189
rect 111977 273184 209287 273186
rect 111977 273128 111982 273184
rect 112038 273128 209226 273184
rect 209282 273128 209287 273184
rect 111977 273126 209287 273128
rect 111977 273123 112043 273126
rect 209221 273123 209287 273126
rect 368657 273186 368723 273189
rect 533981 273186 534047 273189
rect 368657 273184 534047 273186
rect 368657 273128 368662 273184
rect 368718 273128 533986 273184
rect 534042 273128 534047 273184
rect 368657 273126 534047 273128
rect 368657 273123 368723 273126
rect 533981 273123 534047 273126
rect 107193 273050 107259 273053
rect 203517 273050 203583 273053
rect 107193 273048 203583 273050
rect 107193 272992 107198 273048
rect 107254 272992 203522 273048
rect 203578 272992 203583 273048
rect 107193 272990 203583 272992
rect 107193 272987 107259 272990
rect 203517 272987 203583 272990
rect 371233 273050 371299 273053
rect 539869 273050 539935 273053
rect 371233 273048 539935 273050
rect 371233 272992 371238 273048
rect 371294 272992 539874 273048
rect 539930 272992 539935 273048
rect 371233 272990 539935 272992
rect 371233 272987 371299 272990
rect 539869 272987 539935 272990
rect 105997 272914 106063 272917
rect 207473 272914 207539 272917
rect 105997 272912 207539 272914
rect 105997 272856 106002 272912
rect 106058 272856 207478 272912
rect 207534 272856 207539 272912
rect 105997 272854 207539 272856
rect 105997 272851 106063 272854
rect 207473 272851 207539 272854
rect 371325 272914 371391 272917
rect 541065 272914 541131 272917
rect 371325 272912 541131 272914
rect 371325 272856 371330 272912
rect 371386 272856 541070 272912
rect 541126 272856 541131 272912
rect 371325 272854 541131 272856
rect 371325 272851 371391 272854
rect 541065 272851 541131 272854
rect 97717 272778 97783 272781
rect 201309 272778 201375 272781
rect 97717 272776 201375 272778
rect 97717 272720 97722 272776
rect 97778 272720 201314 272776
rect 201370 272720 201375 272776
rect 97717 272718 201375 272720
rect 97717 272715 97783 272718
rect 201309 272715 201375 272718
rect 373993 272778 374059 272781
rect 548149 272778 548215 272781
rect 373993 272776 548215 272778
rect 373993 272720 373998 272776
rect 374054 272720 548154 272776
rect 548210 272720 548215 272776
rect 373993 272718 548215 272720
rect 373993 272715 374059 272718
rect 548149 272715 548215 272718
rect 100109 272642 100175 272645
rect 205725 272642 205791 272645
rect 100109 272640 205791 272642
rect 100109 272584 100114 272640
rect 100170 272584 205730 272640
rect 205786 272584 205791 272640
rect 100109 272582 205791 272584
rect 100109 272579 100175 272582
rect 205725 272579 205791 272582
rect 379329 272642 379395 272645
rect 562409 272642 562475 272645
rect 379329 272640 562475 272642
rect 379329 272584 379334 272640
rect 379390 272584 562414 272640
rect 562470 272584 562475 272640
rect 379329 272582 562475 272584
rect 379329 272579 379395 272582
rect 562409 272579 562475 272582
rect 98913 272506 98979 272509
rect 204805 272506 204871 272509
rect 98913 272504 204871 272506
rect 98913 272448 98918 272504
rect 98974 272448 204810 272504
rect 204866 272448 204871 272504
rect 98913 272446 204871 272448
rect 98913 272443 98979 272446
rect 204805 272443 204871 272446
rect 392761 272506 392827 272509
rect 597829 272506 597895 272509
rect 392761 272504 597895 272506
rect 392761 272448 392766 272504
rect 392822 272448 597834 272504
rect 597890 272448 597895 272504
rect 392761 272446 597895 272448
rect 392761 272443 392827 272446
rect 597829 272443 597895 272446
rect 41965 272372 42031 272373
rect 41965 272368 42012 272372
rect 42076 272370 42082 272372
rect 91829 272370 91895 272373
rect 202137 272370 202203 272373
rect 41965 272312 41970 272368
rect 41965 272308 42012 272312
rect 42076 272310 42122 272370
rect 91829 272368 202203 272370
rect 91829 272312 91834 272368
rect 91890 272312 202142 272368
rect 202198 272312 202203 272368
rect 91829 272310 202203 272312
rect 42076 272308 42082 272310
rect 41965 272307 42031 272308
rect 91829 272307 91895 272310
rect 202137 272307 202203 272310
rect 398097 272370 398163 272373
rect 611997 272370 612063 272373
rect 398097 272368 612063 272370
rect 398097 272312 398102 272368
rect 398158 272312 612002 272368
rect 612058 272312 612063 272368
rect 398097 272310 612063 272312
rect 398097 272307 398163 272310
rect 611997 272307 612063 272310
rect 85941 272234 86007 272237
rect 199929 272234 199995 272237
rect 85941 272232 199995 272234
rect 85941 272176 85946 272232
rect 86002 272176 199934 272232
rect 199990 272176 199995 272232
rect 85941 272174 199995 272176
rect 85941 272171 86007 272174
rect 199929 272171 199995 272174
rect 403433 272234 403499 272237
rect 626165 272234 626231 272237
rect 403433 272232 626231 272234
rect 403433 272176 403438 272232
rect 403494 272176 626170 272232
rect 626226 272176 626231 272232
rect 403433 272174 626231 272176
rect 403433 272171 403499 272174
rect 626165 272171 626231 272174
rect 83549 272098 83615 272101
rect 199101 272098 199167 272101
rect 83549 272096 199167 272098
rect 83549 272040 83554 272096
rect 83610 272040 199106 272096
rect 199162 272040 199167 272096
rect 83549 272038 199167 272040
rect 83549 272035 83615 272038
rect 199101 272035 199167 272038
rect 408769 272098 408835 272101
rect 640425 272098 640491 272101
rect 408769 272096 640491 272098
rect 408769 272040 408774 272096
rect 408830 272040 640430 272096
rect 640486 272040 640491 272096
rect 408769 272038 640491 272040
rect 408769 272035 408835 272038
rect 640425 272035 640491 272038
rect 76465 271962 76531 271965
rect 196341 271962 196407 271965
rect 76465 271960 196407 271962
rect 76465 271904 76470 271960
rect 76526 271904 196346 271960
rect 196402 271904 196407 271960
rect 76465 271902 196407 271904
rect 76465 271899 76531 271902
rect 196341 271899 196407 271902
rect 410517 271962 410583 271965
rect 645117 271962 645183 271965
rect 410517 271960 645183 271962
rect 410517 271904 410522 271960
rect 410578 271904 645122 271960
rect 645178 271904 645183 271960
rect 410517 271902 645183 271904
rect 410517 271899 410583 271902
rect 645117 271899 645183 271902
rect 70577 271826 70643 271829
rect 194133 271826 194199 271829
rect 70577 271824 194199 271826
rect 70577 271768 70582 271824
rect 70638 271768 194138 271824
rect 194194 271768 194199 271824
rect 70577 271766 194199 271768
rect 70577 271763 70643 271766
rect 194133 271763 194199 271766
rect 194501 271826 194567 271829
rect 208485 271826 208551 271829
rect 194501 271824 208551 271826
rect 194501 271768 194506 271824
rect 194562 271768 208490 271824
rect 208546 271768 208551 271824
rect 194501 271766 208551 271768
rect 194501 271763 194567 271766
rect 208485 271763 208551 271766
rect 410885 271826 410951 271829
rect 646313 271826 646379 271829
rect 410885 271824 646379 271826
rect 410885 271768 410890 271824
rect 410946 271768 646318 271824
rect 646374 271768 646379 271824
rect 410885 271766 646379 271768
rect 410885 271763 410951 271766
rect 646313 271763 646379 271766
rect 115473 271690 115539 271693
rect 210601 271690 210667 271693
rect 115473 271688 210667 271690
rect 115473 271632 115478 271688
rect 115534 271632 210606 271688
rect 210662 271632 210667 271688
rect 115473 271630 210667 271632
rect 115473 271627 115539 271630
rect 210601 271627 210667 271630
rect 365989 271690 366055 271693
rect 526897 271690 526963 271693
rect 365989 271688 526963 271690
rect 365989 271632 365994 271688
rect 366050 271632 526902 271688
rect 526958 271632 526963 271688
rect 365989 271630 526963 271632
rect 365989 271627 366055 271630
rect 526897 271627 526963 271630
rect 122557 271554 122623 271557
rect 213269 271554 213335 271557
rect 122557 271552 213335 271554
rect 122557 271496 122562 271552
rect 122618 271496 213274 271552
rect 213330 271496 213335 271552
rect 122557 271494 213335 271496
rect 122557 271491 122623 271494
rect 213269 271491 213335 271494
rect 365529 271554 365595 271557
rect 525701 271554 525767 271557
rect 365529 271552 525767 271554
rect 365529 271496 365534 271552
rect 365590 271496 525706 271552
rect 525762 271496 525767 271552
rect 365529 271494 525767 271496
rect 365529 271491 365595 271494
rect 525701 271491 525767 271494
rect 363321 271418 363387 271421
rect 519813 271418 519879 271421
rect 363321 271416 519879 271418
rect 363321 271360 363326 271416
rect 363382 271360 519818 271416
rect 519874 271360 519879 271416
rect 363321 271358 519879 271360
rect 363321 271355 363387 271358
rect 519813 271355 519879 271358
rect 42149 270466 42215 270469
rect 42558 270466 42564 270468
rect 42149 270464 42564 270466
rect 42149 270408 42154 270464
rect 42210 270408 42564 270464
rect 42149 270406 42564 270408
rect 42149 270403 42215 270406
rect 42558 270404 42564 270406
rect 42628 270404 42634 270468
rect 121361 270466 121427 270469
rect 213729 270466 213795 270469
rect 121361 270464 213795 270466
rect 121361 270408 121366 270464
rect 121422 270408 213734 270464
rect 213790 270408 213795 270464
rect 121361 270406 213795 270408
rect 121361 270403 121427 270406
rect 213729 270403 213795 270406
rect 366909 270466 366975 270469
rect 529289 270466 529355 270469
rect 366909 270464 529355 270466
rect 366909 270408 366914 270464
rect 366970 270408 529294 270464
rect 529350 270408 529355 270464
rect 366909 270406 529355 270408
rect 366909 270403 366975 270406
rect 529289 270403 529355 270406
rect 108389 270330 108455 270333
rect 207933 270330 207999 270333
rect 108389 270328 207999 270330
rect 108389 270272 108394 270328
rect 108450 270272 207938 270328
rect 207994 270272 207999 270328
rect 108389 270270 207999 270272
rect 108389 270267 108455 270270
rect 207933 270267 207999 270270
rect 369577 270330 369643 270333
rect 536373 270330 536439 270333
rect 369577 270328 536439 270330
rect 369577 270272 369582 270328
rect 369638 270272 536378 270328
rect 536434 270272 536439 270328
rect 369577 270270 536439 270272
rect 369577 270267 369643 270270
rect 536373 270267 536439 270270
rect 103697 270194 103763 270197
rect 207013 270194 207079 270197
rect 103697 270192 207079 270194
rect 103697 270136 103702 270192
rect 103758 270136 207018 270192
rect 207074 270136 207079 270192
rect 103697 270134 207079 270136
rect 103697 270131 103763 270134
rect 207013 270131 207079 270134
rect 372245 270194 372311 270197
rect 543457 270194 543523 270197
rect 372245 270192 543523 270194
rect 372245 270136 372250 270192
rect 372306 270136 543462 270192
rect 543518 270136 543523 270192
rect 372245 270134 543523 270136
rect 372245 270131 372311 270134
rect 543457 270131 543523 270134
rect 42149 270058 42215 270061
rect 42374 270058 42380 270060
rect 42149 270056 42380 270058
rect 42149 270000 42154 270056
rect 42210 270000 42380 270056
rect 42149 269998 42380 270000
rect 42149 269995 42215 269998
rect 42374 269996 42380 269998
rect 42444 269996 42450 270060
rect 101305 270058 101371 270061
rect 205265 270058 205331 270061
rect 101305 270056 205331 270058
rect 101305 270000 101310 270056
rect 101366 270000 205270 270056
rect 205326 270000 205331 270056
rect 101305 269998 205331 270000
rect 101305 269995 101371 269998
rect 205265 269995 205331 269998
rect 378041 270058 378107 270061
rect 558821 270058 558887 270061
rect 378041 270056 558887 270058
rect 378041 270000 378046 270056
rect 378102 270000 558826 270056
rect 558882 270000 558887 270056
rect 378041 269998 558887 270000
rect 378041 269995 378107 269998
rect 558821 269995 558887 269998
rect 96613 269922 96679 269925
rect 204345 269922 204411 269925
rect 96613 269920 204411 269922
rect 96613 269864 96618 269920
rect 96674 269864 204350 269920
rect 204406 269864 204411 269920
rect 96613 269862 204411 269864
rect 96613 269859 96679 269862
rect 204345 269859 204411 269862
rect 383377 269922 383443 269925
rect 572989 269922 573055 269925
rect 383377 269920 573055 269922
rect 383377 269864 383382 269920
rect 383438 269864 572994 269920
rect 573050 269864 573055 269920
rect 383377 269862 573055 269864
rect 383377 269859 383443 269862
rect 572989 269859 573055 269862
rect 90633 269786 90699 269789
rect 201677 269786 201743 269789
rect 90633 269784 201743 269786
rect 90633 269728 90638 269784
rect 90694 269728 201682 269784
rect 201738 269728 201743 269784
rect 90633 269726 201743 269728
rect 90633 269723 90699 269726
rect 201677 269723 201743 269726
rect 391381 269786 391447 269789
rect 594333 269786 594399 269789
rect 391381 269784 594399 269786
rect 391381 269728 391386 269784
rect 391442 269728 594338 269784
rect 594394 269728 594399 269784
rect 391381 269726 594399 269728
rect 391381 269723 391447 269726
rect 594333 269723 594399 269726
rect 87137 269650 87203 269653
rect 200389 269650 200455 269653
rect 87137 269648 200455 269650
rect 87137 269592 87142 269648
rect 87198 269592 200394 269648
rect 200450 269592 200455 269648
rect 87137 269590 200455 269592
rect 87137 269587 87203 269590
rect 200389 269587 200455 269590
rect 402053 269650 402119 269653
rect 622669 269650 622735 269653
rect 402053 269648 622735 269650
rect 402053 269592 402058 269648
rect 402114 269592 622674 269648
rect 622730 269592 622735 269648
rect 402053 269590 622735 269592
rect 402053 269587 402119 269590
rect 622669 269587 622735 269590
rect 84745 269514 84811 269517
rect 199009 269514 199075 269517
rect 84745 269512 199075 269514
rect 84745 269456 84750 269512
rect 84806 269456 199014 269512
rect 199070 269456 199075 269512
rect 84745 269454 199075 269456
rect 84745 269451 84811 269454
rect 199009 269451 199075 269454
rect 404721 269514 404787 269517
rect 629753 269514 629819 269517
rect 404721 269512 629819 269514
rect 404721 269456 404726 269512
rect 404782 269456 629758 269512
rect 629814 269456 629819 269512
rect 404721 269454 629819 269456
rect 404721 269451 404787 269454
rect 629753 269451 629819 269454
rect 42149 269380 42215 269381
rect 42149 269378 42196 269380
rect 42104 269376 42196 269378
rect 42104 269320 42154 269376
rect 42104 269318 42196 269320
rect 42149 269316 42196 269318
rect 42260 269316 42266 269380
rect 78857 269378 78923 269381
rect 197721 269378 197787 269381
rect 78857 269376 197787 269378
rect 78857 269320 78862 269376
rect 78918 269320 197726 269376
rect 197782 269320 197787 269376
rect 78857 269318 197787 269320
rect 42149 269315 42215 269316
rect 78857 269315 78923 269318
rect 197721 269315 197787 269318
rect 407389 269378 407455 269381
rect 636837 269378 636903 269381
rect 407389 269376 636903 269378
rect 407389 269320 407394 269376
rect 407450 269320 636842 269376
rect 636898 269320 636903 269376
rect 407389 269318 636903 269320
rect 407389 269315 407455 269318
rect 636837 269315 636903 269318
rect 77661 269242 77727 269245
rect 196801 269242 196867 269245
rect 77661 269240 196867 269242
rect 77661 269184 77666 269240
rect 77722 269184 196806 269240
rect 196862 269184 196867 269240
rect 77661 269182 196867 269184
rect 77661 269179 77727 269182
rect 196801 269179 196867 269182
rect 409597 269242 409663 269245
rect 642725 269242 642791 269245
rect 409597 269240 642791 269242
rect 409597 269184 409602 269240
rect 409658 269184 642730 269240
rect 642786 269184 642791 269240
rect 409597 269182 642791 269184
rect 409597 269179 409663 269182
rect 642725 269179 642791 269182
rect 69381 269106 69447 269109
rect 193673 269106 193739 269109
rect 69381 269104 193739 269106
rect 69381 269048 69386 269104
rect 69442 269048 193678 269104
rect 193734 269048 193739 269104
rect 69381 269046 193739 269048
rect 69381 269043 69447 269046
rect 193673 269043 193739 269046
rect 410057 269106 410123 269109
rect 643921 269106 643987 269109
rect 410057 269104 643987 269106
rect 410057 269048 410062 269104
rect 410118 269048 643926 269104
rect 643982 269048 643987 269104
rect 410057 269046 643987 269048
rect 410057 269043 410123 269046
rect 643921 269043 643987 269046
rect 128537 268970 128603 268973
rect 216397 268970 216463 268973
rect 128537 268968 216463 268970
rect 128537 268912 128542 268968
rect 128598 268912 216402 268968
rect 216458 268912 216463 268968
rect 128537 268910 216463 268912
rect 128537 268907 128603 268910
rect 216397 268907 216463 268910
rect 364241 268970 364307 268973
rect 522205 268970 522271 268973
rect 364241 268968 522271 268970
rect 364241 268912 364246 268968
rect 364302 268912 522210 268968
rect 522266 268912 522271 268968
rect 364241 268910 522271 268912
rect 364241 268907 364307 268910
rect 522205 268907 522271 268910
rect 127341 268834 127407 268837
rect 215477 268834 215543 268837
rect 127341 268832 215543 268834
rect 127341 268776 127346 268832
rect 127402 268776 215482 268832
rect 215538 268776 215543 268832
rect 127341 268774 215543 268776
rect 127341 268771 127407 268774
rect 215477 268771 215543 268774
rect 362033 268834 362099 268837
rect 516225 268834 516291 268837
rect 362033 268832 516291 268834
rect 362033 268776 362038 268832
rect 362094 268776 516230 268832
rect 516286 268776 516291 268832
rect 362033 268774 516291 268776
rect 362033 268771 362099 268774
rect 516225 268771 516291 268774
rect 142705 268698 142771 268701
rect 221733 268698 221799 268701
rect 142705 268696 221799 268698
rect 142705 268640 142710 268696
rect 142766 268640 221738 268696
rect 221794 268640 221799 268696
rect 142705 268638 221799 268640
rect 142705 268635 142771 268638
rect 221733 268635 221799 268638
rect 358905 268698 358971 268701
rect 507945 268698 508011 268701
rect 358905 268696 508011 268698
rect 358905 268640 358910 268696
rect 358966 268640 507950 268696
rect 508006 268640 508011 268696
rect 358905 268638 508011 268640
rect 358905 268635 358971 268638
rect 507945 268635 508011 268638
rect 153285 268562 153351 268565
rect 225781 268562 225847 268565
rect 153285 268560 225847 268562
rect 153285 268504 153290 268560
rect 153346 268504 225786 268560
rect 225842 268504 225847 268560
rect 153285 268502 225847 268504
rect 153285 268499 153351 268502
rect 225781 268499 225847 268502
rect 359365 268562 359431 268565
rect 509141 268562 509207 268565
rect 359365 268560 509207 268562
rect 359365 268504 359370 268560
rect 359426 268504 509146 268560
rect 509202 268504 509207 268560
rect 359365 268502 509207 268504
rect 359365 268499 359431 268502
rect 509141 268499 509207 268502
rect 676121 268562 676187 268565
rect 676262 268562 676322 268668
rect 676121 268560 676322 268562
rect 676121 268504 676126 268560
rect 676182 268504 676322 268560
rect 676121 268502 676322 268504
rect 676121 268499 676187 268502
rect 184933 268426 184999 268429
rect 203057 268426 203123 268429
rect 184933 268424 203123 268426
rect 184933 268368 184938 268424
rect 184994 268368 203062 268424
rect 203118 268368 203123 268424
rect 184933 268366 203123 268368
rect 184933 268363 184999 268366
rect 203057 268363 203123 268366
rect 356605 268426 356671 268429
rect 502057 268426 502123 268429
rect 356605 268424 502123 268426
rect 356605 268368 356610 268424
rect 356666 268368 502062 268424
rect 502118 268368 502123 268424
rect 356605 268366 502123 268368
rect 356605 268363 356671 268366
rect 502057 268363 502123 268366
rect 353937 268290 354003 268293
rect 494973 268290 495039 268293
rect 353937 268288 495039 268290
rect 353937 268232 353942 268288
rect 353998 268232 494978 268288
rect 495034 268232 495039 268288
rect 353937 268230 495039 268232
rect 353937 268227 354003 268230
rect 494973 268227 495039 268230
rect 676262 268157 676322 268260
rect 203517 268154 203583 268157
rect 208393 268154 208459 268157
rect 203517 268152 208459 268154
rect 203517 268096 203522 268152
rect 203578 268096 208398 268152
rect 208454 268096 208459 268152
rect 203517 268094 208459 268096
rect 203517 268091 203583 268094
rect 208393 268091 208459 268094
rect 676213 268152 676322 268157
rect 676213 268096 676218 268152
rect 676274 268096 676322 268152
rect 676213 268094 676322 268096
rect 676213 268091 676279 268094
rect 676029 267882 676095 267885
rect 676029 267880 676292 267882
rect 676029 267824 676034 267880
rect 676090 267824 676292 267880
rect 676029 267822 676292 267824
rect 676029 267819 676095 267822
rect 387793 267746 387859 267749
rect 584857 267746 584923 267749
rect 387793 267744 584923 267746
rect 387793 267688 387798 267744
rect 387854 267688 584862 267744
rect 584918 267688 584923 267744
rect 387793 267686 584923 267688
rect 387793 267683 387859 267686
rect 584857 267683 584923 267686
rect 386965 267610 387031 267613
rect 582465 267610 582531 267613
rect 386965 267608 582531 267610
rect 386965 267552 386970 267608
rect 387026 267552 582470 267608
rect 582526 267552 582531 267608
rect 386965 267550 582531 267552
rect 386965 267547 387031 267550
rect 582465 267547 582531 267550
rect 389633 267474 389699 267477
rect 589549 267474 589615 267477
rect 389633 267472 589615 267474
rect 389633 267416 389638 267472
rect 389694 267416 589554 267472
rect 589610 267416 589615 267472
rect 389633 267414 589615 267416
rect 389633 267411 389699 267414
rect 589549 267411 589615 267414
rect 675937 267474 676003 267477
rect 675937 267472 676292 267474
rect 675937 267416 675942 267472
rect 675998 267416 676292 267472
rect 675937 267414 676292 267416
rect 675937 267411 676003 267414
rect 390461 267338 390527 267341
rect 591941 267338 592007 267341
rect 390461 267336 592007 267338
rect 390461 267280 390466 267336
rect 390522 267280 591946 267336
rect 592002 267280 592007 267336
rect 390461 267278 592007 267280
rect 390461 267275 390527 267278
rect 591941 267275 592007 267278
rect 391841 267202 391907 267205
rect 595437 267202 595503 267205
rect 391841 267200 595503 267202
rect 391841 267144 391846 267200
rect 391902 267144 595442 267200
rect 595498 267144 595503 267200
rect 391841 267142 595503 267144
rect 391841 267139 391907 267142
rect 595437 267139 595503 267142
rect 393129 267066 393195 267069
rect 599025 267066 599091 267069
rect 393129 267064 599091 267066
rect 393129 267008 393134 267064
rect 393190 267008 599030 267064
rect 599086 267008 599091 267064
rect 393129 267006 599091 267008
rect 393129 267003 393195 267006
rect 599025 267003 599091 267006
rect 675753 267066 675819 267069
rect 675753 267064 676292 267066
rect 675753 267008 675758 267064
rect 675814 267008 676292 267064
rect 675753 267006 676292 267008
rect 675753 267003 675819 267006
rect 394509 266930 394575 266933
rect 602521 266930 602587 266933
rect 394509 266928 602587 266930
rect 394509 266872 394514 266928
rect 394570 266872 602526 266928
rect 602582 266872 602587 266928
rect 394509 266870 602587 266872
rect 394509 266867 394575 266870
rect 602521 266867 602587 266870
rect 395797 266794 395863 266797
rect 606109 266794 606175 266797
rect 395797 266792 606175 266794
rect 395797 266736 395802 266792
rect 395858 266736 606114 266792
rect 606170 266736 606175 266792
rect 395797 266734 606175 266736
rect 395797 266731 395863 266734
rect 606109 266731 606175 266734
rect 397177 266658 397243 266661
rect 609697 266658 609763 266661
rect 397177 266656 609763 266658
rect 397177 266600 397182 266656
rect 397238 266600 609702 266656
rect 609758 266600 609763 266656
rect 397177 266598 609763 266600
rect 397177 266595 397243 266598
rect 609697 266595 609763 266598
rect 676029 266658 676095 266661
rect 676029 266656 676292 266658
rect 676029 266600 676034 266656
rect 676090 266600 676292 266656
rect 676029 266598 676292 266600
rect 676029 266595 676095 266598
rect 398465 266522 398531 266525
rect 613193 266522 613259 266525
rect 398465 266520 613259 266522
rect 398465 266464 398470 266520
rect 398526 266464 613198 266520
rect 613254 266464 613259 266520
rect 398465 266462 613259 266464
rect 398465 266459 398531 266462
rect 613193 266459 613259 266462
rect 399845 266386 399911 266389
rect 616781 266386 616847 266389
rect 399845 266384 616847 266386
rect 399845 266328 399850 266384
rect 399906 266328 616786 266384
rect 616842 266328 616847 266384
rect 399845 266326 616847 266328
rect 399845 266323 399911 266326
rect 616781 266323 616847 266326
rect 386505 266250 386571 266253
rect 581269 266250 581335 266253
rect 386505 266248 581335 266250
rect 386505 266192 386510 266248
rect 386566 266192 581274 266248
rect 581330 266192 581335 266248
rect 386505 266190 581335 266192
rect 386505 266187 386571 266190
rect 581269 266187 581335 266190
rect 676029 266250 676095 266253
rect 676029 266248 676292 266250
rect 676029 266192 676034 266248
rect 676090 266192 676292 266248
rect 676029 266190 676292 266192
rect 676029 266187 676095 266190
rect 385125 266114 385191 266117
rect 577773 266114 577839 266117
rect 385125 266112 577839 266114
rect 385125 266056 385130 266112
rect 385186 266056 577778 266112
rect 577834 266056 577839 266112
rect 385125 266054 577839 266056
rect 385125 266051 385191 266054
rect 577773 266051 577839 266054
rect 676213 266114 676279 266117
rect 676213 266112 676322 266114
rect 676213 266056 676218 266112
rect 676274 266056 676322 266112
rect 676213 266051 676322 266056
rect 405641 265978 405707 265981
rect 466269 265978 466335 265981
rect 405641 265976 466335 265978
rect 405641 265920 405646 265976
rect 405702 265920 466274 265976
rect 466330 265920 466335 265976
rect 405641 265918 466335 265920
rect 405641 265915 405707 265918
rect 466269 265915 466335 265918
rect 408309 265842 408375 265845
rect 459461 265842 459527 265845
rect 408309 265840 459527 265842
rect 408309 265784 408314 265840
rect 408370 265784 459466 265840
rect 459522 265784 459527 265840
rect 676262 265812 676322 266051
rect 408309 265782 459527 265784
rect 408309 265779 408375 265782
rect 459461 265779 459527 265782
rect 675661 265434 675727 265437
rect 675661 265432 676292 265434
rect 675661 265376 675666 265432
rect 675722 265376 676292 265432
rect 675661 265374 676292 265376
rect 675661 265371 675727 265374
rect 676262 264893 676322 264996
rect 676213 264888 676322 264893
rect 676213 264832 676218 264888
rect 676274 264832 676322 264888
rect 676213 264830 676322 264832
rect 676213 264827 676279 264830
rect 674230 264556 674236 264620
rect 674300 264618 674306 264620
rect 674300 264558 676292 264618
rect 674300 264556 674306 264558
rect 676029 264210 676095 264213
rect 676029 264208 676292 264210
rect 676029 264152 676034 264208
rect 676090 264152 676292 264208
rect 676029 264150 676292 264152
rect 676029 264147 676095 264150
rect 676121 263666 676187 263669
rect 676262 263666 676322 263772
rect 676121 263664 676322 263666
rect 676121 263608 676126 263664
rect 676182 263608 676322 263664
rect 676121 263606 676322 263608
rect 676121 263603 676187 263606
rect 675845 263394 675911 263397
rect 675845 263392 676292 263394
rect 675845 263336 675850 263392
rect 675906 263336 676292 263392
rect 675845 263334 676292 263336
rect 675845 263331 675911 263334
rect 676029 262986 676095 262989
rect 676029 262984 676292 262986
rect 676029 262928 676034 262984
rect 676090 262928 676292 262984
rect 676029 262926 676292 262928
rect 676029 262923 676095 262926
rect 658181 262442 658247 262445
rect 674230 262442 674236 262444
rect 658181 262440 674236 262442
rect 658181 262384 658186 262440
rect 658242 262384 674236 262440
rect 658181 262382 674236 262384
rect 658181 262379 658247 262382
rect 674230 262380 674236 262382
rect 674300 262442 674306 262444
rect 675886 262442 675892 262444
rect 674300 262382 675892 262442
rect 674300 262380 674306 262382
rect 675886 262380 675892 262382
rect 675956 262380 675962 262444
rect 676121 262442 676187 262445
rect 676262 262442 676322 262548
rect 676121 262440 676322 262442
rect 676121 262384 676126 262440
rect 676182 262384 676322 262440
rect 676121 262382 676322 262384
rect 676121 262379 676187 262382
rect 416773 262306 416839 262309
rect 412436 262304 416839 262306
rect 412436 262248 416778 262304
rect 416834 262248 416839 262304
rect 412436 262246 416839 262248
rect 416773 262243 416839 262246
rect 676029 262170 676095 262173
rect 676029 262168 676292 262170
rect 676029 262112 676034 262168
rect 676090 262112 676292 262168
rect 676029 262110 676292 262112
rect 676029 262107 676095 262110
rect 676029 261762 676095 261765
rect 676029 261760 676292 261762
rect 676029 261704 676034 261760
rect 676090 261704 676292 261760
rect 676029 261702 676292 261704
rect 676029 261699 676095 261702
rect 676121 261218 676187 261221
rect 676262 261218 676322 261324
rect 676121 261216 676322 261218
rect 676121 261160 676126 261216
rect 676182 261160 676322 261216
rect 676121 261158 676322 261160
rect 676121 261155 676187 261158
rect 675937 260946 676003 260949
rect 675937 260944 676292 260946
rect 675937 260888 675942 260944
rect 675998 260888 676292 260944
rect 675937 260886 676292 260888
rect 675937 260883 676003 260886
rect 675569 260538 675635 260541
rect 675569 260536 676292 260538
rect 675569 260480 675574 260536
rect 675630 260480 676292 260536
rect 675569 260478 676292 260480
rect 675569 260475 675635 260478
rect 675569 260130 675635 260133
rect 675569 260128 676292 260130
rect 675569 260072 675574 260128
rect 675630 260072 676292 260128
rect 675569 260070 676292 260072
rect 675569 260067 675635 260070
rect 676121 259586 676187 259589
rect 676262 259586 676322 259692
rect 676121 259584 676322 259586
rect 676121 259528 676126 259584
rect 676182 259528 676322 259584
rect 676121 259526 676322 259528
rect 676121 259523 676187 259526
rect 676029 259314 676095 259317
rect 676029 259312 676292 259314
rect 676029 259256 676034 259312
rect 676090 259256 676292 259312
rect 676029 259254 676292 259256
rect 676029 259251 676095 259254
rect 416773 259178 416839 259181
rect 412436 259176 416839 259178
rect 412436 259120 416778 259176
rect 416834 259120 416839 259176
rect 412436 259118 416839 259120
rect 416773 259115 416839 259118
rect 676121 258770 676187 258773
rect 676262 258770 676322 258876
rect 676121 258768 676322 258770
rect 676121 258712 676126 258768
rect 676182 258712 676322 258768
rect 676121 258710 676322 258712
rect 676121 258707 676187 258710
rect 184933 258634 184999 258637
rect 184933 258632 191820 258634
rect 184933 258576 184938 258632
rect 184994 258576 191820 258632
rect 184933 258574 191820 258576
rect 184933 258571 184999 258574
rect 679022 258365 679082 258468
rect 41505 258362 41571 258365
rect 41462 258360 41571 258362
rect 41462 258304 41510 258360
rect 41566 258304 41571 258360
rect 41462 258299 41571 258304
rect 678973 258360 679082 258365
rect 678973 258304 678978 258360
rect 679034 258304 679082 258360
rect 678973 258302 679082 258304
rect 678973 258299 679039 258302
rect 41462 258060 41522 258299
rect 41505 257954 41571 257957
rect 41462 257952 41571 257954
rect 41462 257896 41510 257952
rect 41566 257896 41571 257952
rect 41462 257891 41571 257896
rect 41462 257652 41522 257891
rect 684542 257652 684602 258060
rect 41505 257546 41571 257549
rect 41462 257544 41571 257546
rect 41462 257488 41510 257544
rect 41566 257488 41571 257544
rect 41462 257483 41571 257488
rect 678973 257546 679039 257549
rect 678973 257544 679082 257546
rect 678973 257488 678978 257544
rect 679034 257488 679082 257544
rect 678973 257483 679082 257488
rect 41462 257244 41522 257483
rect 679022 257244 679082 257483
rect 41781 256866 41847 256869
rect 42190 256866 42196 256868
rect 41492 256864 42196 256866
rect 41492 256808 41786 256864
rect 41842 256808 42196 256864
rect 41492 256806 42196 256808
rect 41781 256803 41847 256806
rect 42190 256804 42196 256806
rect 42260 256804 42266 256868
rect 41462 256322 41522 256428
rect 41638 256322 41644 256324
rect 41462 256262 41644 256322
rect 41638 256260 41644 256262
rect 41708 256260 41714 256324
rect 43437 256050 43503 256053
rect 41492 256048 43503 256050
rect 41492 255992 43442 256048
rect 43498 255992 43503 256048
rect 41492 255990 43503 255992
rect 43437 255987 43503 255990
rect 416773 255914 416839 255917
rect 412436 255912 416839 255914
rect 412436 255856 416778 255912
rect 416834 255856 416839 255912
rect 412436 255854 416839 255856
rect 416773 255851 416839 255854
rect 43437 255642 43503 255645
rect 41492 255640 43503 255642
rect 41492 255584 43442 255640
rect 43498 255584 43503 255640
rect 41492 255582 43503 255584
rect 43437 255579 43503 255582
rect 42006 255234 42012 255236
rect 41492 255174 42012 255234
rect 42006 255172 42012 255174
rect 42076 255234 42082 255236
rect 45921 255234 45987 255237
rect 42076 255232 45987 255234
rect 42076 255176 45926 255232
rect 45982 255176 45987 255232
rect 42076 255174 45987 255176
rect 42076 255172 42082 255174
rect 45921 255171 45987 255174
rect 41454 255036 41460 255100
rect 41524 255036 41530 255100
rect 41462 254796 41522 255036
rect 45737 254418 45803 254421
rect 41492 254416 45803 254418
rect 41492 254388 45742 254416
rect 41462 254360 45742 254388
rect 45798 254360 45803 254416
rect 41462 254358 45803 254360
rect 41462 254284 41522 254358
rect 45737 254355 45803 254358
rect 41454 254220 41460 254284
rect 41524 254220 41530 254284
rect 41822 254010 41828 254012
rect 41492 253950 41828 254010
rect 41822 253948 41828 253950
rect 41892 253948 41898 254012
rect 42701 253602 42767 253605
rect 41492 253600 42767 253602
rect 41492 253544 42706 253600
rect 42762 253544 42767 253600
rect 41492 253542 42767 253544
rect 42701 253539 42767 253542
rect 31710 253061 31770 253164
rect 31661 253056 31770 253061
rect 31661 253000 31666 253056
rect 31722 253000 31770 253056
rect 31661 252998 31770 253000
rect 31661 252995 31727 252998
rect 42006 252786 42012 252788
rect 41492 252726 42012 252786
rect 42006 252724 42012 252726
rect 42076 252724 42082 252788
rect 416773 252786 416839 252789
rect 412436 252784 416839 252786
rect 412436 252728 416778 252784
rect 416834 252728 416839 252784
rect 412436 252726 416839 252728
rect 416773 252723 416839 252726
rect 42793 252378 42859 252381
rect 41492 252376 42859 252378
rect 41492 252320 42798 252376
rect 42854 252320 42859 252376
rect 41492 252318 42859 252320
rect 42793 252315 42859 252318
rect 32998 251837 33058 251940
rect 32998 251832 33107 251837
rect 32998 251776 33046 251832
rect 33102 251776 33107 251832
rect 32998 251774 33107 251776
rect 33041 251771 33107 251774
rect 43805 251562 43871 251565
rect 41492 251560 43871 251562
rect 41492 251504 43810 251560
rect 43866 251504 43871 251560
rect 41492 251502 43871 251504
rect 43805 251499 43871 251502
rect 43897 251154 43963 251157
rect 41492 251152 43963 251154
rect 41492 251096 43902 251152
rect 43958 251096 43963 251152
rect 41492 251094 43963 251096
rect 43897 251091 43963 251094
rect 32814 250613 32874 250716
rect 32765 250608 32874 250613
rect 32765 250552 32770 250608
rect 32826 250552 32874 250608
rect 32765 250550 32874 250552
rect 32765 250547 32831 250550
rect 32814 250205 32874 250308
rect 32814 250200 32923 250205
rect 32814 250144 32862 250200
rect 32918 250144 32923 250200
rect 32814 250142 32923 250144
rect 32857 250139 32923 250142
rect 32998 249797 33058 249900
rect 32949 249792 33058 249797
rect 32949 249736 32954 249792
rect 33010 249736 33058 249792
rect 32949 249734 33058 249736
rect 32949 249731 33015 249734
rect 43253 249522 43319 249525
rect 416773 249522 416839 249525
rect 41492 249520 43319 249522
rect 41492 249464 43258 249520
rect 43314 249464 43319 249520
rect 41492 249462 43319 249464
rect 412436 249520 416839 249522
rect 412436 249464 416778 249520
rect 416834 249464 416839 249520
rect 412436 249462 416839 249464
rect 43253 249459 43319 249462
rect 416773 249459 416839 249462
rect 43345 249114 43411 249117
rect 41492 249112 43411 249114
rect 41492 249056 43350 249112
rect 43406 249056 43411 249112
rect 41492 249054 43411 249056
rect 43345 249051 43411 249054
rect 43161 248706 43227 248709
rect 41492 248704 43227 248706
rect 41492 248648 43166 248704
rect 43222 248648 43227 248704
rect 41492 248646 43227 248648
rect 43161 248643 43227 248646
rect 38334 248165 38394 248268
rect 38285 248160 38394 248165
rect 38285 248104 38290 248160
rect 38346 248104 38394 248160
rect 38285 248102 38394 248104
rect 38285 248099 38351 248102
rect 184933 248026 184999 248029
rect 184933 248024 191820 248026
rect 184933 247968 184938 248024
rect 184994 247968 191820 248024
rect 184933 247966 191820 247968
rect 184933 247963 184999 247966
rect 41462 247757 41522 247860
rect 41462 247752 41571 247757
rect 41462 247696 41510 247752
rect 41566 247696 41571 247752
rect 41462 247694 41571 247696
rect 41505 247691 41571 247694
rect 41462 247349 41522 247452
rect 41462 247344 41571 247349
rect 41462 247288 41510 247344
rect 41566 247288 41571 247344
rect 41462 247286 41571 247288
rect 41505 247283 41571 247286
rect 41462 246533 41522 246636
rect 41462 246528 41571 246533
rect 41462 246472 41510 246528
rect 41566 246472 41571 246528
rect 41462 246470 41571 246472
rect 41505 246467 41571 246470
rect 416773 246394 416839 246397
rect 412436 246392 416839 246394
rect 412436 246336 416778 246392
rect 416834 246336 416839 246392
rect 412436 246334 416839 246336
rect 416773 246331 416839 246334
rect 418061 243130 418127 243133
rect 412436 243128 418127 243130
rect 412436 243072 418066 243128
rect 418122 243072 418127 243128
rect 412436 243070 418127 243072
rect 418061 243067 418127 243070
rect 418153 240002 418219 240005
rect 412436 240000 418219 240002
rect 412436 239944 418158 240000
rect 418214 239944 418219 240000
rect 412436 239942 418219 239944
rect 418153 239939 418219 239942
rect 184933 237418 184999 237421
rect 184933 237416 191820 237418
rect 184933 237360 184938 237416
rect 184994 237360 191820 237416
rect 184933 237358 191820 237360
rect 184933 237355 184999 237358
rect 418429 236738 418495 236741
rect 412436 236736 418495 236738
rect 412436 236680 418434 236736
rect 418490 236680 418495 236736
rect 412436 236678 418495 236680
rect 418429 236675 418495 236678
rect 418521 233610 418587 233613
rect 412436 233608 418587 233610
rect 412436 233552 418526 233608
rect 418582 233552 418587 233608
rect 412436 233550 418587 233552
rect 418521 233547 418587 233550
rect 93025 228986 93091 228989
rect 210049 228986 210115 228989
rect 93025 228984 210115 228986
rect 93025 228928 93030 228984
rect 93086 228928 210054 228984
rect 210110 228928 210115 228984
rect 93025 228926 210115 228928
rect 93025 228923 93091 228926
rect 210049 228923 210115 228926
rect 256693 228986 256759 228989
rect 261753 228986 261819 228989
rect 256693 228984 261819 228986
rect 256693 228928 256698 228984
rect 256754 228928 261758 228984
rect 261814 228928 261819 228984
rect 256693 228926 261819 228928
rect 256693 228923 256759 228926
rect 261753 228923 261819 228926
rect 383653 228986 383719 228989
rect 504541 228986 504607 228989
rect 383653 228984 504607 228986
rect 383653 228928 383658 228984
rect 383714 228928 504546 228984
rect 504602 228928 504607 228984
rect 383653 228926 504607 228928
rect 383653 228923 383719 228926
rect 504541 228923 504607 228926
rect 84653 228850 84719 228853
rect 206185 228850 206251 228853
rect 84653 228848 206251 228850
rect 84653 228792 84658 228848
rect 84714 228792 206190 228848
rect 206246 228792 206251 228848
rect 84653 228790 206251 228792
rect 84653 228787 84719 228790
rect 206185 228787 206251 228790
rect 246941 228850 247007 228853
rect 261385 228850 261451 228853
rect 246941 228848 261451 228850
rect 246941 228792 246946 228848
rect 247002 228792 261390 228848
rect 261446 228792 261451 228848
rect 246941 228790 261451 228792
rect 246941 228787 247007 228790
rect 261385 228787 261451 228790
rect 381537 228850 381603 228853
rect 499665 228850 499731 228853
rect 381537 228848 499731 228850
rect 381537 228792 381542 228848
rect 381598 228792 499670 228848
rect 499726 228792 499731 228848
rect 381537 228790 499731 228792
rect 381537 228787 381603 228790
rect 499665 228787 499731 228790
rect 86309 228714 86375 228717
rect 207197 228714 207263 228717
rect 86309 228712 207263 228714
rect 86309 228656 86314 228712
rect 86370 228656 207202 228712
rect 207258 228656 207263 228712
rect 86309 228654 207263 228656
rect 86309 228651 86375 228654
rect 207197 228651 207263 228654
rect 385861 228714 385927 228717
rect 509877 228714 509943 228717
rect 385861 228712 509943 228714
rect 385861 228656 385866 228712
rect 385922 228656 509882 228712
rect 509938 228656 509943 228712
rect 385861 228654 509943 228656
rect 385861 228651 385927 228654
rect 509877 228651 509943 228654
rect 88057 228578 88123 228581
rect 207565 228578 207631 228581
rect 88057 228576 207631 228578
rect 88057 228520 88062 228576
rect 88118 228520 207570 228576
rect 207626 228520 207631 228576
rect 88057 228518 207631 228520
rect 88057 228515 88123 228518
rect 207565 228515 207631 228518
rect 237097 228578 237163 228581
rect 259637 228578 259703 228581
rect 237097 228576 259703 228578
rect 237097 228520 237102 228576
rect 237158 228520 259642 228576
rect 259698 228520 259703 228576
rect 237097 228518 259703 228520
rect 237097 228515 237163 228518
rect 259637 228515 259703 228518
rect 387977 228578 388043 228581
rect 514661 228578 514727 228581
rect 387977 228576 514727 228578
rect 387977 228520 387982 228576
rect 388038 228520 514666 228576
rect 514722 228520 514727 228576
rect 387977 228518 514727 228520
rect 387977 228515 388043 228518
rect 514661 228515 514727 228518
rect 82721 228442 82787 228445
rect 205817 228442 205883 228445
rect 82721 228440 205883 228442
rect 82721 228384 82726 228440
rect 82782 228384 205822 228440
rect 205878 228384 205883 228440
rect 82721 228382 205883 228384
rect 82721 228379 82787 228382
rect 205817 228379 205883 228382
rect 235533 228442 235599 228445
rect 262489 228442 262555 228445
rect 235533 228440 262555 228442
rect 235533 228384 235538 228440
rect 235594 228384 262494 228440
rect 262550 228384 262555 228440
rect 235533 228382 262555 228384
rect 235533 228379 235599 228382
rect 262489 228379 262555 228382
rect 389081 228442 389147 228445
rect 517237 228442 517303 228445
rect 389081 228440 517303 228442
rect 389081 228384 389086 228440
rect 389142 228384 517242 228440
rect 517298 228384 517303 228440
rect 389081 228382 517303 228384
rect 389081 228379 389147 228382
rect 517237 228379 517303 228382
rect 76281 228306 76347 228309
rect 202965 228306 203031 228309
rect 76281 228304 203031 228306
rect 76281 228248 76286 228304
rect 76342 228248 202970 228304
rect 203026 228248 203031 228304
rect 76281 228246 203031 228248
rect 76281 228243 76347 228246
rect 202965 228243 203031 228246
rect 225965 228306 226031 228309
rect 266077 228306 266143 228309
rect 225965 228304 266143 228306
rect 225965 228248 225970 228304
rect 226026 228248 266082 228304
rect 266138 228248 266143 228304
rect 225965 228246 266143 228248
rect 225965 228243 226031 228246
rect 266077 228243 266143 228246
rect 391197 228306 391263 228309
rect 522481 228306 522547 228309
rect 391197 228304 522547 228306
rect 391197 228248 391202 228304
rect 391258 228248 522486 228304
rect 522542 228248 522547 228304
rect 391197 228246 522547 228248
rect 391197 228243 391263 228246
rect 522481 228243 522547 228246
rect 71221 228170 71287 228173
rect 200481 228170 200547 228173
rect 71221 228168 200547 228170
rect 71221 228112 71226 228168
rect 71282 228112 200486 228168
rect 200542 228112 200547 228168
rect 71221 228110 200547 228112
rect 71221 228107 71287 228110
rect 200481 228107 200547 228110
rect 220721 228170 220787 228173
rect 264237 228170 264303 228173
rect 220721 228168 264303 228170
rect 220721 228112 220726 228168
rect 220782 228112 264242 228168
rect 264298 228112 264303 228168
rect 220721 228110 264303 228112
rect 220721 228107 220787 228110
rect 264237 228107 264303 228110
rect 393313 228170 393379 228173
rect 527541 228170 527607 228173
rect 393313 228168 527607 228170
rect 393313 228112 393318 228168
rect 393374 228112 527546 228168
rect 527602 228112 527607 228168
rect 393313 228110 527607 228112
rect 393313 228107 393379 228110
rect 527541 228107 527607 228110
rect 69473 228034 69539 228037
rect 200113 228034 200179 228037
rect 69473 228032 200179 228034
rect 69473 227976 69478 228032
rect 69534 227976 200118 228032
rect 200174 227976 200179 228032
rect 69473 227974 200179 227976
rect 69473 227971 69539 227974
rect 200113 227971 200179 227974
rect 219249 228034 219315 228037
rect 263225 228034 263291 228037
rect 219249 228032 263291 228034
rect 219249 227976 219254 228032
rect 219310 227976 263230 228032
rect 263286 227976 263291 228032
rect 219249 227974 263291 227976
rect 219249 227971 219315 227974
rect 263225 227971 263291 227974
rect 397637 228034 397703 228037
rect 535453 228034 535519 228037
rect 397637 228032 535519 228034
rect 397637 227976 397642 228032
rect 397698 227976 535458 228032
rect 535514 227976 535519 228032
rect 397637 227974 535519 227976
rect 397637 227971 397703 227974
rect 535453 227971 535519 227974
rect 62757 227898 62823 227901
rect 197261 227898 197327 227901
rect 62757 227896 197327 227898
rect 62757 227840 62762 227896
rect 62818 227840 197266 227896
rect 197322 227840 197327 227896
rect 62757 227838 197327 227840
rect 62757 227835 62823 227838
rect 197261 227835 197327 227838
rect 217593 227898 217659 227901
rect 262857 227898 262923 227901
rect 217593 227896 262923 227898
rect 217593 227840 217598 227896
rect 217654 227840 262862 227896
rect 262918 227840 262923 227896
rect 217593 227838 262923 227840
rect 217593 227835 217659 227838
rect 262857 227835 262923 227838
rect 395429 227898 395495 227901
rect 532693 227898 532759 227901
rect 395429 227896 532759 227898
rect 395429 227840 395434 227896
rect 395490 227840 532698 227896
rect 532754 227840 532759 227896
rect 395429 227838 532759 227840
rect 395429 227835 395495 227838
rect 532693 227835 532759 227838
rect 57605 227762 57671 227765
rect 194777 227762 194843 227765
rect 57605 227760 194843 227762
rect 57605 227704 57610 227760
rect 57666 227704 194782 227760
rect 194838 227704 194843 227760
rect 57605 227702 194843 227704
rect 57605 227699 57671 227702
rect 194777 227699 194843 227702
rect 210785 227762 210851 227765
rect 260005 227762 260071 227765
rect 210785 227760 260071 227762
rect 210785 227704 210790 227760
rect 210846 227704 260010 227760
rect 260066 227704 260071 227760
rect 210785 227702 260071 227704
rect 210785 227699 210851 227702
rect 260005 227699 260071 227702
rect 402973 227762 403039 227765
rect 550265 227762 550331 227765
rect 402973 227760 550331 227762
rect 402973 227704 402978 227760
rect 403034 227704 550270 227760
rect 550326 227704 550331 227760
rect 402973 227702 550331 227704
rect 402973 227699 403039 227702
rect 550265 227699 550331 227702
rect 56041 227626 56107 227629
rect 194409 227626 194475 227629
rect 56041 227624 194475 227626
rect 56041 227568 56046 227624
rect 56102 227568 194414 227624
rect 194470 227568 194475 227624
rect 56041 227566 194475 227568
rect 56041 227563 56107 227566
rect 194409 227563 194475 227566
rect 212349 227626 212415 227629
rect 260373 227626 260439 227629
rect 212349 227624 260439 227626
rect 212349 227568 212354 227624
rect 212410 227568 260378 227624
rect 260434 227568 260439 227624
rect 212349 227566 260439 227568
rect 212349 227563 212415 227566
rect 260373 227563 260439 227566
rect 405089 227626 405155 227629
rect 555049 227626 555115 227629
rect 405089 227624 555115 227626
rect 405089 227568 405094 227624
rect 405150 227568 555054 227624
rect 555110 227568 555115 227624
rect 405089 227566 555115 227568
rect 405089 227563 405155 227566
rect 555049 227563 555115 227566
rect 94773 227490 94839 227493
rect 210417 227490 210483 227493
rect 94773 227488 210483 227490
rect 94773 227432 94778 227488
rect 94834 227432 210422 227488
rect 210478 227432 210483 227488
rect 94773 227430 210483 227432
rect 94773 227427 94839 227430
rect 210417 227427 210483 227430
rect 381169 227490 381235 227493
rect 496813 227490 496879 227493
rect 381169 227488 496879 227490
rect 381169 227432 381174 227488
rect 381230 227432 496818 227488
rect 496874 227432 496879 227488
rect 381169 227430 496879 227432
rect 381169 227427 381235 227430
rect 496813 227427 496879 227430
rect 101489 227354 101555 227357
rect 213269 227354 213335 227357
rect 101489 227352 213335 227354
rect 101489 227296 101494 227352
rect 101550 227296 213274 227352
rect 213330 227296 213335 227352
rect 101489 227294 213335 227296
rect 101489 227291 101555 227294
rect 213269 227291 213335 227294
rect 378317 227354 378383 227357
rect 492305 227354 492371 227357
rect 378317 227352 492371 227354
rect 378317 227296 378322 227352
rect 378378 227296 492310 227352
rect 492366 227296 492371 227352
rect 378317 227294 492371 227296
rect 378317 227291 378383 227294
rect 492305 227291 492371 227294
rect 99833 227218 99899 227221
rect 212901 227218 212967 227221
rect 99833 227216 212967 227218
rect 99833 227160 99838 227216
rect 99894 227160 212906 227216
rect 212962 227160 212967 227216
rect 99833 227158 212967 227160
rect 99833 227155 99899 227158
rect 212901 227155 212967 227158
rect 375833 227218 375899 227221
rect 486049 227218 486115 227221
rect 375833 227216 486115 227218
rect 375833 227160 375838 227216
rect 375894 227160 486054 227216
rect 486110 227160 486115 227216
rect 375833 227158 486115 227160
rect 375833 227155 375899 227158
rect 486049 227155 486115 227158
rect 106549 227082 106615 227085
rect 215753 227082 215819 227085
rect 106549 227080 215819 227082
rect 106549 227024 106554 227080
rect 106610 227024 215758 227080
rect 215814 227024 215819 227080
rect 106549 227022 215819 227024
rect 106549 227019 106615 227022
rect 215753 227019 215819 227022
rect 410057 227082 410123 227085
rect 516133 227082 516199 227085
rect 410057 227080 516199 227082
rect 410057 227024 410062 227080
rect 410118 227024 516138 227080
rect 516194 227024 516199 227080
rect 410057 227022 516199 227024
rect 410057 227019 410123 227022
rect 516133 227019 516199 227022
rect 113081 226946 113147 226949
rect 218605 226946 218671 226949
rect 113081 226944 218671 226946
rect 113081 226888 113086 226944
rect 113142 226888 218610 226944
rect 218666 226888 218671 226944
rect 113081 226886 218671 226888
rect 113081 226883 113147 226886
rect 218605 226883 218671 226886
rect 114921 226810 114987 226813
rect 218973 226810 219039 226813
rect 114921 226808 219039 226810
rect 114921 226752 114926 226808
rect 114982 226752 218978 226808
rect 219034 226752 219039 226808
rect 114921 226750 219039 226752
rect 114921 226747 114987 226750
rect 218973 226747 219039 226750
rect 98913 226266 98979 226269
rect 211153 226266 211219 226269
rect 98913 226264 211219 226266
rect 98913 226208 98918 226264
rect 98974 226208 211158 226264
rect 211214 226208 211219 226264
rect 98913 226206 211219 226208
rect 98913 226203 98979 226206
rect 211153 226203 211219 226206
rect 372245 226266 372311 226269
rect 478505 226266 478571 226269
rect 372245 226264 478571 226266
rect 372245 226208 372250 226264
rect 372306 226208 478510 226264
rect 478566 226208 478571 226264
rect 372245 226206 478571 226208
rect 372245 226203 372311 226206
rect 478505 226203 478571 226206
rect 102041 226130 102107 226133
rect 212533 226130 212599 226133
rect 102041 226128 212599 226130
rect 102041 226072 102046 226128
rect 102102 226072 212538 226128
rect 212594 226072 212599 226128
rect 102041 226070 212599 226072
rect 102041 226067 102107 226070
rect 212533 226067 212599 226070
rect 408309 226130 408375 226133
rect 513465 226130 513531 226133
rect 408309 226128 513531 226130
rect 408309 226072 408314 226128
rect 408370 226072 513470 226128
rect 513526 226072 513531 226128
rect 408309 226070 513531 226072
rect 408309 226067 408375 226070
rect 513465 226067 513531 226070
rect 41965 225996 42031 225997
rect 41965 225992 42012 225996
rect 42076 225994 42082 225996
rect 92197 225994 92263 225997
rect 208301 225994 208367 225997
rect 41965 225936 41970 225992
rect 41965 225932 42012 225936
rect 42076 225934 42122 225994
rect 92197 225992 208367 225994
rect 92197 225936 92202 225992
rect 92258 225936 208306 225992
rect 208362 225936 208367 225992
rect 92197 225934 208367 225936
rect 42076 225932 42082 225934
rect 41965 225931 42031 225932
rect 92197 225931 92263 225934
rect 208301 225931 208367 225934
rect 408401 225994 408467 225997
rect 518709 225994 518775 225997
rect 408401 225992 518775 225994
rect 408401 225936 408406 225992
rect 408462 225936 518714 225992
rect 518770 225936 518775 225992
rect 408401 225934 518775 225936
rect 408401 225931 408467 225934
rect 518709 225931 518775 225934
rect 80421 225858 80487 225861
rect 203701 225858 203767 225861
rect 80421 225856 203767 225858
rect 80421 225800 80426 225856
rect 80482 225800 203706 225856
rect 203762 225800 203767 225856
rect 80421 225798 203767 225800
rect 80421 225795 80487 225798
rect 203701 225795 203767 225798
rect 411161 225858 411227 225861
rect 530669 225858 530735 225861
rect 411161 225856 530735 225858
rect 411161 225800 411166 225856
rect 411222 225800 530674 225856
rect 530730 225800 530735 225856
rect 411161 225798 530735 225800
rect 411161 225795 411227 225798
rect 530669 225795 530735 225798
rect 83825 225722 83891 225725
rect 205081 225722 205147 225725
rect 83825 225720 205147 225722
rect 83825 225664 83830 225720
rect 83886 225664 205086 225720
rect 205142 225664 205147 225720
rect 83825 225662 205147 225664
rect 83825 225659 83891 225662
rect 205081 225659 205147 225662
rect 390461 225722 390527 225725
rect 520825 225722 520891 225725
rect 390461 225720 520891 225722
rect 390461 225664 390466 225720
rect 390522 225664 520830 225720
rect 520886 225664 520891 225720
rect 390461 225662 520891 225664
rect 390461 225659 390527 225662
rect 520825 225659 520891 225662
rect 77109 225586 77175 225589
rect 202229 225586 202295 225589
rect 77109 225584 202295 225586
rect 77109 225528 77114 225584
rect 77170 225528 202234 225584
rect 202290 225528 202295 225584
rect 77109 225526 202295 225528
rect 77109 225523 77175 225526
rect 202229 225523 202295 225526
rect 392577 225586 392643 225589
rect 525793 225586 525859 225589
rect 392577 225584 525859 225586
rect 392577 225528 392582 225584
rect 392638 225528 525798 225584
rect 525854 225528 525859 225584
rect 392577 225526 525859 225528
rect 392577 225523 392643 225526
rect 525793 225523 525859 225526
rect 70393 225450 70459 225453
rect 199377 225450 199443 225453
rect 70393 225448 199443 225450
rect 70393 225392 70398 225448
rect 70454 225392 199382 225448
rect 199438 225392 199443 225448
rect 70393 225390 199443 225392
rect 70393 225387 70459 225390
rect 199377 225387 199443 225390
rect 391565 225450 391631 225453
rect 523401 225450 523467 225453
rect 391565 225448 523467 225450
rect 391565 225392 391570 225448
rect 391626 225392 523406 225448
rect 523462 225392 523467 225448
rect 391565 225390 523467 225392
rect 391565 225387 391631 225390
rect 523401 225387 523467 225390
rect 66989 225314 67055 225317
rect 197997 225314 198063 225317
rect 66989 225312 198063 225314
rect 66989 225256 66994 225312
rect 67050 225256 198002 225312
rect 198058 225256 198063 225312
rect 66989 225254 198063 225256
rect 66989 225251 67055 225254
rect 197997 225251 198063 225254
rect 397913 225314 397979 225317
rect 538857 225314 538923 225317
rect 397913 225312 538923 225314
rect 397913 225256 397918 225312
rect 397974 225256 538862 225312
rect 538918 225256 538923 225312
rect 397913 225254 538923 225256
rect 397913 225251 397979 225254
rect 538857 225251 538923 225254
rect 63401 225178 63467 225181
rect 196525 225178 196591 225181
rect 63401 225176 196591 225178
rect 63401 225120 63406 225176
rect 63462 225120 196530 225176
rect 196586 225120 196591 225176
rect 63401 225118 196591 225120
rect 63401 225115 63467 225118
rect 196525 225115 196591 225118
rect 400121 225178 400187 225181
rect 543549 225178 543615 225181
rect 400121 225176 543615 225178
rect 400121 225120 400126 225176
rect 400182 225120 543554 225176
rect 543610 225120 543615 225176
rect 400121 225118 543615 225120
rect 400121 225115 400187 225118
rect 543549 225115 543615 225118
rect 55121 225042 55187 225045
rect 192569 225042 192635 225045
rect 55121 225040 192635 225042
rect 55121 224984 55126 225040
rect 55182 224984 192574 225040
rect 192630 224984 192635 225040
rect 55121 224982 192635 224984
rect 55121 224979 55187 224982
rect 192569 224979 192635 224982
rect 403341 225042 403407 225045
rect 549345 225042 549411 225045
rect 403341 225040 549411 225042
rect 403341 224984 403346 225040
rect 403402 224984 549350 225040
rect 549406 224984 549411 225040
rect 403341 224982 549411 224984
rect 403341 224979 403407 224982
rect 549345 224979 549411 224982
rect 56869 224906 56935 224909
rect 193673 224906 193739 224909
rect 56869 224904 193739 224906
rect 56869 224848 56874 224904
rect 56930 224848 193678 224904
rect 193734 224848 193739 224904
rect 56869 224846 193739 224848
rect 56869 224843 56935 224846
rect 193673 224843 193739 224846
rect 404353 224906 404419 224909
rect 552013 224906 552079 224909
rect 404353 224904 552079 224906
rect 404353 224848 404358 224904
rect 404414 224848 552018 224904
rect 552074 224848 552079 224904
rect 404353 224846 552079 224848
rect 404353 224843 404419 224846
rect 552013 224843 552079 224846
rect 97257 224770 97323 224773
rect 210509 224770 210575 224773
rect 97257 224768 210575 224770
rect 97257 224712 97262 224768
rect 97318 224712 210514 224768
rect 210570 224712 210575 224768
rect 97257 224710 210575 224712
rect 97257 224707 97323 224710
rect 210509 224707 210575 224710
rect 373717 224770 373783 224773
rect 481909 224770 481975 224773
rect 373717 224768 481975 224770
rect 373717 224712 373722 224768
rect 373778 224712 481914 224768
rect 481970 224712 481975 224768
rect 373717 224710 481975 224712
rect 373717 224707 373783 224710
rect 481909 224707 481975 224710
rect 109033 224634 109099 224637
rect 215385 224634 215451 224637
rect 109033 224632 215451 224634
rect 109033 224576 109038 224632
rect 109094 224576 215390 224632
rect 215446 224576 215451 224632
rect 109033 224574 215451 224576
rect 109033 224571 109099 224574
rect 215385 224571 215451 224574
rect 370865 224634 370931 224637
rect 475101 224634 475167 224637
rect 370865 224632 475167 224634
rect 370865 224576 370870 224632
rect 370926 224576 475106 224632
rect 475162 224576 475167 224632
rect 370865 224574 475167 224576
rect 370865 224571 370931 224574
rect 475101 224571 475167 224574
rect 112437 224498 112503 224501
rect 216857 224498 216923 224501
rect 112437 224496 216923 224498
rect 112437 224440 112442 224496
rect 112498 224440 216862 224496
rect 216918 224440 216923 224496
rect 112437 224438 216923 224440
rect 112437 224435 112503 224438
rect 216857 224435 216923 224438
rect 369393 224498 369459 224501
rect 471973 224498 472039 224501
rect 369393 224496 472039 224498
rect 369393 224440 369398 224496
rect 369454 224440 471978 224496
rect 472034 224440 472039 224496
rect 369393 224438 472039 224440
rect 369393 224435 369459 224438
rect 471973 224435 472039 224438
rect 115749 224362 115815 224365
rect 218237 224362 218303 224365
rect 115749 224360 218303 224362
rect 115749 224304 115754 224360
rect 115810 224304 218242 224360
rect 218298 224304 218303 224360
rect 115749 224302 218303 224304
rect 115749 224299 115815 224302
rect 218237 224299 218303 224302
rect 395981 224362 396047 224365
rect 480253 224362 480319 224365
rect 395981 224360 480319 224362
rect 395981 224304 395986 224360
rect 396042 224304 480258 224360
rect 480314 224304 480319 224360
rect 395981 224302 480319 224304
rect 395981 224299 396047 224302
rect 480253 224299 480319 224302
rect 110689 224226 110755 224229
rect 216489 224226 216555 224229
rect 110689 224224 216555 224226
rect 110689 224168 110694 224224
rect 110750 224168 216494 224224
rect 216550 224168 216555 224224
rect 110689 224166 216555 224168
rect 110689 224163 110755 224166
rect 216489 224163 216555 224166
rect 120809 224090 120875 224093
rect 220813 224090 220879 224093
rect 120809 224088 220879 224090
rect 120809 224032 120814 224088
rect 120870 224032 220818 224088
rect 220874 224032 220879 224088
rect 120809 224030 220879 224032
rect 120809 224027 120875 224030
rect 220813 224027 220879 224030
rect 104801 223546 104867 223549
rect 214465 223546 214531 223549
rect 104801 223544 214531 223546
rect 104801 223488 104806 223544
rect 104862 223488 214470 223544
rect 214526 223488 214531 223544
rect 104801 223486 214531 223488
rect 104801 223483 104867 223486
rect 214465 223483 214531 223486
rect 376937 223546 377003 223549
rect 488625 223546 488691 223549
rect 376937 223544 488691 223546
rect 376937 223488 376942 223544
rect 376998 223488 488630 223544
rect 488686 223488 488691 223544
rect 376937 223486 488691 223488
rect 376937 223483 377003 223486
rect 488625 223483 488691 223486
rect 675937 223546 676003 223549
rect 675937 223544 676292 223546
rect 675937 223488 675942 223544
rect 675998 223488 676292 223544
rect 675937 223486 676292 223488
rect 675937 223483 676003 223486
rect 98085 223410 98151 223413
rect 211889 223410 211955 223413
rect 98085 223408 211955 223410
rect 98085 223352 98090 223408
rect 98146 223352 211894 223408
rect 211950 223352 211955 223408
rect 98085 223350 211955 223352
rect 98085 223347 98151 223350
rect 211889 223347 211955 223350
rect 377305 223410 377371 223413
rect 489453 223410 489519 223413
rect 377305 223408 489519 223410
rect 377305 223352 377310 223408
rect 377366 223352 489458 223408
rect 489514 223352 489519 223408
rect 377305 223350 489519 223352
rect 377305 223347 377371 223350
rect 489453 223347 489519 223350
rect 96429 223274 96495 223277
rect 211521 223274 211587 223277
rect 96429 223272 211587 223274
rect 96429 223216 96434 223272
rect 96490 223216 211526 223272
rect 211582 223216 211587 223272
rect 96429 223214 211587 223216
rect 96429 223211 96495 223214
rect 211521 223211 211587 223214
rect 379789 223274 379855 223277
rect 495341 223274 495407 223277
rect 379789 223272 495407 223274
rect 379789 223216 379794 223272
rect 379850 223216 495346 223272
rect 495402 223216 495407 223272
rect 379789 223214 495407 223216
rect 379789 223211 379855 223214
rect 495341 223211 495407 223214
rect 89713 223138 89779 223141
rect 208669 223138 208735 223141
rect 89713 223136 208735 223138
rect 89713 223080 89718 223136
rect 89774 223080 208674 223136
rect 208730 223080 208735 223136
rect 89713 223078 208735 223080
rect 89713 223075 89779 223078
rect 208669 223075 208735 223078
rect 380157 223138 380223 223141
rect 494053 223138 494119 223141
rect 380157 223136 494119 223138
rect 380157 223080 380162 223136
rect 380218 223080 494058 223136
rect 494114 223080 494119 223136
rect 380157 223078 494119 223080
rect 380157 223075 380223 223078
rect 494053 223075 494119 223078
rect 675661 223138 675727 223141
rect 675661 223136 676292 223138
rect 675661 223080 675666 223136
rect 675722 223080 676292 223136
rect 675661 223078 676292 223080
rect 675661 223075 675727 223078
rect 81249 223002 81315 223005
rect 204713 223002 204779 223005
rect 81249 223000 204779 223002
rect 81249 222944 81254 223000
rect 81310 222944 204718 223000
rect 204774 222944 204779 223000
rect 81249 222942 204779 222944
rect 81249 222939 81315 222942
rect 204713 222939 204779 222942
rect 332685 223002 332751 223005
rect 381813 223002 381879 223005
rect 332685 223000 381879 223002
rect 332685 222944 332690 223000
rect 332746 222944 381818 223000
rect 381874 222944 381879 223000
rect 332685 222942 381879 222944
rect 332685 222939 332751 222942
rect 381813 222939 381879 222942
rect 384757 223002 384823 223005
rect 507117 223002 507183 223005
rect 384757 223000 507183 223002
rect 384757 222944 384762 223000
rect 384818 222944 507122 223000
rect 507178 222944 507183 223000
rect 384757 222942 507183 222944
rect 384757 222939 384823 222942
rect 507117 222939 507183 222942
rect 79593 222866 79659 222869
rect 204345 222866 204411 222869
rect 79593 222864 204411 222866
rect 79593 222808 79598 222864
rect 79654 222808 204350 222864
rect 204406 222808 204411 222864
rect 79593 222806 204411 222808
rect 79593 222803 79659 222806
rect 204345 222803 204411 222806
rect 330937 222866 331003 222869
rect 381077 222866 381143 222869
rect 330937 222864 381143 222866
rect 330937 222808 330942 222864
rect 330998 222808 381082 222864
rect 381138 222808 381143 222864
rect 330937 222806 381143 222808
rect 330937 222803 331003 222806
rect 381077 222803 381143 222806
rect 382641 222866 382707 222869
rect 502701 222866 502767 222869
rect 382641 222864 502767 222866
rect 382641 222808 382646 222864
rect 382702 222808 502706 222864
rect 502762 222808 502767 222864
rect 382641 222806 502767 222808
rect 382641 222803 382707 222806
rect 502701 222803 502767 222806
rect 72877 222730 72943 222733
rect 201493 222730 201559 222733
rect 72877 222728 201559 222730
rect 72877 222672 72882 222728
rect 72938 222672 201498 222728
rect 201554 222672 201559 222728
rect 72877 222670 201559 222672
rect 72877 222667 72943 222670
rect 201493 222667 201559 222670
rect 335813 222730 335879 222733
rect 388529 222730 388595 222733
rect 335813 222728 388595 222730
rect 335813 222672 335818 222728
rect 335874 222672 388534 222728
rect 388590 222672 388595 222728
rect 335813 222670 388595 222672
rect 335813 222667 335879 222670
rect 388529 222667 388595 222670
rect 390093 222730 390159 222733
rect 409781 222730 409847 222733
rect 510613 222730 510679 222733
rect 390093 222728 401610 222730
rect 390093 222672 390098 222728
rect 390154 222672 401610 222728
rect 390093 222670 401610 222672
rect 390093 222667 390159 222670
rect 74441 222594 74507 222597
rect 201861 222594 201927 222597
rect 74441 222592 201927 222594
rect 74441 222536 74446 222592
rect 74502 222536 201866 222592
rect 201922 222536 201927 222592
rect 74441 222534 201927 222536
rect 74441 222531 74507 222534
rect 201861 222531 201927 222534
rect 332317 222594 332383 222597
rect 384297 222594 384363 222597
rect 332317 222592 384363 222594
rect 332317 222536 332322 222592
rect 332378 222536 384302 222592
rect 384358 222536 384363 222592
rect 332317 222534 384363 222536
rect 332317 222531 332383 222534
rect 384297 222531 384363 222534
rect 392209 222594 392275 222597
rect 401550 222594 401610 222670
rect 409781 222728 510679 222730
rect 409781 222672 409786 222728
rect 409842 222672 510618 222728
rect 510674 222672 510679 222728
rect 409781 222670 510679 222672
rect 409781 222667 409847 222670
rect 510613 222667 510679 222670
rect 676029 222730 676095 222733
rect 676029 222728 676292 222730
rect 676029 222672 676034 222728
rect 676090 222672 676292 222728
rect 676029 222670 676292 222672
rect 676029 222667 676095 222670
rect 519721 222594 519787 222597
rect 392209 222592 401426 222594
rect 392209 222536 392214 222592
rect 392270 222536 401426 222592
rect 392209 222534 401426 222536
rect 401550 222592 519787 222594
rect 401550 222536 519726 222592
rect 519782 222536 519787 222592
rect 401550 222534 519787 222536
rect 392209 222531 392275 222534
rect 67817 222458 67883 222461
rect 198733 222458 198799 222461
rect 67817 222456 198799 222458
rect 67817 222400 67822 222456
rect 67878 222400 198738 222456
rect 198794 222400 198799 222456
rect 67817 222398 198799 222400
rect 67817 222395 67883 222398
rect 198733 222395 198799 222398
rect 333789 222458 333855 222461
rect 387701 222458 387767 222461
rect 333789 222456 387767 222458
rect 333789 222400 333794 222456
rect 333850 222400 387706 222456
rect 387762 222400 387767 222456
rect 333789 222398 387767 222400
rect 333789 222395 333855 222398
rect 387701 222395 387767 222398
rect 396533 222458 396599 222461
rect 401366 222458 401426 222534
rect 519721 222531 519787 222534
rect 525057 222458 525123 222461
rect 396533 222456 400230 222458
rect 396533 222400 396538 222456
rect 396594 222400 400230 222456
rect 396533 222398 400230 222400
rect 401366 222456 525123 222458
rect 401366 222400 525062 222456
rect 525118 222400 525123 222456
rect 401366 222398 525123 222400
rect 396533 222395 396599 222398
rect 61101 222322 61167 222325
rect 196157 222322 196223 222325
rect 61101 222320 196223 222322
rect 61101 222264 61106 222320
rect 61162 222264 196162 222320
rect 196218 222264 196223 222320
rect 61101 222262 196223 222264
rect 61101 222259 61167 222262
rect 196157 222259 196223 222262
rect 338757 222322 338823 222325
rect 396901 222322 396967 222325
rect 338757 222320 396967 222322
rect 338757 222264 338762 222320
rect 338818 222264 396906 222320
rect 396962 222264 396967 222320
rect 338757 222262 396967 222264
rect 400170 222322 400230 222398
rect 525057 222395 525123 222398
rect 534901 222322 534967 222325
rect 400170 222320 534967 222322
rect 400170 222264 534906 222320
rect 534962 222264 534967 222320
rect 400170 222262 534967 222264
rect 338757 222259 338823 222262
rect 396901 222259 396967 222262
rect 534901 222259 534967 222262
rect 675753 222322 675819 222325
rect 675753 222320 676292 222322
rect 675753 222264 675758 222320
rect 675814 222264 676292 222320
rect 675753 222262 676292 222264
rect 675753 222259 675819 222262
rect 54385 222186 54451 222189
rect 193305 222186 193371 222189
rect 54385 222184 193371 222186
rect 54385 222128 54390 222184
rect 54446 222128 193310 222184
rect 193366 222128 193371 222184
rect 54385 222126 193371 222128
rect 54385 222123 54451 222126
rect 193305 222123 193371 222126
rect 335905 222186 335971 222189
rect 390185 222186 390251 222189
rect 335905 222184 390251 222186
rect 335905 222128 335910 222184
rect 335966 222128 390190 222184
rect 390246 222128 390251 222184
rect 335905 222126 390251 222128
rect 335905 222123 335971 222126
rect 390185 222123 390251 222126
rect 394417 222186 394483 222189
rect 529933 222186 529999 222189
rect 394417 222184 529999 222186
rect 394417 222128 394422 222184
rect 394478 222128 529938 222184
rect 529994 222128 529999 222184
rect 394417 222126 529999 222128
rect 394417 222123 394483 222126
rect 529933 222123 529999 222126
rect 103145 222050 103211 222053
rect 214373 222050 214439 222053
rect 103145 222048 214439 222050
rect 103145 221992 103150 222048
rect 103206 221992 214378 222048
rect 214434 221992 214439 222048
rect 103145 221990 214439 221992
rect 103145 221987 103211 221990
rect 214373 221987 214439 221990
rect 375097 222050 375163 222053
rect 483565 222050 483631 222053
rect 375097 222048 483631 222050
rect 375097 221992 375102 222048
rect 375158 221992 483570 222048
rect 483626 221992 483631 222048
rect 375097 221990 483631 221992
rect 375097 221987 375163 221990
rect 483565 221987 483631 221990
rect 109861 221914 109927 221917
rect 217225 221914 217291 221917
rect 109861 221912 217291 221914
rect 109861 221856 109866 221912
rect 109922 221856 217230 221912
rect 217286 221856 217291 221912
rect 109861 221854 217291 221856
rect 109861 221851 109927 221854
rect 217225 221851 217291 221854
rect 397453 221914 397519 221917
rect 491385 221914 491451 221917
rect 397453 221912 491451 221914
rect 397453 221856 397458 221912
rect 397514 221856 491390 221912
rect 491446 221856 491451 221912
rect 397453 221854 491451 221856
rect 397453 221851 397519 221854
rect 491385 221851 491451 221854
rect 522481 221914 522547 221917
rect 627085 221914 627151 221917
rect 522481 221912 627151 221914
rect 522481 221856 522486 221912
rect 522542 221856 627090 221912
rect 627146 221856 627151 221912
rect 522481 221854 627151 221856
rect 522481 221851 522547 221854
rect 627085 221851 627151 221854
rect 675753 221914 675819 221917
rect 675753 221912 676292 221914
rect 675753 221856 675758 221912
rect 675814 221856 676292 221912
rect 675753 221854 676292 221856
rect 675753 221851 675819 221854
rect 111609 221778 111675 221781
rect 217317 221778 217383 221781
rect 111609 221776 217383 221778
rect 111609 221720 111614 221776
rect 111670 221720 217322 221776
rect 217378 221720 217383 221776
rect 111609 221718 217383 221720
rect 111609 221715 111675 221718
rect 217317 221715 217383 221718
rect 386873 221778 386939 221781
rect 409781 221778 409847 221781
rect 386873 221776 409847 221778
rect 386873 221720 386878 221776
rect 386934 221720 409786 221776
rect 409842 221720 409847 221776
rect 386873 221718 409847 221720
rect 386873 221715 386939 221718
rect 409781 221715 409847 221718
rect 510613 221778 510679 221781
rect 512453 221778 512519 221781
rect 625245 221778 625311 221781
rect 510613 221776 625311 221778
rect 510613 221720 510618 221776
rect 510674 221720 512458 221776
rect 512514 221720 625250 221776
rect 625306 221720 625311 221776
rect 510613 221718 625311 221720
rect 510613 221715 510679 221718
rect 512453 221715 512519 221718
rect 625245 221715 625311 221718
rect 121361 221642 121427 221645
rect 221825 221642 221891 221645
rect 121361 221640 221891 221642
rect 121361 221584 121366 221640
rect 121422 221584 221830 221640
rect 221886 221584 221891 221640
rect 121361 221582 221891 221584
rect 121361 221579 121427 221582
rect 221825 221579 221891 221582
rect 502701 221642 502767 221645
rect 623405 221642 623471 221645
rect 502701 221640 623471 221642
rect 502701 221584 502706 221640
rect 502762 221584 623410 221640
rect 623466 221584 623471 221640
rect 502701 221582 623471 221584
rect 502701 221579 502767 221582
rect 623405 221579 623471 221582
rect 118325 221506 118391 221509
rect 220445 221506 220511 221509
rect 118325 221504 220511 221506
rect 118325 221448 118330 221504
rect 118386 221448 220450 221504
rect 220506 221448 220511 221504
rect 118325 221446 220511 221448
rect 118325 221443 118391 221446
rect 220445 221443 220511 221446
rect 507117 221506 507183 221509
rect 624325 221506 624391 221509
rect 507117 221504 624391 221506
rect 507117 221448 507122 221504
rect 507178 221448 624330 221504
rect 624386 221448 624391 221504
rect 507117 221446 624391 221448
rect 507117 221443 507183 221446
rect 624325 221443 624391 221446
rect 675845 221506 675911 221509
rect 675845 221504 676292 221506
rect 675845 221448 675850 221504
rect 675906 221448 676292 221504
rect 675845 221446 676292 221448
rect 675845 221443 675911 221446
rect 496813 221370 496879 221373
rect 499297 221370 499363 221373
rect 622945 221370 623011 221373
rect 496813 221368 623011 221370
rect 496813 221312 496818 221368
rect 496874 221312 499302 221368
rect 499358 221312 622950 221368
rect 623006 221312 623011 221368
rect 496813 221310 623011 221312
rect 496813 221307 496879 221310
rect 499297 221307 499363 221310
rect 622945 221307 623011 221310
rect 488625 221234 488691 221237
rect 621473 221234 621539 221237
rect 488625 221232 621539 221234
rect 488625 221176 488630 221232
rect 488686 221176 621478 221232
rect 621534 221176 621539 221232
rect 488625 221174 621539 221176
rect 488625 221171 488691 221174
rect 621473 221171 621539 221174
rect 494053 221098 494119 221101
rect 496445 221098 496511 221101
rect 637389 221098 637455 221101
rect 494053 221096 637455 221098
rect 494053 221040 494058 221096
rect 494114 221040 496450 221096
rect 496506 221040 637394 221096
rect 637450 221040 637455 221096
rect 494053 221038 637455 221040
rect 494053 221035 494119 221038
rect 496445 221035 496511 221038
rect 637389 221035 637455 221038
rect 675753 221098 675819 221101
rect 675753 221096 676292 221098
rect 675753 221040 675758 221096
rect 675814 221040 676292 221096
rect 675753 221038 676292 221040
rect 675753 221035 675819 221038
rect 491385 220962 491451 220965
rect 493041 220962 493107 220965
rect 636929 220962 636995 220965
rect 491385 220960 636995 220962
rect 491385 220904 491390 220960
rect 491446 220904 493046 220960
rect 493102 220904 636934 220960
rect 636990 220904 636995 220960
rect 491385 220902 636995 220904
rect 491385 220899 491451 220902
rect 493041 220899 493107 220902
rect 636929 220899 636995 220902
rect 675569 220690 675635 220693
rect 675569 220688 676292 220690
rect 675569 220632 675574 220688
rect 675630 220632 676292 220688
rect 675569 220630 676292 220632
rect 675569 220627 675635 220630
rect 676029 220282 676095 220285
rect 676029 220280 676292 220282
rect 676029 220224 676034 220280
rect 676090 220224 676292 220280
rect 676029 220222 676292 220224
rect 676029 220219 676095 220222
rect 676070 219948 676076 220012
rect 676140 219948 676146 220012
rect 676078 219874 676138 219948
rect 676078 219814 676292 219874
rect 676029 219466 676095 219469
rect 676029 219464 676292 219466
rect 676029 219408 676034 219464
rect 676090 219408 676292 219464
rect 676029 219406 676292 219408
rect 676029 219403 676095 219406
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 675937 218650 676003 218653
rect 675937 218648 676292 218650
rect 675937 218592 675942 218648
rect 675998 218592 676292 218648
rect 675937 218590 676292 218592
rect 675937 218587 676003 218590
rect 676029 218242 676095 218245
rect 676029 218240 676292 218242
rect 676029 218184 676034 218240
rect 676090 218184 676292 218240
rect 676029 218182 676292 218184
rect 676029 218179 676095 218182
rect 676029 217834 676095 217837
rect 676029 217832 676292 217834
rect 676029 217776 676034 217832
rect 676090 217776 676292 217832
rect 676029 217774 676292 217776
rect 676029 217771 676095 217774
rect 675937 217426 676003 217429
rect 675937 217424 676292 217426
rect 675937 217368 675942 217424
rect 675998 217368 676292 217424
rect 675937 217366 676292 217368
rect 675937 217363 676003 217366
rect 675937 217018 676003 217021
rect 675937 217016 676292 217018
rect 675937 216960 675942 217016
rect 675998 216960 676292 217016
rect 675937 216958 676292 216960
rect 675937 216955 676003 216958
rect 676029 216610 676095 216613
rect 676029 216608 676292 216610
rect 676029 216552 676034 216608
rect 676090 216552 676292 216608
rect 676029 216550 676292 216552
rect 676029 216547 676095 216550
rect 580165 216202 580231 216205
rect 576380 216200 580231 216202
rect 576380 216144 580170 216200
rect 580226 216144 580231 216200
rect 576380 216142 580231 216144
rect 580165 216139 580231 216142
rect 675937 216202 676003 216205
rect 675937 216200 676292 216202
rect 675937 216144 675942 216200
rect 675998 216144 676292 216200
rect 675937 216142 676292 216144
rect 675937 216139 676003 216142
rect 675845 215794 675911 215797
rect 675845 215792 676292 215794
rect 675845 215736 675850 215792
rect 675906 215736 676292 215792
rect 675845 215734 676292 215736
rect 675845 215731 675911 215734
rect 675385 215386 675451 215389
rect 675385 215384 676292 215386
rect 675385 215328 675390 215384
rect 675446 215328 676292 215384
rect 675385 215326 676292 215328
rect 675385 215323 675451 215326
rect 41505 215114 41571 215117
rect 41462 215112 41571 215114
rect 41462 215056 41510 215112
rect 41566 215056 41571 215112
rect 41462 215051 41571 215056
rect 41462 214948 41522 215051
rect 676029 214978 676095 214981
rect 676029 214976 676292 214978
rect 676029 214920 676034 214976
rect 676090 214920 676292 214976
rect 676029 214918 676292 214920
rect 676029 214915 676095 214918
rect 41597 214706 41663 214709
rect 582281 214706 582347 214709
rect 41462 214704 41663 214706
rect 41462 214648 41602 214704
rect 41658 214648 41663 214704
rect 41462 214646 41663 214648
rect 576380 214704 582347 214706
rect 576380 214648 582286 214704
rect 582342 214648 582347 214704
rect 576380 214646 582347 214648
rect 41462 214540 41522 214646
rect 41597 214643 41663 214646
rect 582281 214643 582347 214646
rect 676029 214570 676095 214573
rect 676029 214568 676292 214570
rect 676029 214512 676034 214568
rect 676090 214512 676292 214568
rect 676029 214510 676292 214512
rect 676029 214507 676095 214510
rect 41413 214298 41479 214301
rect 41413 214296 41522 214298
rect 41413 214240 41418 214296
rect 41474 214240 41522 214296
rect 41413 214235 41522 214240
rect 41462 214132 41522 214235
rect 675937 214162 676003 214165
rect 675937 214160 676292 214162
rect 675937 214104 675942 214160
rect 675998 214104 676292 214160
rect 675937 214102 676292 214104
rect 675937 214099 676003 214102
rect 41413 213890 41479 213893
rect 41413 213888 41522 213890
rect 41413 213832 41418 213888
rect 41474 213832 41522 213888
rect 41413 213827 41522 213832
rect 41462 213724 41522 213827
rect 676029 213754 676095 213757
rect 676029 213752 676292 213754
rect 676029 213696 676034 213752
rect 676090 213696 676292 213752
rect 676029 213694 676292 213696
rect 676029 213691 676095 213694
rect 42190 213346 42196 213348
rect 41492 213286 42196 213346
rect 42190 213284 42196 213286
rect 42260 213284 42266 213348
rect 676078 213286 676292 213346
rect 580257 213210 580323 213213
rect 576380 213208 580323 213210
rect 576380 213152 580262 213208
rect 580318 213152 580323 213208
rect 576380 213150 580323 213152
rect 580257 213147 580323 213150
rect 41505 213074 41571 213077
rect 41462 213072 41571 213074
rect 41462 213016 41510 213072
rect 41566 213016 41571 213072
rect 41462 213011 41571 213016
rect 41462 212908 41522 213011
rect 46933 212530 46999 212533
rect 41492 212528 46999 212530
rect 41492 212472 46938 212528
rect 46994 212472 46999 212528
rect 41492 212470 46999 212472
rect 46933 212467 46999 212470
rect 676078 212125 676138 213286
rect 679022 212500 679082 212908
rect 45645 212122 45711 212125
rect 676029 212122 676138 212125
rect 41492 212120 45711 212122
rect 41492 212064 45650 212120
rect 45706 212064 45711 212120
rect 41492 212062 45711 212064
rect 675948 212120 676292 212122
rect 675948 212064 676034 212120
rect 676090 212064 676292 212120
rect 675948 212062 676292 212064
rect 45645 212059 45711 212062
rect 676029 212059 676095 212062
rect 41822 211714 41828 211716
rect 41492 211654 41828 211714
rect 41822 211652 41828 211654
rect 41892 211652 41898 211716
rect 581637 211714 581703 211717
rect 576380 211712 581703 211714
rect 576380 211656 581642 211712
rect 581698 211656 581703 211712
rect 576380 211654 581703 211656
rect 581637 211651 581703 211654
rect 45461 211306 45527 211309
rect 41492 211304 45527 211306
rect 41492 211248 45466 211304
rect 45522 211248 45527 211304
rect 41492 211246 45527 211248
rect 45461 211243 45527 211246
rect 41454 210972 41460 211036
rect 41524 210972 41530 211036
rect 41462 210868 41522 210972
rect 42742 210490 42748 210492
rect 41492 210430 42748 210490
rect 42742 210428 42748 210430
rect 42812 210428 42818 210492
rect 580533 210218 580599 210221
rect 576380 210216 580599 210218
rect 576380 210160 580538 210216
rect 580594 210160 580599 210216
rect 576380 210158 580599 210160
rect 580533 210155 580599 210158
rect 32998 209813 33058 210052
rect 32949 209808 33058 209813
rect 32949 209752 32954 209808
rect 33010 209752 33058 209808
rect 32949 209750 33058 209752
rect 32949 209747 33015 209750
rect 41822 209674 41828 209676
rect 41492 209614 41828 209674
rect 41822 209612 41828 209614
rect 41892 209612 41898 209676
rect 599761 209538 599827 209541
rect 599761 209536 606556 209538
rect 599761 209480 599766 209536
rect 599822 209480 606556 209536
rect 599761 209478 606556 209480
rect 599761 209475 599827 209478
rect 42374 209266 42380 209268
rect 41492 209206 42380 209266
rect 42374 209204 42380 209206
rect 42444 209204 42450 209268
rect 671061 209266 671127 209269
rect 666356 209264 671127 209266
rect 666356 209208 671066 209264
rect 671122 209208 671127 209264
rect 666356 209206 671127 209208
rect 671061 209203 671127 209206
rect 42558 208858 42564 208860
rect 41492 208798 42564 208858
rect 42558 208796 42564 208798
rect 42628 208796 42634 208860
rect 579705 208722 579771 208725
rect 576380 208720 579771 208722
rect 576380 208664 579710 208720
rect 579766 208664 579771 208720
rect 576380 208662 579771 208664
rect 579705 208659 579771 208662
rect 599945 208586 600011 208589
rect 599945 208584 606556 208586
rect 599945 208528 599950 208584
rect 600006 208528 606556 208584
rect 599945 208526 606556 208528
rect 599945 208523 600011 208526
rect 32998 208181 33058 208420
rect 32998 208176 33107 208181
rect 32998 208120 33046 208176
rect 33102 208120 33107 208176
rect 32998 208118 33107 208120
rect 33041 208115 33107 208118
rect 41462 207770 41522 208012
rect 41638 207770 41644 207772
rect 41462 207710 41644 207770
rect 41638 207708 41644 207710
rect 41708 207708 41714 207772
rect 42006 207634 42012 207636
rect 41492 207574 42012 207634
rect 42006 207572 42012 207574
rect 42076 207572 42082 207636
rect 599853 207498 599919 207501
rect 599853 207496 606556 207498
rect 599853 207440 599858 207496
rect 599914 207440 606556 207496
rect 599853 207438 606556 207440
rect 599853 207435 599919 207438
rect 42190 207226 42196 207228
rect 41492 207166 42196 207226
rect 42190 207164 42196 207166
rect 42260 207164 42266 207228
rect 582281 207090 582347 207093
rect 576380 207088 582347 207090
rect 576380 207032 582286 207088
rect 582342 207032 582347 207088
rect 576380 207030 582347 207032
rect 582281 207027 582347 207030
rect 42885 206818 42951 206821
rect 41492 206816 42951 206818
rect 41492 206760 42890 206816
rect 42946 206760 42951 206816
rect 41492 206758 42951 206760
rect 42885 206755 42951 206758
rect 600037 206546 600103 206549
rect 600037 206544 606556 206546
rect 600037 206488 600042 206544
rect 600098 206488 606556 206544
rect 600037 206486 606556 206488
rect 600037 206483 600103 206486
rect 43069 206410 43135 206413
rect 41492 206408 43135 206410
rect 41492 206352 43074 206408
rect 43130 206352 43135 206408
rect 41492 206350 43135 206352
rect 43069 206347 43135 206350
rect 675569 206002 675635 206005
rect 674606 206000 675635 206002
rect 41462 205732 41522 205972
rect 674606 205944 675574 206000
rect 675630 205944 675635 206000
rect 674606 205942 675635 205944
rect 671061 205866 671127 205869
rect 666356 205864 671127 205866
rect 666356 205808 671066 205864
rect 671122 205808 671127 205864
rect 666356 205806 671127 205808
rect 671061 205803 671127 205806
rect 41454 205668 41460 205732
rect 41524 205668 41530 205732
rect 42977 205594 43043 205597
rect 582281 205594 582347 205597
rect 41492 205592 43043 205594
rect 41492 205536 42982 205592
rect 43038 205536 43043 205592
rect 41492 205534 43043 205536
rect 576380 205592 582347 205594
rect 576380 205536 582286 205592
rect 582342 205536 582347 205592
rect 576380 205534 582347 205536
rect 42977 205531 43043 205534
rect 582281 205531 582347 205534
rect 599117 205458 599183 205461
rect 599117 205456 606556 205458
rect 599117 205400 599122 205456
rect 599178 205400 606556 205456
rect 599117 205398 606556 205400
rect 599117 205395 599183 205398
rect 42793 205186 42859 205189
rect 41492 205184 42859 205186
rect 41492 205128 42798 205184
rect 42854 205128 42859 205184
rect 41492 205126 42859 205128
rect 42793 205123 42859 205126
rect 674465 205050 674531 205053
rect 674606 205050 674666 205942
rect 675569 205939 675635 205942
rect 674465 205048 674666 205050
rect 674465 204992 674470 205048
rect 674526 204992 674666 205048
rect 674465 204990 674666 204992
rect 674465 204987 674531 204990
rect 48221 204778 48287 204781
rect 41492 204776 48287 204778
rect 41492 204720 48226 204776
rect 48282 204720 48287 204776
rect 41492 204718 48287 204720
rect 48221 204715 48287 204718
rect 29177 204506 29243 204509
rect 29134 204504 29243 204506
rect 29134 204448 29182 204504
rect 29238 204448 29243 204504
rect 29134 204443 29243 204448
rect 601509 204506 601575 204509
rect 601509 204504 606556 204506
rect 601509 204448 601514 204504
rect 601570 204448 606556 204504
rect 601509 204446 606556 204448
rect 601509 204443 601575 204446
rect 29134 204340 29194 204443
rect 670969 204234 671035 204237
rect 666356 204232 671035 204234
rect 666356 204176 670974 204232
rect 671030 204176 671035 204232
rect 666356 204174 671035 204176
rect 670969 204171 671035 204174
rect 580717 204098 580783 204101
rect 576380 204096 580783 204098
rect 576380 204040 580722 204096
rect 580778 204040 580783 204096
rect 576380 204038 580783 204040
rect 580717 204035 580783 204038
rect 31661 203690 31727 203693
rect 31661 203688 31770 203690
rect 31661 203632 31666 203688
rect 31722 203632 31770 203688
rect 31661 203627 31770 203632
rect 31710 203524 31770 203627
rect 601417 203418 601483 203421
rect 601417 203416 606556 203418
rect 601417 203360 601422 203416
rect 601478 203360 606556 203416
rect 601417 203358 606556 203360
rect 601417 203355 601483 203358
rect 581085 202602 581151 202605
rect 576380 202600 581151 202602
rect 576380 202544 581090 202600
rect 581146 202544 581151 202600
rect 576380 202542 581151 202544
rect 581085 202539 581151 202542
rect 599945 202466 600011 202469
rect 599945 202464 606556 202466
rect 599945 202408 599950 202464
rect 600006 202408 606556 202464
rect 599945 202406 606556 202408
rect 599945 202403 600011 202406
rect 598933 201378 598999 201381
rect 598933 201376 606556 201378
rect 598933 201320 598938 201376
rect 598994 201320 606556 201376
rect 598933 201318 606556 201320
rect 598933 201315 598999 201318
rect 581085 201106 581151 201109
rect 576380 201104 581151 201106
rect 576380 201048 581090 201104
rect 581146 201048 581151 201104
rect 576380 201046 581151 201048
rect 581085 201043 581151 201046
rect 670969 200834 671035 200837
rect 666356 200832 671035 200834
rect 666356 200776 670974 200832
rect 671030 200776 671035 200832
rect 666356 200774 671035 200776
rect 670969 200771 671035 200774
rect 599945 200426 600011 200429
rect 599945 200424 606556 200426
rect 599945 200368 599950 200424
rect 600006 200368 606556 200424
rect 599945 200366 606556 200368
rect 599945 200363 600011 200366
rect 582281 199610 582347 199613
rect 576380 199608 582347 199610
rect 576380 199552 582286 199608
rect 582342 199552 582347 199608
rect 576380 199550 582347 199552
rect 582281 199547 582347 199550
rect 599945 199338 600011 199341
rect 599945 199336 606556 199338
rect 599945 199280 599950 199336
rect 600006 199280 606556 199336
rect 599945 199278 606556 199280
rect 599945 199275 600011 199278
rect 670877 199066 670943 199069
rect 666356 199064 670943 199066
rect 666356 199008 670882 199064
rect 670938 199008 670943 199064
rect 666356 199006 670943 199008
rect 670877 199003 670943 199006
rect 599117 198386 599183 198389
rect 599117 198384 606556 198386
rect 599117 198328 599122 198384
rect 599178 198328 606556 198384
rect 599117 198326 606556 198328
rect 599117 198323 599183 198326
rect 582281 197978 582347 197981
rect 576380 197976 582347 197978
rect 576380 197920 582286 197976
rect 582342 197920 582347 197976
rect 576380 197918 582347 197920
rect 582281 197915 582347 197918
rect 599945 197298 600011 197301
rect 599945 197296 606556 197298
rect 599945 197240 599950 197296
rect 600006 197240 606556 197296
rect 599945 197238 606556 197240
rect 599945 197235 600011 197238
rect 580717 196482 580783 196485
rect 576380 196480 580783 196482
rect 576380 196424 580722 196480
rect 580778 196424 580783 196480
rect 576380 196422 580783 196424
rect 580717 196419 580783 196422
rect 599853 196346 599919 196349
rect 599853 196344 606556 196346
rect 599853 196288 599858 196344
rect 599914 196288 606556 196344
rect 599853 196286 606556 196288
rect 599853 196283 599919 196286
rect 670877 195666 670943 195669
rect 666356 195664 670943 195666
rect 666356 195608 670882 195664
rect 670938 195608 670943 195664
rect 666356 195606 670943 195608
rect 670877 195603 670943 195606
rect 599945 195258 600011 195261
rect 599945 195256 606556 195258
rect 599945 195200 599950 195256
rect 600006 195200 606556 195256
rect 599945 195198 606556 195200
rect 599945 195195 600011 195198
rect 582281 194986 582347 194989
rect 576380 194984 582347 194986
rect 576380 194928 582286 194984
rect 582342 194928 582347 194984
rect 576380 194926 582347 194928
rect 582281 194923 582347 194926
rect 599117 194306 599183 194309
rect 599117 194304 606556 194306
rect 599117 194248 599122 194304
rect 599178 194248 606556 194304
rect 599117 194246 606556 194248
rect 599117 194243 599183 194246
rect 670785 194034 670851 194037
rect 666356 194032 670851 194034
rect 666356 193976 670790 194032
rect 670846 193976 670851 194032
rect 666356 193974 670851 193976
rect 670785 193971 670851 193974
rect 582189 193490 582255 193493
rect 576380 193488 582255 193490
rect 576380 193432 582194 193488
rect 582250 193432 582255 193488
rect 576380 193430 582255 193432
rect 582189 193427 582255 193430
rect 599945 193218 600011 193221
rect 599945 193216 606556 193218
rect 599945 193160 599950 193216
rect 600006 193160 606556 193216
rect 599945 193158 606556 193160
rect 599945 193155 600011 193158
rect 599117 192266 599183 192269
rect 599117 192264 606556 192266
rect 599117 192208 599122 192264
rect 599178 192208 606556 192264
rect 599117 192206 606556 192208
rect 599117 192203 599183 192206
rect 582281 191994 582347 191997
rect 576380 191992 582347 191994
rect 576380 191936 582286 191992
rect 582342 191936 582347 191992
rect 576380 191934 582347 191936
rect 582281 191931 582347 191934
rect 599853 191178 599919 191181
rect 599853 191176 606556 191178
rect 599853 191120 599858 191176
rect 599914 191120 606556 191176
rect 599853 191118 606556 191120
rect 599853 191115 599919 191118
rect 670785 190634 670851 190637
rect 666356 190632 670851 190634
rect 666356 190576 670790 190632
rect 670846 190576 670851 190632
rect 666356 190574 670851 190576
rect 670785 190571 670851 190574
rect 582189 190498 582255 190501
rect 576380 190496 582255 190498
rect 576380 190440 582194 190496
rect 582250 190440 582255 190496
rect 576380 190438 582255 190440
rect 582189 190435 582255 190438
rect 42149 190226 42215 190229
rect 42558 190226 42564 190228
rect 42149 190224 42564 190226
rect 42149 190168 42154 190224
rect 42210 190168 42564 190224
rect 42149 190166 42564 190168
rect 42149 190163 42215 190166
rect 42558 190164 42564 190166
rect 42628 190164 42634 190228
rect 600957 190226 601023 190229
rect 600957 190224 606556 190226
rect 600957 190168 600962 190224
rect 601018 190168 606556 190224
rect 600957 190166 606556 190168
rect 600957 190163 601023 190166
rect 601601 189138 601667 189141
rect 601601 189136 606556 189138
rect 601601 189080 601606 189136
rect 601662 189080 606556 189136
rect 601601 189078 606556 189080
rect 601601 189075 601667 189078
rect 670693 189002 670759 189005
rect 666356 189000 670759 189002
rect 666356 188944 670698 189000
rect 670754 188944 670759 189000
rect 666356 188942 670759 188944
rect 670693 188939 670759 188942
rect 579797 188866 579863 188869
rect 576380 188864 579863 188866
rect 576380 188808 579802 188864
rect 579858 188808 579863 188864
rect 576380 188806 579863 188808
rect 579797 188803 579863 188806
rect 601417 188186 601483 188189
rect 601417 188184 606556 188186
rect 601417 188128 601422 188184
rect 601478 188128 606556 188184
rect 601417 188126 606556 188128
rect 601417 188123 601483 188126
rect 41454 187580 41460 187644
rect 41524 187642 41530 187644
rect 41873 187642 41939 187645
rect 41524 187640 41939 187642
rect 41524 187584 41878 187640
rect 41934 187584 41939 187640
rect 41524 187582 41939 187584
rect 41524 187580 41530 187582
rect 41873 187579 41939 187582
rect 582281 187370 582347 187373
rect 576380 187368 582347 187370
rect 576380 187312 582286 187368
rect 582342 187312 582347 187368
rect 576380 187310 582347 187312
rect 582281 187307 582347 187310
rect 42149 187100 42215 187101
rect 42149 187098 42196 187100
rect 42104 187096 42196 187098
rect 42104 187040 42154 187096
rect 42104 187038 42196 187040
rect 42149 187036 42196 187038
rect 42260 187036 42266 187100
rect 599945 187098 600011 187101
rect 599945 187096 606556 187098
rect 599945 187040 599950 187096
rect 600006 187040 606556 187096
rect 599945 187038 606556 187040
rect 42149 187035 42215 187036
rect 599945 187035 600011 187038
rect 41965 186420 42031 186421
rect 41965 186416 42012 186420
rect 42076 186418 42082 186420
rect 41965 186360 41970 186416
rect 41965 186356 42012 186360
rect 42076 186358 42122 186418
rect 42076 186356 42082 186358
rect 41965 186355 42031 186356
rect 600037 186146 600103 186149
rect 600037 186144 606556 186146
rect 600037 186088 600042 186144
rect 600098 186088 606556 186144
rect 600037 186086 606556 186088
rect 600037 186083 600103 186086
rect 42149 185874 42215 185877
rect 42374 185874 42380 185876
rect 42149 185872 42380 185874
rect 42149 185816 42154 185872
rect 42210 185816 42380 185872
rect 42149 185814 42380 185816
rect 42149 185811 42215 185814
rect 42374 185812 42380 185814
rect 42444 185812 42450 185876
rect 582189 185874 582255 185877
rect 576380 185872 582255 185874
rect 576380 185816 582194 185872
rect 582250 185816 582255 185872
rect 576380 185814 582255 185816
rect 582189 185811 582255 185814
rect 670693 185602 670759 185605
rect 666356 185600 670759 185602
rect 666356 185544 670698 185600
rect 670754 185544 670759 185600
rect 666356 185542 670759 185544
rect 670693 185539 670759 185542
rect 599853 185058 599919 185061
rect 599853 185056 606556 185058
rect 599853 185000 599858 185056
rect 599914 185000 606556 185056
rect 599853 184998 606556 185000
rect 599853 184995 599919 184998
rect 580901 184378 580967 184381
rect 576380 184376 580967 184378
rect 576380 184320 580906 184376
rect 580962 184320 580967 184376
rect 576380 184318 580967 184320
rect 580901 184315 580967 184318
rect 42149 184242 42215 184245
rect 42742 184242 42748 184244
rect 42149 184240 42748 184242
rect 42149 184184 42154 184240
rect 42210 184184 42748 184240
rect 42149 184182 42748 184184
rect 42149 184179 42215 184182
rect 42742 184180 42748 184182
rect 42812 184180 42818 184244
rect 599761 184106 599827 184109
rect 599761 184104 606556 184106
rect 599761 184048 599766 184104
rect 599822 184048 606556 184104
rect 599761 184046 606556 184048
rect 599761 184043 599827 184046
rect 666645 183834 666711 183837
rect 672073 183834 672139 183837
rect 666356 183832 672139 183834
rect 666356 183776 666650 183832
rect 666706 183776 672078 183832
rect 672134 183776 672139 183832
rect 666356 183774 672139 183776
rect 666645 183771 666711 183774
rect 672073 183771 672139 183774
rect 41638 183636 41644 183700
rect 41708 183698 41714 183700
rect 41781 183698 41847 183701
rect 41708 183696 41847 183698
rect 41708 183640 41786 183696
rect 41842 183640 41847 183696
rect 41708 183638 41847 183640
rect 41708 183636 41714 183638
rect 41781 183635 41847 183638
rect 599945 183018 600011 183021
rect 599945 183016 606556 183018
rect 599945 182960 599950 183016
rect 600006 182960 606556 183016
rect 599945 182958 606556 182960
rect 599945 182955 600011 182958
rect 580257 182882 580323 182885
rect 576380 182880 580323 182882
rect 576380 182824 580262 182880
rect 580318 182824 580323 182880
rect 576380 182822 580323 182824
rect 580257 182819 580323 182822
rect 41781 182748 41847 182749
rect 41781 182744 41828 182748
rect 41892 182746 41898 182748
rect 41781 182688 41786 182744
rect 41781 182684 41828 182688
rect 41892 182686 41938 182746
rect 41892 182684 41898 182686
rect 41781 182683 41847 182684
rect 600037 182066 600103 182069
rect 600037 182064 606556 182066
rect 600037 182008 600042 182064
rect 600098 182008 606556 182064
rect 600037 182006 606556 182008
rect 600037 182003 600103 182006
rect 580625 181386 580691 181389
rect 576380 181384 580691 181386
rect 576380 181328 580630 181384
rect 580686 181328 580691 181384
rect 576380 181326 580691 181328
rect 580625 181323 580691 181326
rect 600129 180978 600195 180981
rect 600129 180976 606556 180978
rect 600129 180920 600134 180976
rect 600190 180920 606556 180976
rect 600129 180918 606556 180920
rect 600129 180915 600195 180918
rect 666645 180434 666711 180437
rect 666356 180432 666711 180434
rect 666356 180376 666650 180432
rect 666706 180376 666711 180432
rect 666356 180374 666711 180376
rect 666645 180371 666711 180374
rect 599853 180026 599919 180029
rect 599853 180024 606556 180026
rect 599853 179968 599858 180024
rect 599914 179968 606556 180024
rect 599853 179966 606556 179968
rect 599853 179963 599919 179966
rect 580533 179754 580599 179757
rect 576380 179752 580599 179754
rect 576380 179696 580538 179752
rect 580594 179696 580599 179752
rect 576380 179694 580599 179696
rect 580533 179691 580599 179694
rect 703813 179210 703879 179213
rect 708965 179210 709031 179213
rect 703813 179150 709031 179210
rect 703813 179147 703879 179150
rect 708965 179147 709031 179150
rect 599669 178938 599735 178941
rect 599669 178936 606556 178938
rect 599669 178880 599674 178936
rect 599730 178880 606556 178936
rect 599669 178878 606556 178880
rect 599669 178875 599735 178878
rect 666645 178802 666711 178805
rect 672165 178802 672231 178805
rect 666356 178800 672231 178802
rect 666356 178744 666650 178800
rect 666706 178744 672170 178800
rect 672226 178744 672231 178800
rect 666356 178742 672231 178744
rect 666645 178739 666711 178742
rect 672165 178739 672231 178742
rect 675753 178530 675819 178533
rect 675753 178528 676292 178530
rect 675753 178472 675758 178528
rect 675814 178472 676292 178528
rect 675753 178470 676292 178472
rect 675753 178467 675819 178470
rect 581085 178258 581151 178261
rect 576380 178256 581151 178258
rect 576380 178200 581090 178256
rect 581146 178200 581151 178256
rect 576380 178198 581151 178200
rect 581085 178195 581151 178198
rect 675937 178122 676003 178125
rect 675937 178120 676292 178122
rect 675937 178064 675942 178120
rect 675998 178064 676292 178120
rect 675937 178062 676292 178064
rect 675937 178059 676003 178062
rect 599761 177986 599827 177989
rect 599761 177984 606556 177986
rect 599761 177928 599766 177984
rect 599822 177928 606556 177984
rect 599761 177926 606556 177928
rect 599761 177923 599827 177926
rect 676029 177714 676095 177717
rect 676029 177712 676292 177714
rect 676029 177656 676034 177712
rect 676090 177656 676292 177712
rect 676029 177654 676292 177656
rect 676029 177651 676095 177654
rect 675845 177306 675911 177309
rect 675845 177304 676292 177306
rect 675845 177248 675850 177304
rect 675906 177248 676292 177304
rect 675845 177246 676292 177248
rect 675845 177243 675911 177246
rect 598933 176898 598999 176901
rect 675937 176898 676003 176901
rect 598933 176896 606556 176898
rect 598933 176840 598938 176896
rect 598994 176840 606556 176896
rect 598933 176838 606556 176840
rect 675937 176896 676292 176898
rect 675937 176840 675942 176896
rect 675998 176840 676292 176896
rect 675937 176838 676292 176840
rect 598933 176835 598999 176838
rect 675937 176835 676003 176838
rect 580717 176762 580783 176765
rect 576380 176760 580783 176762
rect 576380 176704 580722 176760
rect 580778 176704 580783 176760
rect 576380 176702 580783 176704
rect 580717 176699 580783 176702
rect 676029 176490 676095 176493
rect 676029 176488 676292 176490
rect 676029 176432 676034 176488
rect 676090 176432 676292 176488
rect 676029 176430 676292 176432
rect 676029 176427 676095 176430
rect 675937 176082 676003 176085
rect 675937 176080 676292 176082
rect 675937 176024 675942 176080
rect 675998 176024 676292 176080
rect 675937 176022 676292 176024
rect 675937 176019 676003 176022
rect 600313 175946 600379 175949
rect 600313 175944 606556 175946
rect 600313 175888 600318 175944
rect 600374 175888 606556 175944
rect 600313 175886 606556 175888
rect 600313 175883 600379 175886
rect 676029 175674 676095 175677
rect 676029 175672 676292 175674
rect 676029 175616 676034 175672
rect 676090 175616 676292 175672
rect 676029 175614 676292 175616
rect 676029 175611 676095 175614
rect 666645 175402 666711 175405
rect 666356 175400 666711 175402
rect 666356 175344 666650 175400
rect 666706 175344 666711 175400
rect 666356 175342 666711 175344
rect 666645 175339 666711 175342
rect 581453 175266 581519 175269
rect 576380 175264 581519 175266
rect 576380 175208 581458 175264
rect 581514 175208 581519 175264
rect 576380 175206 581519 175208
rect 581453 175203 581519 175206
rect 675937 175266 676003 175269
rect 675937 175264 676292 175266
rect 675937 175208 675942 175264
rect 675998 175208 676292 175264
rect 675937 175206 676292 175208
rect 675937 175203 676003 175206
rect 599945 174858 600011 174861
rect 676029 174858 676095 174861
rect 599945 174856 606556 174858
rect 599945 174800 599950 174856
rect 600006 174800 606556 174856
rect 599945 174798 606556 174800
rect 676029 174856 676292 174858
rect 676029 174800 676034 174856
rect 676090 174800 676292 174856
rect 676029 174798 676292 174800
rect 599945 174795 600011 174798
rect 676029 174795 676095 174798
rect 676029 174450 676095 174453
rect 676029 174448 676292 174450
rect 676029 174392 676034 174448
rect 676090 174392 676292 174448
rect 676029 174390 676292 174392
rect 676029 174387 676095 174390
rect 676029 174042 676095 174045
rect 676029 174040 676292 174042
rect 676029 173984 676034 174040
rect 676090 173984 676292 174040
rect 676029 173982 676292 173984
rect 676029 173979 676095 173982
rect 601141 173906 601207 173909
rect 601141 173904 606556 173906
rect 601141 173848 601146 173904
rect 601202 173848 606556 173904
rect 601141 173846 606556 173848
rect 601141 173843 601207 173846
rect 582281 173770 582347 173773
rect 576380 173768 582347 173770
rect 576380 173712 582286 173768
rect 582342 173712 582347 173768
rect 576380 173710 582347 173712
rect 582281 173707 582347 173710
rect 666645 173634 666711 173637
rect 671797 173634 671863 173637
rect 666356 173632 671863 173634
rect 666356 173576 666650 173632
rect 666706 173576 671802 173632
rect 671858 173576 671863 173632
rect 666356 173574 671863 173576
rect 666645 173571 666711 173574
rect 671797 173571 671863 173574
rect 675886 173572 675892 173636
rect 675956 173634 675962 173636
rect 675956 173574 676292 173634
rect 675956 173572 675962 173574
rect 675753 173226 675819 173229
rect 675753 173224 676292 173226
rect 675753 173168 675758 173224
rect 675814 173168 676292 173224
rect 675753 173166 676292 173168
rect 675753 173163 675819 173166
rect 599853 172818 599919 172821
rect 676029 172818 676095 172821
rect 599853 172816 606556 172818
rect 599853 172760 599858 172816
rect 599914 172760 606556 172816
rect 599853 172758 606556 172760
rect 676029 172816 676292 172818
rect 676029 172760 676034 172816
rect 676090 172760 676292 172816
rect 676029 172758 676292 172760
rect 599853 172755 599919 172758
rect 676029 172755 676095 172758
rect 675937 172410 676003 172413
rect 675937 172408 676292 172410
rect 675937 172352 675942 172408
rect 675998 172352 676292 172408
rect 675937 172350 676292 172352
rect 675937 172347 676003 172350
rect 579705 172274 579771 172277
rect 576380 172272 579771 172274
rect 576380 172216 579710 172272
rect 579766 172216 579771 172272
rect 576380 172214 579771 172216
rect 579705 172211 579771 172214
rect 676078 171942 676292 172002
rect 599945 171866 600011 171869
rect 676078 171868 676138 171942
rect 599945 171864 606556 171866
rect 599945 171808 599950 171864
rect 600006 171808 606556 171864
rect 599945 171806 606556 171808
rect 599945 171803 600011 171806
rect 676070 171804 676076 171868
rect 676140 171804 676146 171868
rect 676029 171594 676095 171597
rect 676029 171592 676292 171594
rect 676029 171536 676034 171592
rect 676090 171536 676292 171592
rect 676029 171534 676292 171536
rect 676029 171531 676095 171534
rect 675937 171186 676003 171189
rect 675937 171184 676292 171186
rect 675937 171128 675942 171184
rect 675998 171128 676292 171184
rect 675937 171126 676292 171128
rect 675937 171123 676003 171126
rect 599945 170778 600011 170781
rect 599945 170776 606556 170778
rect 599945 170720 599950 170776
rect 600006 170720 606556 170776
rect 599945 170718 606556 170720
rect 599945 170715 600011 170718
rect 675702 170716 675708 170780
rect 675772 170778 675778 170780
rect 675772 170718 676292 170778
rect 675772 170716 675778 170718
rect 580533 170642 580599 170645
rect 576380 170640 580599 170642
rect 576380 170584 580538 170640
rect 580594 170584 580599 170640
rect 576380 170582 580599 170584
rect 580533 170579 580599 170582
rect 675937 170370 676003 170373
rect 675937 170368 676292 170370
rect 675937 170312 675942 170368
rect 675998 170312 676292 170368
rect 675937 170310 676292 170312
rect 675937 170307 676003 170310
rect 666645 170234 666711 170237
rect 666356 170232 666711 170234
rect 666356 170176 666650 170232
rect 666706 170176 666711 170232
rect 666356 170174 666711 170176
rect 666645 170171 666711 170174
rect 675937 169962 676003 169965
rect 675937 169960 676292 169962
rect 675937 169904 675942 169960
rect 675998 169904 676292 169960
rect 675937 169902 676292 169904
rect 675937 169899 676003 169902
rect 599761 169826 599827 169829
rect 599761 169824 606556 169826
rect 599761 169768 599766 169824
rect 599822 169768 606556 169824
rect 599761 169766 606556 169768
rect 599761 169763 599827 169766
rect 676029 169554 676095 169557
rect 676029 169552 676292 169554
rect 676029 169496 676034 169552
rect 676090 169496 676292 169552
rect 676029 169494 676292 169496
rect 676029 169491 676095 169494
rect 582005 169146 582071 169149
rect 576380 169144 582071 169146
rect 576380 169088 582010 169144
rect 582066 169088 582071 169144
rect 576380 169086 582071 169088
rect 582005 169083 582071 169086
rect 675937 169146 676003 169149
rect 675937 169144 676292 169146
rect 675937 169088 675942 169144
rect 675998 169088 676292 169144
rect 675937 169086 676292 169088
rect 675937 169083 676003 169086
rect 599025 168738 599091 168741
rect 675845 168738 675911 168741
rect 599025 168736 606556 168738
rect 599025 168680 599030 168736
rect 599086 168680 606556 168736
rect 599025 168678 606556 168680
rect 675845 168736 676292 168738
rect 675845 168680 675850 168736
rect 675906 168680 676292 168736
rect 675845 168678 676292 168680
rect 599025 168675 599091 168678
rect 675845 168675 675911 168678
rect 666645 168602 666711 168605
rect 672349 168602 672415 168605
rect 666356 168600 672415 168602
rect 666356 168544 666650 168600
rect 666706 168544 672354 168600
rect 672410 168544 672415 168600
rect 666356 168542 672415 168544
rect 666645 168539 666711 168542
rect 672349 168539 672415 168542
rect 676029 168330 676095 168333
rect 676029 168328 676292 168330
rect 676029 168272 676034 168328
rect 676090 168272 676292 168328
rect 676029 168270 676292 168272
rect 676029 168267 676095 168270
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 599853 167786 599919 167789
rect 599853 167784 606556 167786
rect 599853 167728 599858 167784
rect 599914 167728 606556 167784
rect 599853 167726 606556 167728
rect 599853 167723 599919 167726
rect 580993 167650 581059 167653
rect 576380 167648 581059 167650
rect 576380 167592 580998 167648
rect 581054 167592 581059 167648
rect 576380 167590 581059 167592
rect 580993 167587 581059 167590
rect 676029 167106 676095 167109
rect 676029 167104 676292 167106
rect 676029 167048 676034 167104
rect 676090 167048 676292 167104
rect 676029 167046 676292 167048
rect 676029 167043 676095 167046
rect 600037 166698 600103 166701
rect 600037 166696 606556 166698
rect 600037 166640 600042 166696
rect 600098 166640 606556 166696
rect 600037 166638 606556 166640
rect 600037 166635 600103 166638
rect 582281 166154 582347 166157
rect 576380 166152 582347 166154
rect 576380 166096 582286 166152
rect 582342 166096 582347 166152
rect 576380 166094 582347 166096
rect 582281 166091 582347 166094
rect 599945 165746 600011 165749
rect 599945 165744 606556 165746
rect 599945 165688 599950 165744
rect 600006 165688 606556 165744
rect 599945 165686 606556 165688
rect 599945 165683 600011 165686
rect 666645 165202 666711 165205
rect 666356 165200 666711 165202
rect 666356 165144 666650 165200
rect 666706 165144 666711 165200
rect 666356 165142 666711 165144
rect 666645 165139 666711 165142
rect 580809 164658 580875 164661
rect 576380 164656 580875 164658
rect 576380 164600 580814 164656
rect 580870 164600 580875 164656
rect 576380 164598 580875 164600
rect 580809 164595 580875 164598
rect 599853 164658 599919 164661
rect 599853 164656 606556 164658
rect 599853 164600 599858 164656
rect 599914 164600 606556 164656
rect 599853 164598 606556 164600
rect 599853 164595 599919 164598
rect 599945 163706 600011 163709
rect 599945 163704 606556 163706
rect 599945 163648 599950 163704
rect 600006 163648 606556 163704
rect 599945 163646 606556 163648
rect 599945 163643 600011 163646
rect 666645 163570 666711 163573
rect 672441 163570 672507 163573
rect 666356 163568 672507 163570
rect 666356 163512 666650 163568
rect 666706 163512 672446 163568
rect 672502 163512 672507 163568
rect 666356 163510 672507 163512
rect 666645 163507 666711 163510
rect 672441 163507 672507 163510
rect 581821 163162 581887 163165
rect 576380 163160 581887 163162
rect 576380 163104 581826 163160
rect 581882 163104 581887 163160
rect 576380 163102 581887 163104
rect 581821 163099 581887 163102
rect 599853 162618 599919 162621
rect 599853 162616 606556 162618
rect 599853 162560 599858 162616
rect 599914 162560 606556 162616
rect 599853 162558 606556 162560
rect 599853 162555 599919 162558
rect 600037 161666 600103 161669
rect 600037 161664 606556 161666
rect 600037 161608 600042 161664
rect 600098 161608 606556 161664
rect 600037 161606 606556 161608
rect 600037 161603 600103 161606
rect 579889 161530 579955 161533
rect 576380 161528 579955 161530
rect 576380 161472 579894 161528
rect 579950 161472 579955 161528
rect 576380 161470 579955 161472
rect 579889 161467 579955 161470
rect 599945 160578 600011 160581
rect 599945 160576 606556 160578
rect 599945 160520 599950 160576
rect 600006 160520 606556 160576
rect 599945 160518 606556 160520
rect 599945 160515 600011 160518
rect 666645 160170 666711 160173
rect 666356 160168 666711 160170
rect 666356 160112 666650 160168
rect 666706 160112 666711 160168
rect 666356 160110 666711 160112
rect 666645 160107 666711 160110
rect 582189 160034 582255 160037
rect 576380 160032 582255 160034
rect 576380 159976 582194 160032
rect 582250 159976 582255 160032
rect 576380 159974 582255 159976
rect 582189 159971 582255 159974
rect 598933 159626 598999 159629
rect 598933 159624 606556 159626
rect 598933 159568 598938 159624
rect 598994 159568 606556 159624
rect 598933 159566 606556 159568
rect 598933 159563 598999 159566
rect 579705 158538 579771 158541
rect 576380 158536 579771 158538
rect 576380 158480 579710 158536
rect 579766 158480 579771 158536
rect 576380 158478 579771 158480
rect 579705 158475 579771 158478
rect 599853 158538 599919 158541
rect 599853 158536 606556 158538
rect 599853 158480 599858 158536
rect 599914 158480 606556 158536
rect 599853 158478 606556 158480
rect 599853 158475 599919 158478
rect 666645 158402 666711 158405
rect 672533 158402 672599 158405
rect 666356 158400 672599 158402
rect 666356 158344 666650 158400
rect 666706 158344 672538 158400
rect 672594 158344 672599 158400
rect 666356 158342 672599 158344
rect 666645 158339 666711 158342
rect 672533 158339 672599 158342
rect 599945 157586 600011 157589
rect 599945 157584 606556 157586
rect 599945 157528 599950 157584
rect 600006 157528 606556 157584
rect 599945 157526 606556 157528
rect 599945 157523 600011 157526
rect 580165 157042 580231 157045
rect 576380 157040 580231 157042
rect 576380 156984 580170 157040
rect 580226 156984 580231 157040
rect 576380 156982 580231 156984
rect 580165 156979 580231 156982
rect 599853 156498 599919 156501
rect 675753 156500 675819 156501
rect 599853 156496 606556 156498
rect 599853 156440 599858 156496
rect 599914 156440 606556 156496
rect 599853 156438 606556 156440
rect 599853 156435 599919 156438
rect 675702 156436 675708 156500
rect 675772 156498 675819 156500
rect 675772 156496 675864 156498
rect 675814 156440 675864 156496
rect 675772 156438 675864 156440
rect 675772 156436 675819 156438
rect 675753 156435 675819 156436
rect 582097 155546 582163 155549
rect 576380 155544 582163 155546
rect 576380 155488 582102 155544
rect 582158 155488 582163 155544
rect 576380 155486 582163 155488
rect 582097 155483 582163 155486
rect 599945 155546 600011 155549
rect 599945 155544 606556 155546
rect 599945 155488 599950 155544
rect 600006 155488 606556 155544
rect 599945 155486 606556 155488
rect 599945 155483 600011 155486
rect 666645 155002 666711 155005
rect 666356 155000 666711 155002
rect 666356 154944 666650 155000
rect 666706 154944 666711 155000
rect 666356 154942 666711 154944
rect 666645 154939 666711 154942
rect 600037 154458 600103 154461
rect 600037 154456 606556 154458
rect 600037 154400 600042 154456
rect 600098 154400 606556 154456
rect 600037 154398 606556 154400
rect 600037 154395 600103 154398
rect 581269 154050 581335 154053
rect 576380 154048 581335 154050
rect 576380 153992 581274 154048
rect 581330 153992 581335 154048
rect 576380 153990 581335 153992
rect 581269 153987 581335 153990
rect 599853 153506 599919 153509
rect 599853 153504 606556 153506
rect 599853 153448 599858 153504
rect 599914 153448 606556 153504
rect 599853 153446 606556 153448
rect 599853 153443 599919 153446
rect 666645 153370 666711 153373
rect 672625 153370 672691 153373
rect 666356 153368 672691 153370
rect 666356 153312 666650 153368
rect 666706 153312 672630 153368
rect 672686 153312 672691 153368
rect 666356 153310 672691 153312
rect 666645 153307 666711 153310
rect 672625 153307 672691 153310
rect 580349 152418 580415 152421
rect 576380 152416 580415 152418
rect 576380 152360 580354 152416
rect 580410 152360 580415 152416
rect 576380 152358 580415 152360
rect 580349 152355 580415 152358
rect 599945 152418 600011 152421
rect 599945 152416 606556 152418
rect 599945 152360 599950 152416
rect 600006 152360 606556 152416
rect 599945 152358 606556 152360
rect 599945 152355 600011 152358
rect 598933 151466 598999 151469
rect 598933 151464 606556 151466
rect 598933 151408 598938 151464
rect 598994 151408 606556 151464
rect 598933 151406 606556 151408
rect 598933 151403 598999 151406
rect 581913 150922 581979 150925
rect 576380 150920 581979 150922
rect 576380 150864 581918 150920
rect 581974 150864 581979 150920
rect 576380 150862 581979 150864
rect 581913 150859 581979 150862
rect 599853 150378 599919 150381
rect 599853 150376 606556 150378
rect 599853 150320 599858 150376
rect 599914 150320 606556 150376
rect 599853 150318 606556 150320
rect 599853 150315 599919 150318
rect 666645 149970 666711 149973
rect 666356 149968 666711 149970
rect 666356 149912 666650 149968
rect 666706 149912 666711 149968
rect 666356 149910 666711 149912
rect 666645 149907 666711 149910
rect 581453 149426 581519 149429
rect 576380 149424 581519 149426
rect 576380 149368 581458 149424
rect 581514 149368 581519 149424
rect 576380 149366 581519 149368
rect 581453 149363 581519 149366
rect 599945 149426 600011 149429
rect 599945 149424 606556 149426
rect 599945 149368 599950 149424
rect 600006 149368 606556 149424
rect 599945 149366 606556 149368
rect 599945 149363 600011 149366
rect 675753 148474 675819 148477
rect 675886 148474 675892 148476
rect 675753 148472 675892 148474
rect 675753 148416 675758 148472
rect 675814 148416 675892 148472
rect 675753 148414 675892 148416
rect 675753 148411 675819 148414
rect 675886 148412 675892 148414
rect 675956 148412 675962 148476
rect 599853 148338 599919 148341
rect 599853 148336 606556 148338
rect 599853 148280 599858 148336
rect 599914 148280 606556 148336
rect 599853 148278 606556 148280
rect 599853 148275 599919 148278
rect 666645 148202 666711 148205
rect 672717 148202 672783 148205
rect 666356 148200 672783 148202
rect 666356 148144 666650 148200
rect 666706 148144 672722 148200
rect 672778 148144 672783 148200
rect 666356 148142 672783 148144
rect 666645 148139 666711 148142
rect 672717 148139 672783 148142
rect 580993 147930 581059 147933
rect 576380 147928 581059 147930
rect 576380 147872 580998 147928
rect 581054 147872 581059 147928
rect 576380 147870 581059 147872
rect 580993 147867 581059 147870
rect 599945 147386 600011 147389
rect 599945 147384 606556 147386
rect 599945 147328 599950 147384
rect 600006 147328 606556 147384
rect 599945 147326 606556 147328
rect 599945 147323 600011 147326
rect 580533 146434 580599 146437
rect 576380 146432 580599 146434
rect 576380 146376 580538 146432
rect 580594 146376 580599 146432
rect 576380 146374 580599 146376
rect 580533 146371 580599 146374
rect 600037 146298 600103 146301
rect 675753 146298 675819 146301
rect 676070 146298 676076 146300
rect 600037 146296 606556 146298
rect 600037 146240 600042 146296
rect 600098 146240 606556 146296
rect 600037 146238 606556 146240
rect 675753 146296 676076 146298
rect 675753 146240 675758 146296
rect 675814 146240 676076 146296
rect 675753 146238 676076 146240
rect 600037 146235 600103 146238
rect 675753 146235 675819 146238
rect 676070 146236 676076 146238
rect 676140 146236 676146 146300
rect 599853 145346 599919 145349
rect 599853 145344 606556 145346
rect 599853 145288 599858 145344
rect 599914 145288 606556 145344
rect 599853 145286 606556 145288
rect 599853 145283 599919 145286
rect 581177 144938 581243 144941
rect 666645 144938 666711 144941
rect 576380 144936 581243 144938
rect 576380 144880 581182 144936
rect 581238 144880 581243 144936
rect 576380 144878 581243 144880
rect 666356 144936 666711 144938
rect 666356 144880 666650 144936
rect 666706 144880 666711 144936
rect 666356 144878 666711 144880
rect 581177 144875 581243 144878
rect 666645 144875 666711 144878
rect 599945 144258 600011 144261
rect 599945 144256 606556 144258
rect 599945 144200 599950 144256
rect 600006 144200 606556 144256
rect 599945 144198 606556 144200
rect 599945 144195 600011 144198
rect 581085 143306 581151 143309
rect 576380 143304 581151 143306
rect 576380 143248 581090 143304
rect 581146 143248 581151 143304
rect 576380 143246 581151 143248
rect 581085 143243 581151 143246
rect 599853 143306 599919 143309
rect 599853 143304 606556 143306
rect 599853 143248 599858 143304
rect 599914 143248 606556 143304
rect 599853 143246 606556 143248
rect 599853 143243 599919 143246
rect 666645 143170 666711 143173
rect 672901 143170 672967 143173
rect 666356 143168 672967 143170
rect 666356 143112 666650 143168
rect 666706 143112 672906 143168
rect 672962 143112 672967 143168
rect 666356 143110 672967 143112
rect 666645 143107 666711 143110
rect 672901 143107 672967 143110
rect 599945 142218 600011 142221
rect 599945 142216 606556 142218
rect 599945 142160 599950 142216
rect 600006 142160 606556 142216
rect 599945 142158 606556 142160
rect 599945 142155 600011 142158
rect 580809 141810 580875 141813
rect 576380 141808 580875 141810
rect 576380 141752 580814 141808
rect 580870 141752 580875 141808
rect 576380 141750 580875 141752
rect 580809 141747 580875 141750
rect 599301 141266 599367 141269
rect 599301 141264 606556 141266
rect 599301 141208 599306 141264
rect 599362 141208 606556 141264
rect 599301 141206 606556 141208
rect 599301 141203 599367 141206
rect 580901 140314 580967 140317
rect 576380 140312 580967 140314
rect 576380 140256 580906 140312
rect 580962 140256 580967 140312
rect 576380 140254 580967 140256
rect 580901 140251 580967 140254
rect 599853 140178 599919 140181
rect 599853 140176 606556 140178
rect 599853 140120 599858 140176
rect 599914 140120 606556 140176
rect 599853 140118 606556 140120
rect 599853 140115 599919 140118
rect 666645 139770 666711 139773
rect 666356 139768 666711 139770
rect 666356 139712 666650 139768
rect 666706 139712 666711 139768
rect 666356 139710 666711 139712
rect 666645 139707 666711 139710
rect 599761 139226 599827 139229
rect 599761 139224 606556 139226
rect 599761 139168 599766 139224
rect 599822 139168 606556 139224
rect 599761 139166 606556 139168
rect 599761 139163 599827 139166
rect 580717 138818 580783 138821
rect 576380 138816 580783 138818
rect 576380 138760 580722 138816
rect 580778 138760 580783 138816
rect 576380 138758 580783 138760
rect 580717 138755 580783 138758
rect 599945 138138 600011 138141
rect 670693 138138 670759 138141
rect 672993 138138 673059 138141
rect 599945 138136 606556 138138
rect 599945 138080 599950 138136
rect 600006 138080 606556 138136
rect 599945 138078 606556 138080
rect 666356 138136 673059 138138
rect 666356 138080 670698 138136
rect 670754 138080 672998 138136
rect 673054 138080 673059 138136
rect 666356 138078 673059 138080
rect 599945 138075 600011 138078
rect 670693 138075 670759 138078
rect 672993 138075 673059 138078
rect 582005 137322 582071 137325
rect 576380 137320 582071 137322
rect 576380 137264 582010 137320
rect 582066 137264 582071 137320
rect 576380 137262 582071 137264
rect 582005 137259 582071 137262
rect 599853 137186 599919 137189
rect 599853 137184 606556 137186
rect 599853 137128 599858 137184
rect 599914 137128 606556 137184
rect 599853 137126 606556 137128
rect 599853 137123 599919 137126
rect 599945 136098 600011 136101
rect 599945 136096 606556 136098
rect 599945 136040 599950 136096
rect 600006 136040 606556 136096
rect 599945 136038 606556 136040
rect 599945 136035 600011 136038
rect 582189 135826 582255 135829
rect 576380 135824 582255 135826
rect 576380 135768 582194 135824
rect 582250 135768 582255 135824
rect 576380 135766 582255 135768
rect 582189 135763 582255 135766
rect 600037 135146 600103 135149
rect 600037 135144 606556 135146
rect 600037 135088 600042 135144
rect 600098 135088 606556 135144
rect 600037 135086 606556 135088
rect 600037 135083 600103 135086
rect 670693 134738 670759 134741
rect 666356 134736 670759 134738
rect 666356 134680 670698 134736
rect 670754 134680 670759 134736
rect 666356 134678 670759 134680
rect 670693 134675 670759 134678
rect 582097 134194 582163 134197
rect 576380 134192 582163 134194
rect 576380 134136 582102 134192
rect 582158 134136 582163 134192
rect 576380 134134 582163 134136
rect 582097 134131 582163 134134
rect 703813 134194 703879 134197
rect 709057 134194 709123 134197
rect 703813 134134 709123 134194
rect 703813 134131 703879 134134
rect 709057 134131 709123 134134
rect 599853 134058 599919 134061
rect 599853 134056 606556 134058
rect 599853 134000 599858 134056
rect 599914 134000 606556 134056
rect 599853 133998 606556 134000
rect 599853 133995 599919 133998
rect 599945 133106 600011 133109
rect 676121 133106 676187 133109
rect 676262 133106 676322 133348
rect 599945 133104 606556 133106
rect 599945 133048 599950 133104
rect 600006 133048 606556 133104
rect 599945 133046 606556 133048
rect 676121 133104 676322 133106
rect 676121 133048 676126 133104
rect 676182 133048 676322 133104
rect 676121 133046 676322 133048
rect 599945 133043 600011 133046
rect 676121 133043 676187 133046
rect 666645 132970 666711 132973
rect 673085 132970 673151 132973
rect 666356 132968 673151 132970
rect 666356 132912 666650 132968
rect 666706 132912 673090 132968
rect 673146 132912 673151 132968
rect 666356 132910 673151 132912
rect 666645 132907 666711 132910
rect 673085 132907 673151 132910
rect 676029 132970 676095 132973
rect 676029 132968 676292 132970
rect 676029 132912 676034 132968
rect 676090 132912 676292 132968
rect 676029 132910 676292 132912
rect 676029 132907 676095 132910
rect 582281 132698 582347 132701
rect 576380 132696 582347 132698
rect 576380 132640 582286 132696
rect 582342 132640 582347 132696
rect 576380 132638 582347 132640
rect 582281 132635 582347 132638
rect 676213 132698 676279 132701
rect 676213 132696 676322 132698
rect 676213 132640 676218 132696
rect 676274 132640 676322 132696
rect 676213 132635 676322 132640
rect 676262 132532 676322 132635
rect 676213 132290 676279 132293
rect 676213 132288 676322 132290
rect 676213 132232 676218 132288
rect 676274 132232 676322 132288
rect 676213 132227 676322 132232
rect 676262 132124 676322 132227
rect 599853 132018 599919 132021
rect 599853 132016 606556 132018
rect 599853 131960 599858 132016
rect 599914 131960 606556 132016
rect 599853 131958 606556 131960
rect 599853 131955 599919 131958
rect 676029 131746 676095 131749
rect 676029 131744 676292 131746
rect 676029 131688 676034 131744
rect 676090 131688 676292 131744
rect 676029 131686 676292 131688
rect 676029 131683 676095 131686
rect 676213 131474 676279 131477
rect 676213 131472 676322 131474
rect 676213 131416 676218 131472
rect 676274 131416 676322 131472
rect 676213 131411 676322 131416
rect 676262 131308 676322 131411
rect 581821 131202 581887 131205
rect 576380 131200 581887 131202
rect 576380 131144 581826 131200
rect 581882 131144 581887 131200
rect 576380 131142 581887 131144
rect 581821 131139 581887 131142
rect 599761 131066 599827 131069
rect 599761 131064 606556 131066
rect 599761 131008 599766 131064
rect 599822 131008 606556 131064
rect 599761 131006 606556 131008
rect 599761 131003 599827 131006
rect 676029 130930 676095 130933
rect 676029 130928 676292 130930
rect 676029 130872 676034 130928
rect 676090 130872 676292 130928
rect 676029 130870 676292 130872
rect 676029 130867 676095 130870
rect 676213 130658 676279 130661
rect 676213 130656 676322 130658
rect 676213 130600 676218 130656
rect 676274 130600 676322 130656
rect 676213 130595 676322 130600
rect 676262 130492 676322 130595
rect 676029 130114 676095 130117
rect 676029 130112 676292 130114
rect 676029 130056 676034 130112
rect 676090 130056 676292 130112
rect 676029 130054 676292 130056
rect 676029 130051 676095 130054
rect 599945 129978 600011 129981
rect 599945 129976 606556 129978
rect 599945 129920 599950 129976
rect 600006 129920 606556 129976
rect 599945 129918 606556 129920
rect 599945 129915 600011 129918
rect 581913 129706 581979 129709
rect 576380 129704 581979 129706
rect 576380 129648 581918 129704
rect 581974 129648 581979 129704
rect 576380 129646 581979 129648
rect 581913 129643 581979 129646
rect 676029 129706 676095 129709
rect 676029 129704 676292 129706
rect 676029 129648 676034 129704
rect 676090 129648 676292 129704
rect 676029 129646 676292 129648
rect 676029 129643 676095 129646
rect 666645 129570 666711 129573
rect 666356 129568 666711 129570
rect 666356 129512 666650 129568
rect 666706 129512 666711 129568
rect 666356 129510 666711 129512
rect 666645 129507 666711 129510
rect 676213 129434 676279 129437
rect 676213 129432 676322 129434
rect 676213 129376 676218 129432
rect 676274 129376 676322 129432
rect 676213 129371 676322 129376
rect 676262 129268 676322 129371
rect 599853 129026 599919 129029
rect 599853 129024 606556 129026
rect 599853 128968 599858 129024
rect 599914 128968 606556 129024
rect 599853 128966 606556 128968
rect 599853 128963 599919 128966
rect 676029 128890 676095 128893
rect 676029 128888 676292 128890
rect 676029 128832 676034 128888
rect 676090 128832 676292 128888
rect 676029 128830 676292 128832
rect 676029 128827 676095 128830
rect 675886 128420 675892 128484
rect 675956 128482 675962 128484
rect 675956 128422 676292 128482
rect 675956 128420 675962 128422
rect 580625 128210 580691 128213
rect 576380 128208 580691 128210
rect 576380 128152 580630 128208
rect 580686 128152 580691 128208
rect 576380 128150 580691 128152
rect 580625 128147 580691 128150
rect 675753 128074 675819 128077
rect 675753 128072 676292 128074
rect 675753 128016 675758 128072
rect 675814 128016 676292 128072
rect 675753 128014 676292 128016
rect 675753 128011 675819 128014
rect 599945 127938 600011 127941
rect 666645 127938 666711 127941
rect 672809 127938 672875 127941
rect 599945 127936 606556 127938
rect 599945 127880 599950 127936
rect 600006 127880 606556 127936
rect 599945 127878 606556 127880
rect 666356 127936 672875 127938
rect 666356 127880 666650 127936
rect 666706 127880 672814 127936
rect 672870 127880 672875 127936
rect 666356 127878 672875 127880
rect 599945 127875 600011 127878
rect 666645 127875 666711 127878
rect 672809 127875 672875 127878
rect 676029 127666 676095 127669
rect 676029 127664 676292 127666
rect 676029 127608 676034 127664
rect 676090 127608 676292 127664
rect 676029 127606 676292 127608
rect 676029 127603 676095 127606
rect 675937 127258 676003 127261
rect 675937 127256 676292 127258
rect 675937 127200 675942 127256
rect 675998 127200 676292 127256
rect 675937 127198 676292 127200
rect 675937 127195 676003 127198
rect 599761 126986 599827 126989
rect 599761 126984 606556 126986
rect 599761 126928 599766 126984
rect 599822 126928 606556 126984
rect 599761 126926 606556 126928
rect 599761 126923 599827 126926
rect 581361 126714 581427 126717
rect 576380 126712 581427 126714
rect 576380 126656 581366 126712
rect 581422 126656 581427 126712
rect 576380 126654 581427 126656
rect 581361 126651 581427 126654
rect 676070 126516 676076 126580
rect 676140 126578 676146 126580
rect 676262 126578 676322 126820
rect 676140 126518 676322 126578
rect 676140 126516 676146 126518
rect 676029 126442 676095 126445
rect 676029 126440 676292 126442
rect 676029 126384 676034 126440
rect 676090 126384 676292 126440
rect 676029 126382 676292 126384
rect 676029 126379 676095 126382
rect 675937 126034 676003 126037
rect 675937 126032 676292 126034
rect 675937 125976 675942 126032
rect 675998 125976 676292 126032
rect 675937 125974 676292 125976
rect 675937 125971 676003 125974
rect 600037 125898 600103 125901
rect 600037 125896 606556 125898
rect 600037 125840 600042 125896
rect 600098 125840 606556 125896
rect 600037 125838 606556 125840
rect 600037 125835 600103 125838
rect 676121 125354 676187 125357
rect 676262 125354 676322 125596
rect 676121 125352 676322 125354
rect 676121 125296 676126 125352
rect 676182 125296 676322 125352
rect 676121 125294 676322 125296
rect 676121 125291 676187 125294
rect 675845 125218 675911 125221
rect 675845 125216 676292 125218
rect 675845 125160 675850 125216
rect 675906 125160 676292 125216
rect 675845 125158 676292 125160
rect 675845 125155 675911 125158
rect 581545 125082 581611 125085
rect 576380 125080 581611 125082
rect 576380 125024 581550 125080
rect 581606 125024 581611 125080
rect 576380 125022 581611 125024
rect 581545 125019 581611 125022
rect 599945 124946 600011 124949
rect 599945 124944 606556 124946
rect 599945 124888 599950 124944
rect 600006 124888 606556 124944
rect 599945 124886 606556 124888
rect 599945 124883 600011 124886
rect 675661 124810 675727 124813
rect 675661 124808 676292 124810
rect 675661 124752 675666 124808
rect 675722 124752 676292 124808
rect 675661 124750 676292 124752
rect 675661 124747 675727 124750
rect 666645 124538 666711 124541
rect 666356 124536 666711 124538
rect 666356 124480 666650 124536
rect 666706 124480 666711 124536
rect 666356 124478 666711 124480
rect 666645 124475 666711 124478
rect 675937 124402 676003 124405
rect 675937 124400 676292 124402
rect 675937 124344 675942 124400
rect 675998 124344 676292 124400
rect 675937 124342 676292 124344
rect 675937 124339 676003 124342
rect 676029 123994 676095 123997
rect 676029 123992 676292 123994
rect 676029 123936 676034 123992
rect 676090 123936 676292 123992
rect 676029 123934 676292 123936
rect 676029 123931 676095 123934
rect 600037 123858 600103 123861
rect 600037 123856 606556 123858
rect 600037 123800 600042 123856
rect 600098 123800 606556 123856
rect 600037 123798 606556 123800
rect 600037 123795 600103 123798
rect 581453 123586 581519 123589
rect 576380 123584 581519 123586
rect 576380 123528 581458 123584
rect 581514 123528 581519 123584
rect 576380 123526 581519 123528
rect 581453 123523 581519 123526
rect 675937 123586 676003 123589
rect 675937 123584 676292 123586
rect 675937 123528 675942 123584
rect 675998 123528 676292 123584
rect 675937 123526 676292 123528
rect 675937 123523 676003 123526
rect 676029 123178 676095 123181
rect 676029 123176 676292 123178
rect 676029 123120 676034 123176
rect 676090 123120 676292 123176
rect 676029 123118 676292 123120
rect 676029 123115 676095 123118
rect 599853 122906 599919 122909
rect 666645 122906 666711 122909
rect 673177 122906 673243 122909
rect 599853 122904 606556 122906
rect 599853 122848 599858 122904
rect 599914 122848 606556 122904
rect 599853 122846 606556 122848
rect 666356 122904 673243 122906
rect 666356 122848 666650 122904
rect 666706 122848 673182 122904
rect 673238 122848 673243 122904
rect 666356 122846 673243 122848
rect 599853 122843 599919 122846
rect 666645 122843 666711 122846
rect 673177 122843 673243 122846
rect 676029 122770 676095 122773
rect 676029 122768 676292 122770
rect 676029 122712 676034 122768
rect 676090 122712 676292 122768
rect 676029 122710 676292 122712
rect 676029 122707 676095 122710
rect 579705 122090 579771 122093
rect 576380 122088 579771 122090
rect 576380 122032 579710 122088
rect 579766 122032 579771 122088
rect 576380 122030 579771 122032
rect 579705 122027 579771 122030
rect 676029 121954 676095 121957
rect 676029 121952 676292 121954
rect 676029 121896 676034 121952
rect 676090 121896 676292 121952
rect 676029 121894 676292 121896
rect 676029 121891 676095 121894
rect 599945 121818 600011 121821
rect 599945 121816 606556 121818
rect 599945 121760 599950 121816
rect 600006 121760 606556 121816
rect 599945 121758 606556 121760
rect 599945 121755 600011 121758
rect 600037 120866 600103 120869
rect 600037 120864 606556 120866
rect 600037 120808 600042 120864
rect 600098 120808 606556 120864
rect 600037 120806 606556 120808
rect 600037 120803 600103 120806
rect 581269 120594 581335 120597
rect 576380 120592 581335 120594
rect 576380 120536 581274 120592
rect 581330 120536 581335 120592
rect 576380 120534 581335 120536
rect 581269 120531 581335 120534
rect 599945 119778 600011 119781
rect 599945 119776 606556 119778
rect 599945 119720 599950 119776
rect 600006 119720 606556 119776
rect 599945 119718 606556 119720
rect 599945 119715 600011 119718
rect 666645 119506 666711 119509
rect 666356 119504 666711 119506
rect 666356 119448 666650 119504
rect 666706 119448 666711 119504
rect 666356 119446 666711 119448
rect 666645 119443 666711 119446
rect 581729 119098 581795 119101
rect 576380 119096 581795 119098
rect 576380 119040 581734 119096
rect 581790 119040 581795 119096
rect 576380 119038 581795 119040
rect 581729 119035 581795 119038
rect 599853 118826 599919 118829
rect 599853 118824 606556 118826
rect 599853 118768 599858 118824
rect 599914 118768 606556 118824
rect 599853 118766 606556 118768
rect 599853 118763 599919 118766
rect 599853 117738 599919 117741
rect 672165 117738 672231 117741
rect 599853 117736 606556 117738
rect 599853 117680 599858 117736
rect 599914 117680 606556 117736
rect 599853 117678 606556 117680
rect 666356 117736 672231 117738
rect 666356 117680 672170 117736
rect 672226 117680 672231 117736
rect 666356 117678 672231 117680
rect 599853 117675 599919 117678
rect 672165 117675 672231 117678
rect 581637 117602 581703 117605
rect 576380 117600 581703 117602
rect 576380 117544 581642 117600
rect 581698 117544 581703 117600
rect 576380 117542 581703 117544
rect 581637 117539 581703 117542
rect 599945 116786 600011 116789
rect 599945 116784 606556 116786
rect 599945 116728 599950 116784
rect 600006 116728 606556 116784
rect 599945 116726 606556 116728
rect 599945 116723 600011 116726
rect 672349 116106 672415 116109
rect 666356 116104 672415 116106
rect 666356 116048 672354 116104
rect 672410 116048 672415 116104
rect 666356 116046 672415 116048
rect 672349 116043 672415 116046
rect 580993 115970 581059 115973
rect 576380 115968 581059 115970
rect 576380 115912 580998 115968
rect 581054 115912 581059 115968
rect 576380 115910 581059 115912
rect 580993 115907 581059 115910
rect 599853 115698 599919 115701
rect 599853 115696 606556 115698
rect 599853 115640 599858 115696
rect 599914 115640 606556 115696
rect 599853 115638 606556 115640
rect 599853 115635 599919 115638
rect 599945 114746 600011 114749
rect 599945 114744 606556 114746
rect 599945 114688 599950 114744
rect 600006 114688 606556 114744
rect 599945 114686 606556 114688
rect 599945 114683 600011 114686
rect 581177 114474 581243 114477
rect 576380 114472 581243 114474
rect 576380 114416 581182 114472
rect 581238 114416 581243 114472
rect 576380 114414 581243 114416
rect 581177 114411 581243 114414
rect 672073 114338 672139 114341
rect 666356 114336 672139 114338
rect 666356 114280 672078 114336
rect 672134 114280 672139 114336
rect 666356 114278 672139 114280
rect 672073 114275 672139 114278
rect 593370 113598 606556 113658
rect 580942 113188 580948 113252
rect 581012 113250 581018 113252
rect 593370 113250 593430 113598
rect 581012 113190 593430 113250
rect 581012 113188 581018 113190
rect 579797 112978 579863 112981
rect 576380 112976 579863 112978
rect 576380 112920 579802 112976
rect 579858 112920 579863 112976
rect 576380 112918 579863 112920
rect 579797 112915 579863 112918
rect 599945 112706 600011 112709
rect 672901 112706 672967 112709
rect 599945 112704 606556 112706
rect 599945 112648 599950 112704
rect 600006 112648 606556 112704
rect 599945 112646 606556 112648
rect 666356 112704 672967 112706
rect 666356 112648 672906 112704
rect 672962 112648 672967 112704
rect 666356 112646 672967 112648
rect 599945 112643 600011 112646
rect 672901 112643 672967 112646
rect 599761 111618 599827 111621
rect 599761 111616 606556 111618
rect 599761 111560 599766 111616
rect 599822 111560 606556 111616
rect 599761 111558 606556 111560
rect 599761 111555 599827 111558
rect 580073 111482 580139 111485
rect 576380 111480 580139 111482
rect 576380 111424 580078 111480
rect 580134 111424 580139 111480
rect 576380 111422 580139 111424
rect 580073 111419 580139 111422
rect 671613 110938 671679 110941
rect 666356 110936 671679 110938
rect 666356 110880 671618 110936
rect 671674 110880 671679 110936
rect 666356 110878 671679 110880
rect 671613 110875 671679 110878
rect 600221 110666 600287 110669
rect 600221 110664 606556 110666
rect 600221 110608 600226 110664
rect 600282 110608 606556 110664
rect 600221 110606 606556 110608
rect 600221 110603 600287 110606
rect 581085 109986 581151 109989
rect 576380 109984 581151 109986
rect 576380 109928 581090 109984
rect 581146 109928 581151 109984
rect 576380 109926 581151 109928
rect 581085 109923 581151 109926
rect 599945 109578 600011 109581
rect 599945 109576 606556 109578
rect 599945 109520 599950 109576
rect 600006 109520 606556 109576
rect 599945 109518 606556 109520
rect 599945 109515 600011 109518
rect 672257 109306 672323 109309
rect 666356 109304 672323 109306
rect 666356 109248 672262 109304
rect 672318 109248 672323 109304
rect 666356 109246 672323 109248
rect 672257 109243 672323 109246
rect 600313 108626 600379 108629
rect 600313 108624 606556 108626
rect 600313 108568 600318 108624
rect 600374 108568 606556 108624
rect 600313 108566 606556 108568
rect 600313 108563 600379 108566
rect 579889 108490 579955 108493
rect 576380 108488 579955 108490
rect 576380 108432 579894 108488
rect 579950 108432 579955 108488
rect 576380 108430 579955 108432
rect 579889 108427 579955 108430
rect 599945 107538 600011 107541
rect 671153 107538 671219 107541
rect 599945 107536 606556 107538
rect 599945 107480 599950 107536
rect 600006 107480 606556 107536
rect 599945 107478 606556 107480
rect 666356 107536 671219 107538
rect 666356 107480 671158 107536
rect 671214 107480 671219 107536
rect 666356 107478 671219 107480
rect 599945 107475 600011 107478
rect 671153 107475 671219 107478
rect 580165 106858 580231 106861
rect 576380 106856 580231 106858
rect 576380 106800 580170 106856
rect 580226 106800 580231 106856
rect 576380 106798 580231 106800
rect 580165 106795 580231 106798
rect 600589 106586 600655 106589
rect 600589 106584 606556 106586
rect 600589 106528 600594 106584
rect 600650 106528 606556 106584
rect 600589 106526 606556 106528
rect 600589 106523 600655 106526
rect 672441 105906 672507 105909
rect 666356 105904 672507 105906
rect 666356 105848 672446 105904
rect 672502 105848 672507 105904
rect 666356 105846 672507 105848
rect 672441 105843 672507 105846
rect 600405 105498 600471 105501
rect 600405 105496 606556 105498
rect 600405 105440 600410 105496
rect 600466 105440 606556 105496
rect 600405 105438 606556 105440
rect 600405 105435 600471 105438
rect 579981 105362 580047 105365
rect 576380 105360 580047 105362
rect 576380 105304 579986 105360
rect 580042 105304 580047 105360
rect 576380 105302 580047 105304
rect 579981 105299 580047 105302
rect 600681 104546 600747 104549
rect 600681 104544 606556 104546
rect 600681 104488 600686 104544
rect 600742 104488 606556 104544
rect 600681 104486 606556 104488
rect 600681 104483 600747 104486
rect 670785 104138 670851 104141
rect 666356 104136 670851 104138
rect 666356 104080 670790 104136
rect 670846 104080 670851 104136
rect 666356 104078 670851 104080
rect 670785 104075 670851 104078
rect 580901 103866 580967 103869
rect 576380 103864 580967 103866
rect 576380 103808 580906 103864
rect 580962 103808 580967 103864
rect 576380 103806 580967 103808
rect 580901 103803 580967 103806
rect 600497 103458 600563 103461
rect 600497 103456 606556 103458
rect 600497 103400 600502 103456
rect 600558 103400 606556 103456
rect 600497 103398 606556 103400
rect 600497 103395 600563 103398
rect 675753 103322 675819 103325
rect 675886 103322 675892 103324
rect 675753 103320 675892 103322
rect 675753 103264 675758 103320
rect 675814 103264 675892 103320
rect 675753 103262 675892 103264
rect 675753 103259 675819 103262
rect 675886 103260 675892 103262
rect 675956 103260 675962 103324
rect 600865 102506 600931 102509
rect 671981 102506 672047 102509
rect 600865 102504 606556 102506
rect 600865 102448 600870 102504
rect 600926 102448 606556 102504
rect 600865 102446 606556 102448
rect 666356 102504 672047 102506
rect 666356 102448 671986 102504
rect 672042 102448 672047 102504
rect 666356 102446 672047 102448
rect 600865 102443 600931 102446
rect 671981 102443 672047 102446
rect 580257 102370 580323 102373
rect 576380 102368 580323 102370
rect 576380 102312 580262 102368
rect 580318 102312 580323 102368
rect 576380 102310 580323 102312
rect 580257 102307 580323 102310
rect 600773 101418 600839 101421
rect 675753 101418 675819 101421
rect 676070 101418 676076 101420
rect 600773 101416 606556 101418
rect 600773 101360 600778 101416
rect 600834 101360 606556 101416
rect 600773 101358 606556 101360
rect 675753 101416 676076 101418
rect 675753 101360 675758 101416
rect 675814 101360 676076 101416
rect 675753 101358 676076 101360
rect 600773 101355 600839 101358
rect 675753 101355 675819 101358
rect 676070 101356 676076 101358
rect 676140 101356 676146 101420
rect 580349 100874 580415 100877
rect 670877 100874 670943 100877
rect 576380 100872 580415 100874
rect 576380 100816 580354 100872
rect 580410 100816 580415 100872
rect 576380 100814 580415 100816
rect 666356 100872 670943 100874
rect 666356 100816 670882 100872
rect 670938 100816 670943 100872
rect 666356 100814 670943 100816
rect 580349 100811 580415 100814
rect 670877 100811 670943 100814
rect 599945 100466 600011 100469
rect 599945 100464 606556 100466
rect 599945 100408 599950 100464
rect 600006 100408 606556 100464
rect 599945 100406 606556 100408
rect 599945 100403 600011 100406
rect 580717 99378 580783 99381
rect 576380 99376 580783 99378
rect 576380 99320 580722 99376
rect 580778 99320 580783 99376
rect 576380 99318 580783 99320
rect 580717 99315 580783 99318
rect 580533 97746 580599 97749
rect 576380 97744 580599 97746
rect 576380 97688 580538 97744
rect 580594 97688 580599 97744
rect 576380 97686 580599 97688
rect 580533 97683 580599 97686
rect 580441 96250 580507 96253
rect 576380 96248 580507 96250
rect 576380 96192 580446 96248
rect 580502 96192 580507 96248
rect 576380 96190 580507 96192
rect 580441 96187 580507 96190
rect 628281 95978 628347 95981
rect 628238 95976 628347 95978
rect 628238 95920 628286 95976
rect 628342 95920 628347 95976
rect 628238 95915 628347 95920
rect 628238 95404 628298 95915
rect 640517 95706 640583 95709
rect 640517 95704 642466 95706
rect 640517 95648 640522 95704
rect 640578 95648 642466 95704
rect 640517 95646 642466 95648
rect 640517 95643 640583 95646
rect 580809 94754 580875 94757
rect 576380 94752 580875 94754
rect 576380 94696 580814 94752
rect 580870 94696 580875 94752
rect 576380 94694 580875 94696
rect 580809 94691 580875 94694
rect 642406 94588 642466 95646
rect 662086 95508 662092 95572
rect 662156 95570 662162 95572
rect 662229 95570 662295 95573
rect 662156 95568 662295 95570
rect 662156 95512 662234 95568
rect 662290 95512 662295 95568
rect 662156 95510 662295 95512
rect 662156 95508 662162 95510
rect 662229 95507 662295 95510
rect 657353 94754 657419 94757
rect 657310 94752 657419 94754
rect 657310 94696 657358 94752
rect 657414 94696 657419 94752
rect 657310 94691 657419 94696
rect 627913 94482 627979 94485
rect 627913 94480 628268 94482
rect 627913 94424 627918 94480
rect 627974 94424 628268 94480
rect 627913 94422 628268 94424
rect 627913 94419 627979 94422
rect 657310 94180 657370 94691
rect 663241 93802 663307 93805
rect 663198 93800 663307 93802
rect 663198 93744 663246 93800
rect 663302 93744 663307 93800
rect 663198 93739 663307 93744
rect 627269 93530 627335 93533
rect 627269 93528 628268 93530
rect 627269 93472 627274 93528
rect 627330 93472 628268 93528
rect 627269 93470 628268 93472
rect 627269 93467 627335 93470
rect 655329 93394 655395 93397
rect 655329 93392 656788 93394
rect 655329 93336 655334 93392
rect 655390 93336 656788 93392
rect 663198 93364 663258 93739
rect 655329 93334 656788 93336
rect 655329 93331 655395 93334
rect 580625 93258 580691 93261
rect 576380 93256 580691 93258
rect 576380 93200 580630 93256
rect 580686 93200 580691 93256
rect 576380 93198 580691 93200
rect 580625 93195 580691 93198
rect 663333 93122 663399 93125
rect 663333 93120 663442 93122
rect 663333 93064 663338 93120
rect 663394 93064 663442 93120
rect 663333 93059 663442 93064
rect 642725 92714 642791 92717
rect 642725 92712 642834 92714
rect 642725 92656 642730 92712
rect 642786 92656 642834 92712
rect 642725 92651 642834 92656
rect 626441 92578 626507 92581
rect 626441 92576 628268 92578
rect 626441 92520 626446 92576
rect 626502 92520 628268 92576
rect 626441 92518 628268 92520
rect 626441 92515 626507 92518
rect 642774 92140 642834 92651
rect 652753 92578 652819 92581
rect 652753 92576 656788 92578
rect 652753 92520 652758 92576
rect 652814 92520 656788 92576
rect 663382 92548 663442 93059
rect 652753 92518 656788 92520
rect 652753 92515 652819 92518
rect 663425 92306 663491 92309
rect 663382 92304 663491 92306
rect 663382 92248 663430 92304
rect 663486 92248 663491 92304
rect 663382 92243 663491 92248
rect 582281 91762 582347 91765
rect 576380 91760 582347 91762
rect 576380 91704 582286 91760
rect 582342 91704 582347 91760
rect 663382 91732 663442 92243
rect 576380 91702 582347 91704
rect 582281 91699 582347 91702
rect 625889 91626 625955 91629
rect 625889 91624 628268 91626
rect 625889 91568 625894 91624
rect 625950 91568 628268 91624
rect 625889 91566 628268 91568
rect 625889 91563 625955 91566
rect 654041 91490 654107 91493
rect 654041 91488 656788 91490
rect 654041 91432 654046 91488
rect 654102 91432 656788 91488
rect 654041 91430 656788 91432
rect 654041 91427 654107 91430
rect 663241 91082 663307 91085
rect 663198 91080 663307 91082
rect 663198 91024 663246 91080
rect 663302 91024 663307 91080
rect 663198 91019 663307 91024
rect 623773 90674 623839 90677
rect 652937 90674 653003 90677
rect 623773 90672 628268 90674
rect 623773 90616 623778 90672
rect 623834 90616 628268 90672
rect 623773 90614 628268 90616
rect 652937 90672 656788 90674
rect 652937 90616 652942 90672
rect 652998 90616 656788 90672
rect 663198 90644 663258 91019
rect 652937 90614 656788 90616
rect 623773 90611 623839 90614
rect 652937 90611 653003 90614
rect 656985 90402 657051 90405
rect 663701 90402 663767 90405
rect 656942 90400 657051 90402
rect 656942 90344 656990 90400
rect 657046 90344 657051 90400
rect 656942 90339 657051 90344
rect 663566 90400 663767 90402
rect 663566 90344 663706 90400
rect 663762 90344 663767 90400
rect 663566 90342 663767 90344
rect 582005 90266 582071 90269
rect 576380 90264 582071 90266
rect 576380 90208 582010 90264
rect 582066 90208 582071 90264
rect 576380 90206 582071 90208
rect 582005 90203 582071 90206
rect 656942 89828 657002 90339
rect 663566 89828 663626 90342
rect 663701 90339 663767 90342
rect 623957 89722 624023 89725
rect 645945 89722 646011 89725
rect 623957 89720 628268 89722
rect 623957 89664 623962 89720
rect 624018 89664 628268 89720
rect 623957 89662 628268 89664
rect 642988 89720 646011 89722
rect 642988 89664 645950 89720
rect 646006 89664 646011 89720
rect 642988 89662 646011 89664
rect 623957 89659 624023 89662
rect 645945 89659 646011 89662
rect 663425 89586 663491 89589
rect 663382 89584 663491 89586
rect 663382 89528 663430 89584
rect 663486 89528 663491 89584
rect 663382 89523 663491 89528
rect 663382 89012 663442 89523
rect 623129 88906 623195 88909
rect 623129 88904 628268 88906
rect 623129 88848 623134 88904
rect 623190 88848 628268 88904
rect 623129 88846 628268 88848
rect 623129 88843 623195 88846
rect 662137 88772 662203 88773
rect 662086 88708 662092 88772
rect 662156 88770 662203 88772
rect 662156 88768 662248 88770
rect 662198 88712 662248 88768
rect 662156 88710 662248 88712
rect 662156 88708 662203 88710
rect 662137 88707 662203 88708
rect 582189 88634 582255 88637
rect 576380 88632 582255 88634
rect 576380 88576 582194 88632
rect 582250 88576 582255 88632
rect 576380 88574 582255 88576
rect 582189 88571 582255 88574
rect 623221 87954 623287 87957
rect 623221 87952 628268 87954
rect 623221 87896 623226 87952
rect 623282 87896 628268 87952
rect 623221 87894 628268 87896
rect 623221 87891 623287 87894
rect 582097 87138 582163 87141
rect 646037 87138 646103 87141
rect 576380 87136 582163 87138
rect 576380 87080 582102 87136
rect 582158 87080 582163 87136
rect 576380 87078 582163 87080
rect 642988 87136 646103 87138
rect 642988 87080 646042 87136
rect 646098 87080 646103 87136
rect 642988 87078 646103 87080
rect 582097 87075 582163 87078
rect 646037 87075 646103 87078
rect 623497 87002 623563 87005
rect 623497 87000 628268 87002
rect 623497 86944 623502 87000
rect 623558 86944 628268 87000
rect 623497 86942 628268 86944
rect 623497 86939 623563 86942
rect 622117 86050 622183 86053
rect 622117 86048 628268 86050
rect 622117 85992 622122 86048
rect 622178 85992 628268 86048
rect 622117 85990 628268 85992
rect 622117 85987 622183 85990
rect 581913 85642 581979 85645
rect 576380 85640 581979 85642
rect 576380 85584 581918 85640
rect 581974 85584 581979 85640
rect 576380 85582 581979 85584
rect 581913 85579 581979 85582
rect 622669 85098 622735 85101
rect 622669 85096 628268 85098
rect 622669 85040 622674 85096
rect 622730 85040 628268 85096
rect 622669 85038 628268 85040
rect 622669 85035 622735 85038
rect 646129 84690 646195 84693
rect 642988 84688 646195 84690
rect 642988 84632 646134 84688
rect 646190 84632 646195 84688
rect 642988 84630 646195 84632
rect 646129 84627 646195 84630
rect 581821 84146 581887 84149
rect 576380 84144 581887 84146
rect 576380 84088 581826 84144
rect 581882 84088 581887 84144
rect 576380 84086 581887 84088
rect 581821 84083 581887 84086
rect 621933 84146 621999 84149
rect 621933 84144 628268 84146
rect 621933 84088 621938 84144
rect 621994 84088 628268 84144
rect 621933 84086 628268 84088
rect 621933 84083 621999 84086
rect 623313 83194 623379 83197
rect 623313 83192 628268 83194
rect 623313 83136 623318 83192
rect 623374 83136 628268 83192
rect 623313 83134 628268 83136
rect 623313 83131 623379 83134
rect 579613 82650 579679 82653
rect 576380 82648 579679 82650
rect 576380 82592 579618 82648
rect 579674 82592 579679 82648
rect 576380 82590 579679 82592
rect 579613 82587 579679 82590
rect 622301 82242 622367 82245
rect 645853 82242 645919 82245
rect 622301 82240 628268 82242
rect 622301 82184 622306 82240
rect 622362 82184 628268 82240
rect 622301 82182 628268 82184
rect 642988 82240 645919 82242
rect 642988 82184 645858 82240
rect 645914 82184 645919 82240
rect 642988 82182 645919 82184
rect 622301 82179 622367 82182
rect 645853 82179 645919 82182
rect 622485 81426 622551 81429
rect 622485 81424 628268 81426
rect 622485 81368 622490 81424
rect 622546 81368 628268 81424
rect 622485 81366 628268 81368
rect 622485 81363 622551 81366
rect 581545 81154 581611 81157
rect 576380 81152 581611 81154
rect 576380 81096 581550 81152
rect 581606 81096 581611 81152
rect 576380 81094 581611 81096
rect 581545 81091 581611 81094
rect 581729 79522 581795 79525
rect 576380 79520 581795 79522
rect 576380 79464 581734 79520
rect 581790 79464 581795 79520
rect 576380 79462 581795 79464
rect 581729 79459 581795 79462
rect 581269 78026 581335 78029
rect 576380 78024 581335 78026
rect 576380 77968 581274 78024
rect 581330 77968 581335 78024
rect 576380 77966 581335 77968
rect 581269 77963 581335 77966
rect 581453 76530 581519 76533
rect 576380 76528 581519 76530
rect 576380 76472 581458 76528
rect 581514 76472 581519 76528
rect 576380 76470 581519 76472
rect 581453 76467 581519 76470
rect 581637 75034 581703 75037
rect 576380 75032 581703 75034
rect 576380 74976 581642 75032
rect 581698 74976 581703 75032
rect 576380 74974 581703 74976
rect 581637 74971 581703 74974
rect 580942 73538 580948 73540
rect 576380 73478 580948 73538
rect 580942 73476 580948 73478
rect 581012 73476 581018 73540
rect 581361 72042 581427 72045
rect 576380 72040 581427 72042
rect 576380 71984 581366 72040
rect 581422 71984 581427 72040
rect 576380 71982 581427 71984
rect 581361 71979 581427 71982
rect 580993 70410 581059 70413
rect 576380 70408 581059 70410
rect 576380 70352 580998 70408
rect 581054 70352 581059 70408
rect 576380 70350 581059 70352
rect 580993 70347 581059 70350
rect 582281 68914 582347 68917
rect 576380 68912 582347 68914
rect 576380 68856 582286 68912
rect 582342 68856 582347 68912
rect 576380 68854 582347 68856
rect 582281 68851 582347 68854
rect 581177 67418 581243 67421
rect 576380 67416 581243 67418
rect 576380 67360 581182 67416
rect 581238 67360 581243 67416
rect 576380 67358 581243 67360
rect 581177 67355 581243 67358
rect 580533 65922 580599 65925
rect 576380 65920 580599 65922
rect 576380 65864 580538 65920
rect 580594 65864 580599 65920
rect 576380 65862 580599 65864
rect 580533 65859 580599 65862
rect 581085 64426 581151 64429
rect 576380 64424 581151 64426
rect 576380 64368 581090 64424
rect 581146 64368 581151 64424
rect 576380 64366 581151 64368
rect 581085 64363 581151 64366
rect 582005 62930 582071 62933
rect 576380 62928 582071 62930
rect 576380 62872 582010 62928
rect 582066 62872 582071 62928
rect 576380 62870 582071 62872
rect 582005 62867 582071 62870
rect 582189 61298 582255 61301
rect 576380 61296 582255 61298
rect 576380 61240 582194 61296
rect 582250 61240 582255 61296
rect 576380 61238 582255 61240
rect 582189 61235 582255 61238
rect 579613 59802 579679 59805
rect 576380 59800 579679 59802
rect 576380 59744 579618 59800
rect 579674 59744 579679 59800
rect 576380 59742 579679 59744
rect 579613 59739 579679 59742
rect 579613 58306 579679 58309
rect 576380 58304 579679 58306
rect 576380 58248 579618 58304
rect 579674 58248 579679 58304
rect 576380 58246 579679 58248
rect 579613 58243 579679 58246
rect 581913 56810 581979 56813
rect 576380 56808 581979 56810
rect 576380 56752 581918 56808
rect 581974 56752 581979 56808
rect 576380 56750 581979 56752
rect 581913 56747 581979 56750
rect 582097 55314 582163 55317
rect 576380 55312 582163 55314
rect 576380 55256 582102 55312
rect 582158 55256 582163 55312
rect 576380 55254 582163 55256
rect 582097 55251 582163 55254
rect 580901 53818 580967 53821
rect 576380 53816 580967 53818
rect 576380 53760 580906 53816
rect 580962 53760 580967 53816
rect 576380 53758 580967 53760
rect 580901 53755 580967 53758
rect 666553 48514 666619 48517
rect 662094 48512 666619 48514
rect 661480 48456 666558 48512
rect 666614 48456 666619 48512
rect 661480 48454 666619 48456
rect 661480 48452 662154 48454
rect 666553 48451 666619 48454
rect 281441 48242 281507 48245
rect 520406 48242 520412 48244
rect 281441 48240 520412 48242
rect 281441 48184 281446 48240
rect 281502 48184 520412 48240
rect 281441 48182 520412 48184
rect 281441 48179 281507 48182
rect 520406 48180 520412 48182
rect 520476 48180 520482 48244
rect 661174 47565 661234 47761
rect 661125 47560 661234 47565
rect 661125 47504 661130 47560
rect 661186 47504 661234 47560
rect 661125 47502 661234 47504
rect 661125 47499 661191 47502
rect 665173 47426 665239 47429
rect 661388 47424 665239 47426
rect 661388 47368 665178 47424
rect 665234 47368 665239 47424
rect 661388 47366 665239 47368
rect 665173 47363 665239 47366
rect 661125 46242 661191 46245
rect 620186 46240 661191 46242
rect 620186 46184 661130 46240
rect 661186 46184 661191 46240
rect 620186 46182 661191 46184
rect 236372 46102 256804 46162
rect 187601 41850 187667 41853
rect 194409 41850 194475 41853
rect 187601 41848 187710 41850
rect 187601 41792 187606 41848
rect 187662 41792 187710 41848
rect 187601 41787 187710 41792
rect 194409 41848 207030 41850
rect 194409 41792 194414 41848
rect 194470 41792 207030 41848
rect 194409 41790 207030 41792
rect 194409 41787 194475 41790
rect 187650 41306 187710 41787
rect 206970 41442 207030 41790
rect 236372 41442 236432 46102
rect 206970 41382 236432 41442
rect 256744 41442 256804 46102
rect 518801 44298 518867 44301
rect 518801 44296 526178 44298
rect 518801 44240 518806 44296
rect 518862 44240 526178 44296
rect 518801 44238 526178 44240
rect 518801 44235 518867 44238
rect 526118 44165 526178 44238
rect 526118 44160 526227 44165
rect 526118 44104 526166 44160
rect 526222 44104 526227 44160
rect 526118 44102 526227 44104
rect 526161 44099 526227 44102
rect 520457 42124 520523 42125
rect 520406 42060 520412 42124
rect 520476 42122 520523 42124
rect 520476 42120 520568 42122
rect 520518 42064 520568 42120
rect 520476 42062 520568 42064
rect 520476 42060 520523 42062
rect 520457 42059 520523 42060
rect 470047 41986 470113 41989
rect 571333 41986 571399 41989
rect 470047 41984 571399 41986
rect 470047 41928 470052 41984
rect 470108 41928 571338 41984
rect 571394 41928 571399 41984
rect 470047 41926 571399 41928
rect 470047 41923 470113 41926
rect 571333 41923 571399 41926
rect 307293 41850 307359 41853
rect 362033 41850 362099 41853
rect 415485 41850 415551 41853
rect 552013 41850 552079 41853
rect 307293 41848 322950 41850
rect 307293 41792 307298 41848
rect 307354 41792 322950 41848
rect 307293 41790 322950 41792
rect 307293 41787 307359 41790
rect 322890 41578 322950 41790
rect 362033 41848 380910 41850
rect 362033 41792 362038 41848
rect 362094 41792 380910 41848
rect 362033 41790 380910 41792
rect 362033 41787 362099 41790
rect 380850 41714 380910 41790
rect 415485 41848 552079 41850
rect 415485 41792 415490 41848
rect 415546 41792 552018 41848
rect 552074 41792 552079 41848
rect 415485 41790 552079 41792
rect 415485 41787 415551 41790
rect 552013 41787 552079 41790
rect 563605 41714 563671 41717
rect 380850 41712 563671 41714
rect 380850 41656 563610 41712
rect 563666 41656 563671 41712
rect 380850 41654 563671 41656
rect 563605 41651 563671 41654
rect 587985 41578 588051 41581
rect 322890 41576 588051 41578
rect 322890 41520 587990 41576
rect 588046 41520 588051 41576
rect 322890 41518 588051 41520
rect 587985 41515 588051 41518
rect 620186 41442 620246 46182
rect 661125 46179 661191 46182
rect 256744 41382 620246 41442
rect 209773 41306 209839 41309
rect 212441 41306 212507 41309
rect 187650 41304 212507 41306
rect 187650 41248 209778 41304
rect 209834 41248 212446 41304
rect 212502 41248 212507 41304
rect 187650 41246 212507 41248
rect 209773 41243 209839 41246
rect 212441 41243 212507 41246
rect 530209 41306 530275 41309
rect 542997 41306 543063 41309
rect 530209 41304 543063 41306
rect 530209 41248 530214 41304
rect 530270 41248 543002 41304
rect 543058 41248 543063 41304
rect 530209 41246 543063 41248
rect 530209 41243 530275 41246
rect 542997 41243 543063 41246
rect 230933 16690 230999 16693
rect 225676 16688 230999 16690
rect 225676 16632 230938 16688
rect 230994 16632 230999 16688
rect 225676 16630 230999 16632
rect 230933 16627 230999 16630
rect 230841 15194 230907 15197
rect 225676 15192 230907 15194
rect 225676 15136 230846 15192
rect 230902 15136 230907 15192
rect 225676 15134 230907 15136
rect 230841 15131 230907 15134
rect 230749 13698 230815 13701
rect 225676 13696 230815 13698
rect 225676 13640 230754 13696
rect 230810 13640 230815 13696
rect 225676 13638 230815 13640
rect 230749 13635 230815 13638
rect 230565 12202 230631 12205
rect 225676 12200 230631 12202
rect 225676 12144 230570 12200
rect 230626 12144 230631 12200
rect 225676 12142 230631 12144
rect 230565 12139 230631 12142
rect 230657 10706 230723 10709
rect 225676 10704 230723 10706
rect 225676 10648 230662 10704
rect 230718 10648 230723 10704
rect 225676 10646 230723 10648
rect 230657 10643 230723 10646
rect 230473 9210 230539 9213
rect 225676 9208 230539 9210
rect 225676 9152 230478 9208
rect 230534 9152 230539 9208
rect 225676 9150 230539 9152
rect 230473 9147 230539 9150
rect 230381 7714 230447 7717
rect 225676 7712 230447 7714
rect 225676 7656 230386 7712
rect 230442 7656 230447 7712
rect 225676 7654 230447 7656
rect 230381 7651 230447 7654
rect 229369 6218 229435 6221
rect 225676 6216 229435 6218
rect 225676 6160 229374 6216
rect 229430 6160 229435 6216
rect 225676 6158 229435 6160
rect 229369 6155 229435 6158
<< via3 >>
rect 187740 997188 187804 997252
rect 187740 995692 187804 995756
rect 638540 995208 638604 995212
rect 638540 995152 638544 995208
rect 638544 995152 638600 995208
rect 638600 995152 638604 995208
rect 638540 995148 638604 995152
rect 638540 990524 638604 990588
rect 677172 985900 677236 985964
rect 676988 985764 677052 985828
rect 43668 985628 43732 985692
rect 44036 985492 44100 985556
rect 43484 985356 43548 985420
rect 43852 983044 43916 983108
rect 43300 982908 43364 982972
rect 41460 968764 41524 968828
rect 41644 965092 41708 965156
rect 41828 963384 41892 963388
rect 41828 963328 41842 963384
rect 41842 963328 41892 963384
rect 41828 963324 41892 963328
rect 41828 949452 41892 949516
rect 673868 938300 673932 938364
rect 676812 937212 676876 937276
rect 674972 937076 675036 937140
rect 41828 936940 41892 937004
rect 674788 936260 674852 936324
rect 42012 935308 42076 935372
rect 43300 927148 43364 927212
rect 43484 921980 43548 922044
rect 676076 877236 676140 877300
rect 675708 876616 675772 876620
rect 675708 876560 675722 876616
rect 675722 876560 675772 876616
rect 675708 876556 675772 876560
rect 675524 875936 675588 875940
rect 675524 875880 675538 875936
rect 675538 875880 675588 875936
rect 675524 875876 675588 875880
rect 675340 874032 675404 874036
rect 675340 873976 675390 874032
rect 675390 873976 675404 874032
rect 675340 873972 675404 873976
rect 675892 872204 675956 872268
rect 41828 814192 41892 814196
rect 41828 814136 41878 814192
rect 41878 814136 41892 814192
rect 41828 814132 41892 814136
rect 676260 797676 676324 797740
rect 676444 791964 676508 792028
rect 674972 787748 675036 787812
rect 674604 787204 674668 787268
rect 674420 786796 674484 786860
rect 675156 784076 675220 784140
rect 674788 783804 674852 783868
rect 674236 777412 674300 777476
rect 674236 773332 674300 773396
rect 39988 773060 40052 773124
rect 676812 772652 676876 772716
rect 39988 771428 40052 771492
rect 41460 771020 41524 771084
rect 673868 760276 673932 760340
rect 43300 757692 43364 757756
rect 41828 757072 41892 757076
rect 41828 757016 41842 757072
rect 41842 757016 41892 757072
rect 41828 757012 41892 757016
rect 42196 757012 42260 757076
rect 675524 757012 675588 757076
rect 676076 756332 676140 756396
rect 675340 755788 675404 755852
rect 42196 755244 42260 755308
rect 675708 754564 675772 754628
rect 41828 754080 41892 754084
rect 41828 754024 41878 754080
rect 41878 754024 41892 754080
rect 41828 754020 41892 754024
rect 43300 752932 43364 752996
rect 675892 752524 675956 752588
rect 676444 752252 676508 752316
rect 676260 751844 676324 751908
rect 676628 744092 676692 744156
rect 676260 743956 676324 744020
rect 675892 742868 675956 742932
rect 676076 742460 676140 742524
rect 674052 741644 674116 741708
rect 673868 739740 673932 739804
rect 673684 739060 673748 739124
rect 675708 738576 675772 738580
rect 675708 738520 675722 738576
rect 675722 738520 675772 738576
rect 675708 738516 675772 738520
rect 676444 737972 676508 738036
rect 39988 731036 40052 731100
rect 674420 711996 674484 712060
rect 676260 711886 676324 711890
rect 676260 711830 676310 711886
rect 676310 711830 676324 711886
rect 676260 711826 676324 711830
rect 676996 711886 677060 711890
rect 676996 711830 677010 711886
rect 677010 711830 677060 711886
rect 676996 711826 677060 711830
rect 674972 711180 675036 711244
rect 674604 709548 674668 709612
rect 675156 709140 675220 709204
rect 674788 708732 674852 708796
rect 676812 699756 676876 699820
rect 676260 699620 676324 699684
rect 676996 699484 677060 699548
rect 675524 698184 675588 698188
rect 675524 698128 675538 698184
rect 675538 698128 675588 698184
rect 675524 698124 675588 698128
rect 675340 697232 675404 697236
rect 675340 697176 675390 697232
rect 675390 697176 675404 697232
rect 675340 697172 675404 697176
rect 674236 696628 674300 696692
rect 674420 694996 674484 695060
rect 674604 694180 674668 694244
rect 673500 693636 673564 693700
rect 677180 692956 677244 693020
rect 676628 690100 676692 690164
rect 41276 686700 41340 686764
rect 44036 685204 44100 685268
rect 39988 684252 40052 684316
rect 41276 684252 41340 684316
rect 677364 666980 677428 667044
rect 674052 666844 674116 666908
rect 675892 666028 675956 666092
rect 673868 665620 673932 665684
rect 676076 664532 676140 664596
rect 673684 663988 673748 664052
rect 675708 663580 675772 663644
rect 676260 662900 676324 662964
rect 676444 662492 676508 662556
rect 676996 662084 677060 662148
rect 676812 661676 676876 661740
rect 675156 652564 675220 652628
rect 674972 652156 675036 652220
rect 674788 651612 674852 651676
rect 675892 649164 675956 649228
rect 675708 648680 675772 648684
rect 675708 648624 675722 648680
rect 675722 648624 675772 648680
rect 675708 648620 675772 648624
rect 39988 643452 40052 643516
rect 43668 643452 43732 643516
rect 673684 623052 673748 623116
rect 677364 622780 677428 622844
rect 676260 622372 676324 622436
rect 674236 621828 674300 621892
rect 673684 621556 673748 621620
rect 675524 621012 675588 621076
rect 674420 620604 674484 620668
rect 676076 619516 676140 619580
rect 675340 619380 675404 619444
rect 674604 618972 674668 619036
rect 673500 618564 673564 618628
rect 677180 617476 677244 617540
rect 676628 617068 676692 617132
rect 676444 607684 676508 607748
rect 675524 607608 675588 607612
rect 675524 607552 675538 607608
rect 675538 607552 675588 607608
rect 675524 607548 675588 607552
rect 676628 607412 676692 607476
rect 676076 607276 676140 607340
rect 674420 606460 674484 606524
rect 674236 604692 674300 604756
rect 675340 604344 675404 604348
rect 675340 604288 675390 604344
rect 675390 604288 675404 604344
rect 675340 604284 675404 604288
rect 674604 603468 674668 603532
rect 676260 602924 676324 602988
rect 40172 598572 40236 598636
rect 43852 598028 43916 598092
rect 40172 596124 40236 596188
rect 674052 578172 674116 578236
rect 674788 576540 674852 576604
rect 675156 575724 675220 575788
rect 674972 574092 675036 574156
rect 675892 573684 675956 573748
rect 675708 573276 675772 573340
rect 676628 571916 676692 571980
rect 676444 571508 676508 571572
rect 676812 564436 676876 564500
rect 675708 562456 675772 562460
rect 675708 562400 675758 562456
rect 675758 562400 675772 562456
rect 675708 562396 675772 562400
rect 675892 561988 675956 562052
rect 674972 561172 675036 561236
rect 675156 558724 675220 558788
rect 676628 558316 676692 558380
rect 676444 557500 676508 557564
rect 43852 557228 43916 557292
rect 43668 556004 43732 556068
rect 39988 555460 40052 555524
rect 40172 555460 40236 555524
rect 41828 554780 41892 554844
rect 41460 540908 41524 540972
rect 41828 540772 41892 540836
rect 674420 531660 674484 531724
rect 675524 530980 675588 531044
rect 674236 530572 674300 530636
rect 676076 529348 676140 529412
rect 675340 528940 675404 529004
rect 674604 528532 674668 528596
rect 676260 527308 676324 527372
rect 676812 526900 676876 526964
rect 676444 492356 676508 492420
rect 676812 492356 676876 492420
rect 673684 489228 673748 489292
rect 674972 487596 675036 487660
rect 675708 486780 675772 486844
rect 675892 485148 675956 485212
rect 675156 484740 675220 484804
rect 676076 484468 676140 484532
rect 676812 482938 676876 483002
rect 43852 460124 43916 460188
rect 43852 459852 43916 459916
rect 43668 455908 43732 455972
rect 44036 455908 44100 455972
rect 43668 450740 43732 450804
rect 43668 445844 43732 445908
rect 44220 445844 44284 445908
rect 43668 430612 43732 430676
rect 43852 428844 43916 428908
rect 39988 427858 40052 427922
rect 40356 427790 40420 427854
rect 40034 427212 40098 427276
rect 673684 400964 673748 401028
rect 673868 400148 673932 400212
rect 40172 388996 40236 389060
rect 42932 386276 42996 386340
rect 41276 384644 41340 384708
rect 42748 383964 42812 384028
rect 39988 383828 40052 383892
rect 42748 383420 42812 383484
rect 39988 383012 40052 383076
rect 41276 383012 41340 383076
rect 41460 382196 41524 382260
rect 674052 357444 674116 357508
rect 674236 355812 674300 355876
rect 41460 355676 41524 355740
rect 674420 354996 674484 355060
rect 676076 353636 676140 353700
rect 675892 352140 675956 352204
rect 42932 351868 42996 351932
rect 675708 350508 675772 350572
rect 39988 341396 40052 341460
rect 42748 340444 42812 340508
rect 41828 340036 41892 340100
rect 42564 339220 42628 339284
rect 42012 338812 42076 338876
rect 41644 337316 41708 337380
rect 42196 337180 42260 337244
rect 42380 336772 42444 336836
rect 675708 330576 675772 330580
rect 675708 330520 675722 330576
rect 675722 330520 675772 330576
rect 675708 330516 675772 330520
rect 41460 329700 41524 329764
rect 676076 328340 676140 328404
rect 675892 326844 675956 326908
rect 41460 319908 41524 319972
rect 42380 316916 42444 316980
rect 42196 316296 42260 316300
rect 42196 316240 42210 316296
rect 42210 316240 42260 316296
rect 42196 316236 42260 316240
rect 42012 315616 42076 315620
rect 42012 315560 42026 315616
rect 42026 315560 42076 315616
rect 42012 315556 42076 315560
rect 41828 313848 41892 313852
rect 41828 313792 41878 313848
rect 41878 313792 41892 313848
rect 41828 313788 41892 313792
rect 41644 312972 41708 313036
rect 42564 312292 42628 312356
rect 675892 305900 675956 305964
rect 42380 300052 42444 300116
rect 41828 298420 41892 298484
rect 42196 297604 42260 297668
rect 42012 295564 42076 295628
rect 41828 295292 41892 295356
rect 42196 295292 42260 295356
rect 675892 291620 675956 291684
rect 41644 289172 41708 289236
rect 42380 289172 42444 289236
rect 42380 285908 42444 285972
rect 42196 285772 42260 285836
rect 42564 285636 42628 285700
rect 44036 278428 44100 278492
rect 673684 279628 673748 279692
rect 674052 279492 674116 279556
rect 674420 279356 674484 279420
rect 674236 279220 674300 279284
rect 673868 279084 673932 279148
rect 673500 278948 673564 279012
rect 42012 272368 42076 272372
rect 42012 272312 42026 272368
rect 42026 272312 42076 272368
rect 42012 272308 42076 272312
rect 42564 270404 42628 270468
rect 42380 269996 42444 270060
rect 42196 269376 42260 269380
rect 42196 269320 42210 269376
rect 42210 269320 42260 269376
rect 42196 269316 42260 269320
rect 674236 264556 674300 264620
rect 674236 262380 674300 262444
rect 675892 262380 675956 262444
rect 42196 256804 42260 256868
rect 41644 256260 41708 256324
rect 42012 255172 42076 255236
rect 41460 255036 41524 255100
rect 41460 254220 41524 254284
rect 41828 253948 41892 254012
rect 42012 252724 42076 252788
rect 42012 225992 42076 225996
rect 42012 225936 42026 225992
rect 42026 225936 42076 225992
rect 42012 225932 42076 225936
rect 676076 219948 676140 220012
rect 42196 213284 42260 213348
rect 41828 211652 41892 211716
rect 41460 210972 41524 211036
rect 42748 210428 42812 210492
rect 41828 209612 41892 209676
rect 42380 209204 42444 209268
rect 42564 208796 42628 208860
rect 41644 207708 41708 207772
rect 42012 207572 42076 207636
rect 42196 207164 42260 207228
rect 41460 205668 41524 205732
rect 42564 190164 42628 190228
rect 41460 187580 41524 187644
rect 42196 187096 42260 187100
rect 42196 187040 42210 187096
rect 42210 187040 42260 187096
rect 42196 187036 42260 187040
rect 42012 186416 42076 186420
rect 42012 186360 42026 186416
rect 42026 186360 42076 186416
rect 42012 186356 42076 186360
rect 42380 185812 42444 185876
rect 42748 184180 42812 184244
rect 41644 183636 41708 183700
rect 41828 182744 41892 182748
rect 41828 182688 41842 182744
rect 41842 182688 41892 182744
rect 41828 182684 41892 182688
rect 675892 173572 675956 173636
rect 676076 171804 676140 171868
rect 675708 170716 675772 170780
rect 675708 156496 675772 156500
rect 675708 156440 675758 156496
rect 675758 156440 675772 156496
rect 675708 156436 675772 156440
rect 675892 148412 675956 148476
rect 676076 146236 676140 146300
rect 675892 128420 675956 128484
rect 676076 126516 676140 126580
rect 580948 113188 581012 113252
rect 675892 103260 675956 103324
rect 676076 101356 676140 101420
rect 662092 95508 662156 95572
rect 662092 88768 662156 88772
rect 662092 88712 662142 88768
rect 662142 88712 662156 88768
rect 662092 88708 662156 88712
rect 580948 73476 581012 73540
rect 520412 48180 520476 48244
rect 520412 42120 520476 42124
rect 520412 42064 520462 42120
rect 520462 42064 520476 42120
rect 520412 42060 520476 42064
<< metal4 >>
rect 187739 997252 187805 997253
rect 187739 997188 187740 997252
rect 187804 997188 187805 997252
rect 187739 997187 187805 997188
rect 187742 995757 187802 997187
rect 187739 995756 187805 995757
rect 187739 995692 187740 995756
rect 187804 995692 187805 995756
rect 187739 995691 187805 995692
rect 638539 995212 638605 995213
rect 638539 995148 638540 995212
rect 638604 995148 638605 995212
rect 638539 995147 638605 995148
rect 638542 990589 638602 995147
rect 638539 990588 638605 990589
rect 638539 990524 638540 990588
rect 638604 990524 638605 990588
rect 638539 990523 638605 990524
rect 677171 985964 677237 985965
rect 677171 985900 677172 985964
rect 677236 985900 677237 985964
rect 677171 985899 677237 985900
rect 676987 985828 677053 985829
rect 676987 985764 676988 985828
rect 677052 985764 677053 985828
rect 676987 985763 677053 985764
rect 43667 985692 43733 985693
rect 43667 985628 43668 985692
rect 43732 985628 43733 985692
rect 43667 985627 43733 985628
rect 43483 985420 43549 985421
rect 43483 985356 43484 985420
rect 43548 985356 43549 985420
rect 43483 985355 43549 985356
rect 43299 982972 43365 982973
rect 43299 982908 43300 982972
rect 43364 982908 43365 982972
rect 43299 982907 43365 982908
rect 41459 968828 41525 968829
rect 41459 968764 41460 968828
rect 41524 968764 41525 968828
rect 41459 968763 41525 968764
rect 41462 937410 41522 968763
rect 41643 965156 41709 965157
rect 41643 965092 41644 965156
rect 41708 965092 41709 965156
rect 41643 965091 41709 965092
rect 41646 938090 41706 965091
rect 41827 963388 41893 963389
rect 41827 963324 41828 963388
rect 41892 963324 41893 963388
rect 41827 963323 41893 963324
rect 41830 949517 41890 963323
rect 41827 949516 41893 949517
rect 41827 949452 41828 949516
rect 41892 949452 41893 949516
rect 41827 949451 41893 949452
rect 41646 938030 42074 938090
rect 41462 937350 41890 937410
rect 41830 937005 41890 937350
rect 41827 937004 41893 937005
rect 41827 936940 41828 937004
rect 41892 936940 41893 937004
rect 41827 936939 41893 936940
rect 42014 935373 42074 938030
rect 42011 935372 42077 935373
rect 42011 935308 42012 935372
rect 42076 935308 42077 935372
rect 42011 935307 42077 935308
rect 43302 927213 43362 982907
rect 43299 927212 43365 927213
rect 43299 927148 43300 927212
rect 43364 927148 43365 927212
rect 43299 927147 43365 927148
rect 43486 922045 43546 985355
rect 43483 922044 43549 922045
rect 43483 921980 43484 922044
rect 43548 921980 43549 922044
rect 43483 921979 43549 921980
rect 39990 814270 41890 814330
rect 39990 773125 40050 814270
rect 41830 814197 41890 814270
rect 41827 814196 41893 814197
rect 41827 814132 41828 814196
rect 41892 814132 41893 814196
rect 41827 814131 41893 814132
rect 39987 773124 40053 773125
rect 39987 773060 39988 773124
rect 40052 773060 40053 773124
rect 39987 773059 40053 773060
rect 39987 771492 40053 771493
rect 39987 771428 39988 771492
rect 40052 771428 40053 771492
rect 39987 771427 40053 771428
rect 39990 731101 40050 771427
rect 41459 771084 41525 771085
rect 41459 771020 41460 771084
rect 41524 771020 41525 771084
rect 41459 771019 41525 771020
rect 39987 731100 40053 731101
rect 39987 731036 39988 731100
rect 40052 731036 40053 731100
rect 39987 731035 40053 731036
rect 41275 686764 41341 686765
rect 41275 686700 41276 686764
rect 41340 686700 41341 686764
rect 41275 686699 41341 686700
rect 41278 684317 41338 686699
rect 39987 684316 40053 684317
rect 39987 684252 39988 684316
rect 40052 684252 40053 684316
rect 39987 684251 40053 684252
rect 41275 684316 41341 684317
rect 41275 684252 41276 684316
rect 41340 684252 41341 684316
rect 41275 684251 41341 684252
rect 39990 643517 40050 684251
rect 39987 643516 40053 643517
rect 39987 643452 39988 643516
rect 40052 643452 40053 643516
rect 39987 643451 40053 643452
rect 40171 598636 40237 598637
rect 40171 598572 40172 598636
rect 40236 598572 40237 598636
rect 40171 598571 40237 598572
rect 40174 596189 40234 598571
rect 40171 596188 40237 596189
rect 40171 596124 40172 596188
rect 40236 596124 40237 596188
rect 40171 596123 40237 596124
rect 40174 555525 40234 596123
rect 39987 555524 40053 555525
rect 39987 555460 39988 555524
rect 40052 555460 40053 555524
rect 39987 555459 40053 555460
rect 40171 555524 40237 555525
rect 40171 555460 40172 555524
rect 40236 555460 40237 555524
rect 40171 555459 40237 555460
rect 39990 427923 40050 555459
rect 41462 540973 41522 771019
rect 43299 757756 43365 757757
rect 43299 757692 43300 757756
rect 43364 757692 43365 757756
rect 43299 757691 43365 757692
rect 41827 757076 41893 757077
rect 41827 757012 41828 757076
rect 41892 757012 41893 757076
rect 41827 757011 41893 757012
rect 42195 757076 42261 757077
rect 42195 757012 42196 757076
rect 42260 757012 42261 757076
rect 42195 757011 42261 757012
rect 41830 754085 41890 757011
rect 42198 755309 42258 757011
rect 42195 755308 42261 755309
rect 42195 755244 42196 755308
rect 42260 755244 42261 755308
rect 42195 755243 42261 755244
rect 41827 754084 41893 754085
rect 41827 754020 41828 754084
rect 41892 754020 41893 754084
rect 41827 754019 41893 754020
rect 43302 752997 43362 757691
rect 43299 752996 43365 752997
rect 43299 752932 43300 752996
rect 43364 752932 43365 752996
rect 43299 752931 43365 752932
rect 43670 643517 43730 985627
rect 44035 985556 44101 985557
rect 44035 985492 44036 985556
rect 44100 985492 44101 985556
rect 44035 985491 44101 985492
rect 43851 983108 43917 983109
rect 43851 983044 43852 983108
rect 43916 983044 43917 983108
rect 43851 983043 43917 983044
rect 43667 643516 43733 643517
rect 43667 643452 43668 643516
rect 43732 643452 43733 643516
rect 43667 643451 43733 643452
rect 43854 598093 43914 983043
rect 44038 685269 44098 985491
rect 676990 981612 677050 985763
rect 674790 981552 677050 981612
rect 673867 938364 673933 938365
rect 673867 938300 673868 938364
rect 673932 938300 673933 938364
rect 673867 938299 673933 938300
rect 673870 760341 673930 938299
rect 674790 936325 674850 981552
rect 677174 981356 677234 985899
rect 674974 981296 677234 981356
rect 674974 937141 675034 981296
rect 676811 937276 676877 937277
rect 676811 937212 676812 937276
rect 676876 937212 676877 937276
rect 676811 937211 676877 937212
rect 674971 937140 675037 937141
rect 674971 937076 674972 937140
rect 675036 937076 675037 937140
rect 674971 937075 675037 937076
rect 674787 936324 674853 936325
rect 674787 936260 674788 936324
rect 674852 936260 674853 936324
rect 674787 936259 674853 936260
rect 676075 877300 676141 877301
rect 676075 877236 676076 877300
rect 676140 877236 676141 877300
rect 676075 877235 676141 877236
rect 675707 876620 675773 876621
rect 675707 876556 675708 876620
rect 675772 876556 675773 876620
rect 675707 876555 675773 876556
rect 675523 875940 675589 875941
rect 675523 875876 675524 875940
rect 675588 875876 675589 875940
rect 675523 875875 675589 875876
rect 675339 874036 675405 874037
rect 675339 873972 675340 874036
rect 675404 873972 675405 874036
rect 675339 873971 675405 873972
rect 674971 787812 675037 787813
rect 674971 787748 674972 787812
rect 675036 787748 675037 787812
rect 674971 787747 675037 787748
rect 674603 787268 674669 787269
rect 674603 787204 674604 787268
rect 674668 787204 674669 787268
rect 674603 787203 674669 787204
rect 674419 786860 674485 786861
rect 674419 786796 674420 786860
rect 674484 786796 674485 786860
rect 674419 786795 674485 786796
rect 674235 777476 674301 777477
rect 674235 777412 674236 777476
rect 674300 777412 674301 777476
rect 674235 777411 674301 777412
rect 674238 773397 674298 777411
rect 674235 773396 674301 773397
rect 674235 773332 674236 773396
rect 674300 773332 674301 773396
rect 674235 773331 674301 773332
rect 673867 760340 673933 760341
rect 673867 760276 673868 760340
rect 673932 760276 673933 760340
rect 673867 760275 673933 760276
rect 674051 741708 674117 741709
rect 674051 741644 674052 741708
rect 674116 741644 674117 741708
rect 674051 741643 674117 741644
rect 673867 739804 673933 739805
rect 673867 739740 673868 739804
rect 673932 739740 673933 739804
rect 673867 739739 673933 739740
rect 673683 739124 673749 739125
rect 673683 739060 673684 739124
rect 673748 739060 673749 739124
rect 673683 739059 673749 739060
rect 673499 693700 673565 693701
rect 673499 693636 673500 693700
rect 673564 693636 673565 693700
rect 673499 693635 673565 693636
rect 44035 685268 44101 685269
rect 44035 685204 44036 685268
rect 44100 685204 44101 685268
rect 44035 685203 44101 685204
rect 673502 618629 673562 693635
rect 673686 664053 673746 739059
rect 673870 665685 673930 739739
rect 674054 666909 674114 741643
rect 674422 712061 674482 786795
rect 674419 712060 674485 712061
rect 674419 711996 674420 712060
rect 674484 711996 674485 712060
rect 674419 711995 674485 711996
rect 674606 709613 674666 787203
rect 674787 783868 674853 783869
rect 674787 783804 674788 783868
rect 674852 783804 674853 783868
rect 674787 783803 674853 783804
rect 674603 709612 674669 709613
rect 674603 709548 674604 709612
rect 674668 709548 674669 709612
rect 674603 709547 674669 709548
rect 674790 708797 674850 783803
rect 674974 711245 675034 787747
rect 675155 784140 675221 784141
rect 675155 784076 675156 784140
rect 675220 784076 675221 784140
rect 675155 784075 675221 784076
rect 674971 711244 675037 711245
rect 674971 711180 674972 711244
rect 675036 711180 675037 711244
rect 674971 711179 675037 711180
rect 675158 709205 675218 784075
rect 675342 766862 675402 873971
rect 675526 767046 675586 875875
rect 675710 767230 675770 876555
rect 675891 872268 675957 872269
rect 675891 872204 675892 872268
rect 675956 872204 675957 872268
rect 675891 872203 675957 872204
rect 675894 767414 675954 872203
rect 676078 767598 676138 877235
rect 676259 797740 676325 797741
rect 676259 797676 676260 797740
rect 676324 797676 676325 797740
rect 676259 797675 676325 797676
rect 676262 767782 676322 797675
rect 676443 792028 676509 792029
rect 676443 791964 676444 792028
rect 676508 791964 676509 792028
rect 676443 791963 676509 791964
rect 676446 767966 676506 791963
rect 676814 772717 676874 937211
rect 676811 772716 676877 772717
rect 676811 772652 676812 772716
rect 676876 772652 676877 772716
rect 676811 772651 676877 772652
rect 676446 767906 677836 767966
rect 676262 767722 677652 767782
rect 676078 767538 677468 767598
rect 675894 767354 677284 767414
rect 675710 767170 677100 767230
rect 675526 766986 676916 767046
rect 675342 766802 676732 766862
rect 676672 764770 676732 766802
rect 675342 764710 676732 764770
rect 675342 755853 675402 764710
rect 676856 764586 676916 766986
rect 675526 764526 676916 764586
rect 675526 757077 675586 764526
rect 677040 764402 677100 767170
rect 675710 764342 677100 764402
rect 675523 757076 675589 757077
rect 675523 757012 675524 757076
rect 675588 757012 675589 757076
rect 675523 757011 675589 757012
rect 675339 755852 675405 755853
rect 675339 755788 675340 755852
rect 675404 755788 675405 755852
rect 675339 755787 675405 755788
rect 675710 754629 675770 764342
rect 677224 764218 677284 767354
rect 675894 764158 677284 764218
rect 675707 754628 675773 754629
rect 675707 754564 675708 754628
rect 675772 754564 675773 754628
rect 675707 754563 675773 754564
rect 675894 752589 675954 764158
rect 677408 764034 677468 767538
rect 676078 763974 677468 764034
rect 676078 756397 676138 763974
rect 677592 763850 677652 767722
rect 676262 763790 677652 763850
rect 676075 756396 676141 756397
rect 676075 756332 676076 756396
rect 676140 756332 676141 756396
rect 676075 756331 676141 756332
rect 675891 752588 675957 752589
rect 675891 752524 675892 752588
rect 675956 752524 675957 752588
rect 675891 752523 675957 752524
rect 676262 751909 676322 763790
rect 677776 763666 677836 767906
rect 676446 763606 677836 763666
rect 676446 752317 676506 763606
rect 676443 752316 676509 752317
rect 676443 752252 676444 752316
rect 676508 752252 676509 752316
rect 676443 752251 676509 752252
rect 676259 751908 676325 751909
rect 676259 751844 676260 751908
rect 676324 751844 676325 751908
rect 676259 751843 676325 751844
rect 676627 744156 676693 744157
rect 676627 744092 676628 744156
rect 676692 744092 676693 744156
rect 676627 744091 676693 744092
rect 676259 744020 676325 744021
rect 676259 743956 676260 744020
rect 676324 743956 676325 744020
rect 676259 743955 676325 743956
rect 675891 742932 675957 742933
rect 675891 742868 675892 742932
rect 675956 742868 675957 742932
rect 675891 742867 675957 742868
rect 675707 738580 675773 738581
rect 675707 738516 675708 738580
rect 675772 738516 675773 738580
rect 675707 738515 675773 738516
rect 675710 722359 675770 738515
rect 675894 722543 675954 742867
rect 676075 742524 676141 742525
rect 676075 742460 676076 742524
rect 676140 742460 676141 742524
rect 676075 742459 676141 742460
rect 676078 722727 676138 742459
rect 676262 722911 676322 743955
rect 676443 738036 676509 738037
rect 676443 737972 676444 738036
rect 676508 737972 676509 738036
rect 676443 737971 676509 737972
rect 676446 723095 676506 737971
rect 676630 723279 676690 744091
rect 676630 723219 677769 723279
rect 676446 723035 677585 723095
rect 676262 722851 677401 722911
rect 676078 722667 677217 722727
rect 675894 722483 677033 722543
rect 675710 722299 676849 722359
rect 676789 719460 676849 722299
rect 675710 719400 676849 719460
rect 675155 709204 675221 709205
rect 675155 709140 675156 709204
rect 675220 709140 675221 709204
rect 675155 709139 675221 709140
rect 674787 708796 674853 708797
rect 674787 708732 674788 708796
rect 674852 708732 674853 708796
rect 674787 708731 674853 708732
rect 675523 698188 675589 698189
rect 675523 698124 675524 698188
rect 675588 698124 675589 698188
rect 675523 698123 675589 698124
rect 675339 697236 675405 697237
rect 675339 697172 675340 697236
rect 675404 697172 675405 697236
rect 675339 697171 675405 697172
rect 674235 696692 674301 696693
rect 674235 696628 674236 696692
rect 674300 696628 674301 696692
rect 674235 696627 674301 696628
rect 674051 666908 674117 666909
rect 674051 666844 674052 666908
rect 674116 666844 674117 666908
rect 674051 666843 674117 666844
rect 673867 665684 673933 665685
rect 673867 665620 673868 665684
rect 673932 665620 673933 665684
rect 673867 665619 673933 665620
rect 673683 664052 673749 664053
rect 673683 663988 673684 664052
rect 673748 663988 673749 664052
rect 673683 663987 673749 663988
rect 673683 623116 673749 623117
rect 673683 623052 673684 623116
rect 673748 623052 673749 623116
rect 673683 623051 673749 623052
rect 673686 621621 673746 623051
rect 674238 621893 674298 696627
rect 674419 695060 674485 695061
rect 674419 694996 674420 695060
rect 674484 694996 674485 695060
rect 674419 694995 674485 694996
rect 674235 621892 674301 621893
rect 674235 621828 674236 621892
rect 674300 621828 674301 621892
rect 674235 621827 674301 621828
rect 673683 621620 673749 621621
rect 673683 621556 673684 621620
rect 673748 621556 673749 621620
rect 673683 621555 673749 621556
rect 673499 618628 673565 618629
rect 673499 618564 673500 618628
rect 673564 618564 673565 618628
rect 673499 618563 673565 618564
rect 673686 612750 673746 621555
rect 674422 620669 674482 694995
rect 674603 694244 674669 694245
rect 674603 694180 674604 694244
rect 674668 694180 674669 694244
rect 674603 694179 674669 694180
rect 674419 620668 674485 620669
rect 674419 620604 674420 620668
rect 674484 620604 674485 620668
rect 674419 620603 674485 620604
rect 674606 619037 674666 694179
rect 675342 676990 675402 697171
rect 674750 676930 675402 676990
rect 674750 673598 674810 676930
rect 675526 676836 675586 698123
rect 674904 676776 675586 676836
rect 674904 673782 674964 676776
rect 675710 676692 675770 719400
rect 676973 719276 677033 722483
rect 675048 676632 675770 676692
rect 675894 719216 677033 719276
rect 675048 673966 675108 676632
rect 675894 676548 675954 719216
rect 677157 719092 677217 722667
rect 676078 719032 677217 719092
rect 676078 676786 676138 719032
rect 677341 718908 677401 722851
rect 676262 718848 677401 718908
rect 676262 711891 676322 718848
rect 677525 718724 677585 723035
rect 676446 718664 677585 718724
rect 676259 711890 676325 711891
rect 676259 711826 676260 711890
rect 676324 711826 676325 711890
rect 676259 711825 676325 711826
rect 676259 699684 676325 699685
rect 676259 699620 676260 699684
rect 676324 699620 676325 699684
rect 676259 699619 676325 699620
rect 676262 676970 676322 699619
rect 676446 678688 676506 718664
rect 677709 718540 677769 723219
rect 676630 718480 677769 718540
rect 676630 714870 676690 718480
rect 676630 714810 677058 714870
rect 676998 711891 677058 714810
rect 676995 711890 677061 711891
rect 676995 711826 676996 711890
rect 677060 711826 677061 711890
rect 676995 711825 677061 711826
rect 676811 699820 676877 699821
rect 676811 699756 676812 699820
rect 676876 699756 676877 699820
rect 676811 699755 676877 699756
rect 676627 690164 676693 690165
rect 676627 690100 676628 690164
rect 676692 690100 676693 690164
rect 676627 690099 676693 690100
rect 676446 678657 676507 678688
rect 676447 677154 676507 678657
rect 676630 677294 676690 690099
rect 676814 677458 676874 699755
rect 676995 699548 677061 699549
rect 676995 699484 676996 699548
rect 677060 699484 677061 699548
rect 676995 699483 677061 699484
rect 676998 677642 677058 699483
rect 677179 693020 677245 693021
rect 677179 692956 677180 693020
rect 677244 692956 677245 693020
rect 677179 692955 677245 692956
rect 677182 681730 677242 692955
rect 677182 681670 677776 681730
rect 676998 677582 677609 677642
rect 676814 677398 677425 677458
rect 676630 677234 677261 677294
rect 676447 677094 677121 677154
rect 676262 676910 676937 676970
rect 676078 676726 676753 676786
rect 675192 676488 675954 676548
rect 675192 674150 675252 676488
rect 676693 674542 676753 676726
rect 676078 674482 676753 674542
rect 675192 674090 675954 674150
rect 675048 673906 675770 673966
rect 674904 673722 675586 673782
rect 674750 673538 675402 673598
rect 675155 652628 675221 652629
rect 675155 652564 675156 652628
rect 675220 652564 675221 652628
rect 675155 652563 675221 652564
rect 674971 652220 675037 652221
rect 674971 652156 674972 652220
rect 675036 652156 675037 652220
rect 674971 652155 675037 652156
rect 674787 651676 674853 651677
rect 674787 651612 674788 651676
rect 674852 651612 674853 651676
rect 674787 651611 674853 651612
rect 674603 619036 674669 619037
rect 674603 618972 674604 619036
rect 674668 618972 674669 619036
rect 674603 618971 674669 618972
rect 673686 612690 674114 612750
rect 43851 598092 43917 598093
rect 43851 598028 43852 598092
rect 43916 598028 43917 598092
rect 43851 598027 43917 598028
rect 674054 578237 674114 612690
rect 674419 606524 674485 606525
rect 674419 606460 674420 606524
rect 674484 606460 674485 606524
rect 674419 606459 674485 606460
rect 674235 604756 674301 604757
rect 674235 604692 674236 604756
rect 674300 604692 674301 604756
rect 674235 604691 674301 604692
rect 674051 578236 674117 578237
rect 674051 578172 674052 578236
rect 674116 578172 674117 578236
rect 674051 578171 674117 578172
rect 43851 557292 43917 557293
rect 43851 557228 43852 557292
rect 43916 557228 43917 557292
rect 43851 557227 43917 557228
rect 43667 556068 43733 556069
rect 43667 556004 43668 556068
rect 43732 556004 43733 556068
rect 43667 556003 43733 556004
rect 41827 554844 41893 554845
rect 41827 554780 41828 554844
rect 41892 554780 41893 554844
rect 41827 554779 41893 554780
rect 41459 540972 41525 540973
rect 41459 540908 41460 540972
rect 41524 540908 41525 540972
rect 41459 540907 41525 540908
rect 41830 540837 41890 554779
rect 41827 540836 41893 540837
rect 41827 540772 41828 540836
rect 41892 540772 41893 540836
rect 41827 540771 41893 540772
rect 43670 455973 43730 556003
rect 43854 460189 43914 557227
rect 674238 543933 674298 604691
rect 673151 543873 674298 543933
rect 673151 536896 673211 543873
rect 674422 543749 674482 606459
rect 674603 603532 674669 603533
rect 674603 603468 674604 603532
rect 674668 603468 674669 603532
rect 674603 603467 674669 603468
rect 673335 543689 674482 543749
rect 673335 537080 673395 543689
rect 674606 543565 674666 603467
rect 674790 576605 674850 651611
rect 674787 576604 674853 576605
rect 674787 576540 674788 576604
rect 674852 576540 674853 576604
rect 674787 576539 674853 576540
rect 674974 574157 675034 652155
rect 675158 575789 675218 652563
rect 675342 631488 675402 673538
rect 675526 631672 675586 673722
rect 675710 663645 675770 673906
rect 675894 666093 675954 674090
rect 675891 666092 675957 666093
rect 675891 666028 675892 666092
rect 675956 666028 675957 666092
rect 675891 666027 675957 666028
rect 676078 664597 676138 674482
rect 676877 674358 676937 676910
rect 676262 674298 676937 674358
rect 676075 664596 676141 664597
rect 676075 664532 676076 664596
rect 676140 664532 676141 664596
rect 676075 664531 676141 664532
rect 675707 663644 675773 663645
rect 675707 663580 675708 663644
rect 675772 663580 675773 663644
rect 675707 663579 675773 663580
rect 676262 662965 676322 674298
rect 677061 674174 677121 677094
rect 676446 674114 677121 674174
rect 676259 662964 676325 662965
rect 676259 662900 676260 662964
rect 676324 662900 676325 662964
rect 676259 662899 676325 662900
rect 676446 662557 676506 674114
rect 677201 673990 677261 677234
rect 676630 673930 677261 673990
rect 676443 662556 676509 662557
rect 676443 662492 676444 662556
rect 676508 662492 676509 662556
rect 676443 662491 676509 662492
rect 675891 649228 675957 649229
rect 675891 649164 675892 649228
rect 675956 649164 675957 649228
rect 675891 649163 675957 649164
rect 675707 648684 675773 648685
rect 675707 648620 675708 648684
rect 675772 648620 675773 648684
rect 675707 648619 675773 648620
rect 675710 631856 675770 648619
rect 675894 632040 675954 649163
rect 676630 632180 676690 673930
rect 677365 673806 677425 677398
rect 676814 673746 677425 673806
rect 676814 661741 676874 673746
rect 677549 673622 677609 677582
rect 676998 673562 677609 673622
rect 676998 662149 677058 673562
rect 677716 673330 677776 681670
rect 677182 673270 677776 673330
rect 676995 662148 677061 662149
rect 676995 662084 676996 662148
rect 677060 662084 677061 662148
rect 676995 662083 677061 662084
rect 676811 661740 676877 661741
rect 676811 661676 676812 661740
rect 676876 661676 676877 661740
rect 676811 661675 676877 661676
rect 677182 632336 677242 673270
rect 677363 667044 677429 667045
rect 677363 666980 677364 667044
rect 677428 666980 677429 667044
rect 677363 666979 677429 666980
rect 677366 632477 677426 666979
rect 677366 632417 677748 632477
rect 677182 632276 677571 632336
rect 676630 632120 677410 632180
rect 675894 631980 677240 632040
rect 675710 631796 677056 631856
rect 675526 631612 676882 631672
rect 675342 631428 676708 631488
rect 676648 629787 676708 631428
rect 675342 629727 676708 629787
rect 675342 619445 675402 629727
rect 676822 629603 676882 631612
rect 675526 629543 676882 629603
rect 675526 621077 675586 629543
rect 676996 629419 677056 631796
rect 675710 629359 677056 629419
rect 675523 621076 675589 621077
rect 675523 621012 675524 621076
rect 675588 621012 675589 621076
rect 675523 621011 675589 621012
rect 675339 619444 675405 619445
rect 675339 619380 675340 619444
rect 675404 619380 675405 619444
rect 675339 619379 675405 619380
rect 675523 607612 675589 607613
rect 675523 607548 675524 607612
rect 675588 607548 675589 607612
rect 675523 607547 675589 607548
rect 675339 604348 675405 604349
rect 675339 604284 675340 604348
rect 675404 604284 675405 604348
rect 675339 604283 675405 604284
rect 675342 587486 675402 604283
rect 675526 587670 675586 607547
rect 675710 587854 675770 629359
rect 677180 629235 677240 631980
rect 675894 629175 677240 629235
rect 675894 588038 675954 629175
rect 677350 628952 677410 632120
rect 676630 628892 677410 628952
rect 676259 622436 676325 622437
rect 676259 622372 676260 622436
rect 676324 622372 676325 622436
rect 676259 622371 676325 622372
rect 676262 619850 676322 622371
rect 676078 619790 676322 619850
rect 676078 619581 676138 619790
rect 676075 619580 676141 619581
rect 676075 619516 676076 619580
rect 676140 619516 676141 619580
rect 676075 619515 676141 619516
rect 676630 617133 676690 628892
rect 677511 628792 677571 632276
rect 677182 628732 677571 628792
rect 677182 617541 677242 628732
rect 677688 628634 677748 632417
rect 677366 628574 677748 628634
rect 677366 622845 677426 628574
rect 677363 622844 677429 622845
rect 677363 622780 677364 622844
rect 677428 622780 677429 622844
rect 677363 622779 677429 622780
rect 677179 617540 677245 617541
rect 677179 617476 677180 617540
rect 677244 617476 677245 617540
rect 677179 617475 677245 617476
rect 676627 617132 676693 617133
rect 676627 617068 676628 617132
rect 676692 617068 676693 617132
rect 676627 617067 676693 617068
rect 676443 607748 676509 607749
rect 676443 607684 676444 607748
rect 676508 607684 676509 607748
rect 676443 607683 676509 607684
rect 676075 607340 676141 607341
rect 676075 607276 676076 607340
rect 676140 607276 676141 607340
rect 676075 607275 676141 607276
rect 676078 588222 676138 607275
rect 676259 602988 676325 602989
rect 676259 602924 676260 602988
rect 676324 602924 676325 602988
rect 676259 602923 676325 602924
rect 676262 588406 676322 602923
rect 676446 588590 676506 607683
rect 676627 607476 676693 607477
rect 676627 607412 676628 607476
rect 676692 607412 676693 607476
rect 676627 607411 676693 607412
rect 676630 588774 676690 607411
rect 676630 588714 677821 588774
rect 676446 588530 677667 588590
rect 676262 588346 677493 588406
rect 676078 588162 677351 588222
rect 675894 587978 677192 588038
rect 675710 587794 677028 587854
rect 675526 587610 676864 587670
rect 675342 587426 676700 587486
rect 676640 583686 676700 587426
rect 675342 583626 676700 583686
rect 675155 575788 675221 575789
rect 675155 575724 675156 575788
rect 675220 575724 675221 575788
rect 675155 575723 675221 575724
rect 674971 574156 675037 574157
rect 674971 574092 674972 574156
rect 675036 574092 675037 574156
rect 674971 574091 675037 574092
rect 674971 561236 675037 561237
rect 674971 561172 674972 561236
rect 675036 561172 675037 561236
rect 674971 561171 675037 561172
rect 673519 543505 674666 543565
rect 673519 537264 673579 543505
rect 674974 543239 675034 561171
rect 675155 558788 675221 558789
rect 675155 558724 675156 558788
rect 675220 558724 675221 558788
rect 675155 558723 675221 558724
rect 673733 543179 675034 543239
rect 673733 537742 673793 543179
rect 675158 543055 675218 558723
rect 673917 542995 675218 543055
rect 673917 537926 673977 542995
rect 675342 542871 675402 583626
rect 676804 583502 676864 587610
rect 674101 542811 675402 542871
rect 675526 583442 676864 583502
rect 674101 538110 674161 542811
rect 675526 542687 675586 583442
rect 676968 583318 677028 587794
rect 675710 583258 677028 583318
rect 675710 573341 675770 583258
rect 677132 583134 677192 587978
rect 675894 583074 677192 583134
rect 675894 573749 675954 583074
rect 677291 582950 677351 588162
rect 676078 582890 677351 582950
rect 675891 573748 675957 573749
rect 675891 573684 675892 573748
rect 675956 573684 675957 573748
rect 675891 573683 675957 573684
rect 675707 573340 675773 573341
rect 675707 573276 675708 573340
rect 675772 573276 675773 573340
rect 675707 573275 675773 573276
rect 675707 562460 675773 562461
rect 675707 562396 675708 562460
rect 675772 562396 675773 562460
rect 675707 562395 675773 562396
rect 674285 542627 675586 542687
rect 674285 538294 674345 542627
rect 675710 542503 675770 562395
rect 675891 562052 675957 562053
rect 675891 561988 675892 562052
rect 675956 561988 675957 562052
rect 675891 561987 675957 561988
rect 674488 542443 675770 542503
rect 674488 538478 674548 542443
rect 675894 542319 675954 561987
rect 674672 542259 675954 542319
rect 674672 538662 674732 542259
rect 676078 542135 676138 582890
rect 677433 582766 677493 588346
rect 674856 542075 676138 542135
rect 676262 582706 677493 582766
rect 674856 538846 674916 542075
rect 676262 541951 676322 582706
rect 677607 582582 677667 588530
rect 676446 582522 677667 582582
rect 676446 571573 676506 582522
rect 677761 582398 677821 588714
rect 676630 582338 677821 582398
rect 676630 571981 676690 582338
rect 676627 571980 676693 571981
rect 676627 571916 676628 571980
rect 676692 571916 676693 571980
rect 676627 571915 676693 571916
rect 676443 571572 676509 571573
rect 676443 571508 676444 571572
rect 676508 571508 676509 571572
rect 676443 571507 676509 571508
rect 676811 564500 676877 564501
rect 676811 564436 676812 564500
rect 676876 564436 676877 564500
rect 676811 564435 676877 564436
rect 676627 558380 676693 558381
rect 676627 558316 676628 558380
rect 676692 558316 676693 558380
rect 676627 558315 676693 558316
rect 676443 557564 676509 557565
rect 676443 557500 676444 557564
rect 676508 557500 676509 557564
rect 676443 557499 676509 557500
rect 675040 541891 676322 541951
rect 675040 539030 675100 541891
rect 676446 541347 676506 557499
rect 676630 541531 676690 558315
rect 676814 541715 676874 564435
rect 676814 541655 677431 541715
rect 676630 541471 677247 541531
rect 676446 541287 677063 541347
rect 677003 539466 677063 541287
rect 676446 539406 677063 539466
rect 675040 538970 676322 539030
rect 674856 538786 676138 538846
rect 674672 538602 675954 538662
rect 674488 538418 675770 538478
rect 674285 538234 675586 538294
rect 674101 538050 675402 538110
rect 673917 537866 675218 537926
rect 673733 537682 675034 537742
rect 673519 537204 674666 537264
rect 673335 537020 674482 537080
rect 673151 536836 674298 536896
rect 674238 530637 674298 536836
rect 674422 531725 674482 537020
rect 674419 531724 674485 531725
rect 674419 531660 674420 531724
rect 674484 531660 674485 531724
rect 674419 531659 674485 531660
rect 674235 530636 674301 530637
rect 674235 530572 674236 530636
rect 674300 530572 674301 530636
rect 674235 530571 674301 530572
rect 674606 528597 674666 537204
rect 674603 528596 674669 528597
rect 674603 528532 674604 528596
rect 674668 528532 674669 528596
rect 674603 528531 674669 528532
rect 673683 489292 673749 489293
rect 673683 489228 673684 489292
rect 673748 489228 673749 489292
rect 673683 489227 673749 489228
rect 43851 460188 43917 460189
rect 43851 460124 43852 460188
rect 43916 460124 43917 460188
rect 43851 460123 43917 460124
rect 43851 459916 43917 459917
rect 43851 459852 43852 459916
rect 43916 459852 43917 459916
rect 43851 459851 43917 459852
rect 43667 455972 43733 455973
rect 43667 455908 43668 455972
rect 43732 455908 43733 455972
rect 43667 455907 43733 455908
rect 43667 450804 43733 450805
rect 43667 450740 43668 450804
rect 43732 450740 43733 450804
rect 43667 450739 43733 450740
rect 43670 445909 43730 450739
rect 43667 445908 43733 445909
rect 43667 445844 43668 445908
rect 43732 445844 43733 445908
rect 43667 445843 43733 445844
rect 43854 440330 43914 459851
rect 44035 455972 44101 455973
rect 44035 455908 44036 455972
rect 44100 455908 44101 455972
rect 44035 455907 44101 455908
rect 43670 440270 43914 440330
rect 43670 430677 43730 440270
rect 44038 439650 44098 455907
rect 44219 445908 44285 445909
rect 44219 445844 44220 445908
rect 44284 445844 44285 445908
rect 44219 445843 44285 445844
rect 43854 439590 44098 439650
rect 43667 430676 43733 430677
rect 43667 430612 43668 430676
rect 43732 430612 43733 430676
rect 43667 430611 43733 430612
rect 43854 428909 43914 439590
rect 44222 438970 44282 445843
rect 44038 438910 44282 438970
rect 43851 428908 43917 428909
rect 43851 428844 43852 428908
rect 43916 428844 43917 428908
rect 43851 428843 43917 428844
rect 39987 427922 40053 427923
rect 39987 427858 39988 427922
rect 40052 427858 40053 427922
rect 39987 427857 40053 427858
rect 40355 427854 40421 427855
rect 40355 427790 40356 427854
rect 40420 427790 40421 427854
rect 40355 427789 40421 427790
rect 39990 427277 40096 427410
rect 39990 427276 40099 427277
rect 39990 427212 40034 427276
rect 40098 427212 40099 427276
rect 39990 427211 40099 427212
rect 39990 383893 40050 427211
rect 40358 425070 40418 427789
rect 40174 425010 40418 425070
rect 40174 411270 40234 425010
rect 40174 411210 40418 411270
rect 40358 400230 40418 411210
rect 40174 400170 40418 400230
rect 40174 389061 40234 400170
rect 40171 389060 40237 389061
rect 40171 388996 40172 389060
rect 40236 388996 40237 389060
rect 40171 388995 40237 388996
rect 42931 386340 42997 386341
rect 42931 386276 42932 386340
rect 42996 386276 42997 386340
rect 42931 386275 42997 386276
rect 41275 384708 41341 384709
rect 41275 384644 41276 384708
rect 41340 384644 41341 384708
rect 41275 384643 41341 384644
rect 39987 383892 40053 383893
rect 39987 383828 39988 383892
rect 40052 383828 40053 383892
rect 39987 383827 40053 383828
rect 41278 383077 41338 384643
rect 42747 384028 42813 384029
rect 42747 383964 42748 384028
rect 42812 383964 42813 384028
rect 42747 383963 42813 383964
rect 42750 383485 42810 383963
rect 42747 383484 42813 383485
rect 42747 383420 42748 383484
rect 42812 383420 42813 383484
rect 42747 383419 42813 383420
rect 39987 383076 40053 383077
rect 39987 383012 39988 383076
rect 40052 383012 40053 383076
rect 39987 383011 40053 383012
rect 41275 383076 41341 383077
rect 41275 383012 41276 383076
rect 41340 383012 41341 383076
rect 41275 383011 41341 383012
rect 39990 341461 40050 383011
rect 41459 382260 41525 382261
rect 41459 382196 41460 382260
rect 41524 382196 41525 382260
rect 41459 382195 41525 382196
rect 41462 355741 41522 382195
rect 41459 355740 41525 355741
rect 41459 355676 41460 355740
rect 41524 355676 41525 355740
rect 41459 355675 41525 355676
rect 39987 341460 40053 341461
rect 39987 341396 39988 341460
rect 40052 341396 40053 341460
rect 39987 341395 40053 341396
rect 42750 340509 42810 383419
rect 42934 351933 42994 386275
rect 42931 351932 42997 351933
rect 42931 351868 42932 351932
rect 42996 351868 42997 351932
rect 42931 351867 42997 351868
rect 42747 340508 42813 340509
rect 42747 340444 42748 340508
rect 42812 340444 42813 340508
rect 42747 340443 42813 340444
rect 41827 340100 41893 340101
rect 41827 340036 41828 340100
rect 41892 340036 41893 340100
rect 41827 340035 41893 340036
rect 41643 337380 41709 337381
rect 41643 337316 41644 337380
rect 41708 337316 41709 337380
rect 41643 337315 41709 337316
rect 41459 329764 41525 329765
rect 41459 329700 41460 329764
rect 41524 329700 41525 329764
rect 41459 329699 41525 329700
rect 41462 319973 41522 329699
rect 41459 319972 41525 319973
rect 41459 319908 41460 319972
rect 41524 319908 41525 319972
rect 41459 319907 41525 319908
rect 41646 313037 41706 337315
rect 41830 313853 41890 340035
rect 42563 339284 42629 339285
rect 42563 339220 42564 339284
rect 42628 339220 42629 339284
rect 42563 339219 42629 339220
rect 42011 338876 42077 338877
rect 42011 338812 42012 338876
rect 42076 338812 42077 338876
rect 42011 338811 42077 338812
rect 42014 315621 42074 338811
rect 42195 337244 42261 337245
rect 42195 337180 42196 337244
rect 42260 337180 42261 337244
rect 42195 337179 42261 337180
rect 42198 316301 42258 337179
rect 42379 336836 42445 336837
rect 42379 336772 42380 336836
rect 42444 336772 42445 336836
rect 42379 336771 42445 336772
rect 42382 316981 42442 336771
rect 42379 316980 42445 316981
rect 42379 316916 42380 316980
rect 42444 316916 42445 316980
rect 42379 316915 42445 316916
rect 42195 316300 42261 316301
rect 42195 316236 42196 316300
rect 42260 316236 42261 316300
rect 42195 316235 42261 316236
rect 42011 315620 42077 315621
rect 42011 315556 42012 315620
rect 42076 315556 42077 315620
rect 42011 315555 42077 315556
rect 41827 313852 41893 313853
rect 41827 313788 41828 313852
rect 41892 313788 41893 313852
rect 41827 313787 41893 313788
rect 41643 313036 41709 313037
rect 41643 312972 41644 313036
rect 41708 312972 41709 313036
rect 41643 312971 41709 312972
rect 42566 312357 42626 339219
rect 42563 312356 42629 312357
rect 42563 312292 42564 312356
rect 42628 312292 42629 312356
rect 42563 312291 42629 312292
rect 42379 300116 42445 300117
rect 42379 300052 42380 300116
rect 42444 300052 42445 300116
rect 42379 300051 42445 300052
rect 41827 298484 41893 298485
rect 41827 298420 41828 298484
rect 41892 298420 41893 298484
rect 41827 298419 41893 298420
rect 41830 296850 41890 298419
rect 42195 297668 42261 297669
rect 42195 297604 42196 297668
rect 42260 297604 42261 297668
rect 42195 297603 42261 297604
rect 41462 296790 41890 296850
rect 41462 255101 41522 296790
rect 42011 295628 42077 295629
rect 42011 295564 42012 295628
rect 42076 295564 42077 295628
rect 42011 295563 42077 295564
rect 41827 295356 41893 295357
rect 41827 295292 41828 295356
rect 41892 295292 41893 295356
rect 41827 295291 41893 295292
rect 41643 289236 41709 289237
rect 41643 289172 41644 289236
rect 41708 289172 41709 289236
rect 41643 289171 41709 289172
rect 41646 256325 41706 289171
rect 41643 256324 41709 256325
rect 41643 256260 41644 256324
rect 41708 256260 41709 256324
rect 41643 256259 41709 256260
rect 41459 255100 41525 255101
rect 41459 255036 41460 255100
rect 41524 255036 41525 255100
rect 41459 255035 41525 255036
rect 41459 254284 41525 254285
rect 41459 254220 41460 254284
rect 41524 254220 41525 254284
rect 41459 254219 41525 254220
rect 41462 248826 41522 254219
rect 41830 254013 41890 295291
rect 42014 272373 42074 295563
rect 42198 295357 42258 297603
rect 42195 295356 42261 295357
rect 42195 295292 42196 295356
rect 42260 295292 42261 295356
rect 42195 295291 42261 295292
rect 42382 289237 42442 300051
rect 42379 289236 42445 289237
rect 42379 289172 42380 289236
rect 42444 289172 42445 289236
rect 42379 289171 42445 289172
rect 42379 285972 42445 285973
rect 42379 285908 42380 285972
rect 42444 285908 42445 285972
rect 42379 285907 42445 285908
rect 42195 285836 42261 285837
rect 42195 285772 42196 285836
rect 42260 285772 42261 285836
rect 42195 285771 42261 285772
rect 42011 272372 42077 272373
rect 42011 272308 42012 272372
rect 42076 272308 42077 272372
rect 42011 272307 42077 272308
rect 42198 269381 42258 285771
rect 42382 270061 42442 285907
rect 42563 285700 42629 285701
rect 42563 285636 42564 285700
rect 42628 285636 42629 285700
rect 42563 285635 42629 285636
rect 42566 270469 42626 285635
rect 44038 278493 44098 438910
rect 673686 438870 673746 489227
rect 674974 487661 675034 537682
rect 674971 487660 675037 487661
rect 674971 487596 674972 487660
rect 675036 487596 675037 487660
rect 674971 487595 675037 487596
rect 675158 484805 675218 537866
rect 675342 529005 675402 538050
rect 675526 531045 675586 538234
rect 675523 531044 675589 531045
rect 675523 530980 675524 531044
rect 675588 530980 675589 531044
rect 675523 530979 675589 530980
rect 675339 529004 675405 529005
rect 675339 528940 675340 529004
rect 675404 528940 675405 529004
rect 675339 528939 675405 528940
rect 675710 497193 675770 538418
rect 675894 497314 675954 538602
rect 676078 529413 676138 538786
rect 676075 529412 676141 529413
rect 676075 529348 676076 529412
rect 676140 529348 676141 529412
rect 676075 529347 676141 529348
rect 676262 527373 676322 538970
rect 676259 527372 676325 527373
rect 676259 527308 676260 527372
rect 676324 527308 676325 527372
rect 676259 527307 676325 527308
rect 676446 497467 676506 539406
rect 677187 539282 677247 541471
rect 676630 539222 677247 539282
rect 676630 497637 676690 539222
rect 677371 539098 677431 541655
rect 676814 539038 677431 539098
rect 676814 526965 676874 539038
rect 676811 526964 676877 526965
rect 676811 526900 676812 526964
rect 676876 526900 676877 526964
rect 676811 526899 676877 526900
rect 676630 497577 677168 497637
rect 676446 497407 677018 497467
rect 675894 497254 676885 497314
rect 675710 497133 676760 497193
rect 676700 495452 676760 497133
rect 675710 495392 676760 495452
rect 675710 486845 675770 495392
rect 676825 495233 676885 497254
rect 675894 495173 676885 495233
rect 675707 486844 675773 486845
rect 675707 486780 675708 486844
rect 675772 486780 675773 486844
rect 675707 486779 675773 486780
rect 675894 485213 675954 495173
rect 676958 495064 677018 497407
rect 676446 495004 677018 495064
rect 676446 492421 676506 495004
rect 677108 494922 677168 497577
rect 676630 494862 677168 494922
rect 676443 492420 676509 492421
rect 676443 492356 676444 492420
rect 676508 492356 676509 492420
rect 676443 492355 676509 492356
rect 675891 485212 675957 485213
rect 675891 485148 675892 485212
rect 675956 485148 675957 485212
rect 675891 485147 675957 485148
rect 675155 484804 675221 484805
rect 675155 484740 675156 484804
rect 675220 484740 675221 484804
rect 675155 484739 675221 484740
rect 676075 484532 676141 484533
rect 676075 484468 676076 484532
rect 676140 484530 676141 484532
rect 676630 484530 676690 494862
rect 676811 492420 676877 492421
rect 676811 492356 676812 492420
rect 676876 492356 676877 492420
rect 676811 492355 676877 492356
rect 676140 484470 676690 484530
rect 676140 484468 676141 484470
rect 676075 484467 676141 484468
rect 676814 483003 676874 492355
rect 676811 483002 676877 483003
rect 676811 482938 676812 483002
rect 676876 482938 676877 483002
rect 676811 482937 676877 482938
rect 673502 438810 673746 438870
rect 673502 279013 673562 438810
rect 673683 401028 673749 401029
rect 673683 400964 673684 401028
rect 673748 400964 673749 401028
rect 673683 400963 673749 400964
rect 673686 279693 673746 400963
rect 673867 400212 673933 400213
rect 673867 400148 673868 400212
rect 673932 400148 673933 400212
rect 673867 400147 673933 400148
rect 673683 279692 673749 279693
rect 673683 279628 673684 279692
rect 673748 279628 673749 279692
rect 673683 279627 673749 279628
rect 673870 279149 673930 400147
rect 674051 357508 674117 357509
rect 674051 357444 674052 357508
rect 674116 357444 674117 357508
rect 674051 357443 674117 357444
rect 674054 279557 674114 357443
rect 674235 355876 674301 355877
rect 674235 355812 674236 355876
rect 674300 355812 674301 355876
rect 674235 355811 674301 355812
rect 674051 279556 674117 279557
rect 674051 279492 674052 279556
rect 674116 279492 674117 279556
rect 674051 279491 674117 279492
rect 674238 279285 674298 355811
rect 674419 355060 674485 355061
rect 674419 354996 674420 355060
rect 674484 354996 674485 355060
rect 674419 354995 674485 354996
rect 674422 279421 674482 354995
rect 676075 353700 676141 353701
rect 676075 353636 676076 353700
rect 676140 353636 676141 353700
rect 676075 353635 676141 353636
rect 675891 352204 675957 352205
rect 675891 352140 675892 352204
rect 675956 352140 675957 352204
rect 675891 352139 675957 352140
rect 675707 350572 675773 350573
rect 675707 350508 675708 350572
rect 675772 350508 675773 350572
rect 675707 350507 675773 350508
rect 675710 330581 675770 350507
rect 675707 330580 675773 330581
rect 675707 330516 675708 330580
rect 675772 330516 675773 330580
rect 675707 330515 675773 330516
rect 675894 326909 675954 352139
rect 676078 328405 676138 353635
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 675891 326908 675957 326909
rect 675891 326844 675892 326908
rect 675956 326844 675957 326908
rect 675891 326843 675957 326844
rect 675891 305964 675957 305965
rect 675891 305900 675892 305964
rect 675956 305900 675957 305964
rect 675891 305899 675957 305900
rect 675894 291685 675954 305899
rect 675891 291684 675957 291685
rect 675891 291620 675892 291684
rect 675956 291620 675957 291684
rect 675891 291619 675957 291620
rect 674419 279420 674485 279421
rect 674419 279356 674420 279420
rect 674484 279356 674485 279420
rect 674419 279355 674485 279356
rect 674235 279284 674301 279285
rect 674235 279220 674236 279284
rect 674300 279220 674301 279284
rect 674235 279219 674301 279220
rect 673867 279148 673933 279149
rect 673867 279084 673868 279148
rect 673932 279084 673933 279148
rect 673867 279083 673933 279084
rect 673499 279012 673565 279013
rect 673499 278948 673500 279012
rect 673564 278948 673565 279012
rect 673499 278947 673565 278948
rect 44035 278492 44101 278493
rect 44035 278428 44036 278492
rect 44100 278428 44101 278492
rect 44035 278427 44101 278428
rect 42563 270468 42629 270469
rect 42563 270404 42564 270468
rect 42628 270404 42629 270468
rect 42563 270403 42629 270404
rect 42379 270060 42445 270061
rect 42379 269996 42380 270060
rect 42444 269996 42445 270060
rect 42379 269995 42445 269996
rect 42195 269380 42261 269381
rect 42195 269316 42196 269380
rect 42260 269316 42261 269380
rect 42195 269315 42261 269316
rect 674235 264620 674301 264621
rect 674235 264556 674236 264620
rect 674300 264556 674301 264620
rect 674235 264555 674301 264556
rect 674238 262445 674298 264555
rect 674235 262444 674301 262445
rect 674235 262380 674236 262444
rect 674300 262380 674301 262444
rect 674235 262379 674301 262380
rect 675891 262444 675957 262445
rect 675891 262380 675892 262444
rect 675956 262380 675957 262444
rect 675891 262379 675957 262380
rect 42195 256868 42261 256869
rect 42195 256804 42196 256868
rect 42260 256804 42261 256868
rect 42195 256803 42261 256804
rect 42011 255236 42077 255237
rect 42011 255172 42012 255236
rect 42076 255172 42077 255236
rect 42011 255171 42077 255172
rect 41827 254012 41893 254013
rect 41827 253948 41828 254012
rect 41892 253948 41893 254012
rect 41827 253947 41893 253948
rect 42014 253330 42074 255171
rect 40144 248766 41522 248826
rect 41830 253270 42074 253330
rect 40144 236980 40204 248766
rect 41830 248458 41890 253270
rect 42011 252788 42077 252789
rect 42011 252724 42012 252788
rect 42076 252724 42077 252788
rect 42011 252723 42077 252724
rect 40332 248398 41890 248458
rect 40332 237348 40392 248398
rect 42014 248274 42074 252723
rect 40516 248214 42074 248274
rect 40516 237532 40576 248214
rect 42198 248090 42258 256803
rect 675894 252400 675954 262379
rect 675894 252340 676888 252400
rect 40700 248030 42258 248090
rect 40700 237716 40760 248030
rect 675954 245610 676138 245670
rect 40700 237656 42258 237716
rect 40516 237472 42074 237532
rect 40332 237288 41890 237348
rect 40144 236920 41522 236980
rect 41462 211037 41522 236920
rect 41830 211717 41890 237288
rect 42014 225997 42074 237472
rect 42011 225996 42077 225997
rect 42011 225932 42012 225996
rect 42076 225932 42077 225996
rect 42011 225931 42077 225932
rect 42198 213349 42258 237656
rect 676078 228956 676138 245610
rect 676078 226654 676138 226658
rect 676828 226654 676888 252340
rect 676078 226594 676888 226654
rect 676078 220013 676138 226594
rect 676075 220012 676141 220013
rect 676075 219948 676076 220012
rect 676140 219948 676141 220012
rect 676075 219947 676141 219948
rect 42195 213348 42261 213349
rect 42195 213284 42196 213348
rect 42260 213284 42261 213348
rect 42195 213283 42261 213284
rect 41827 211716 41893 211717
rect 41827 211652 41828 211716
rect 41892 211652 41893 211716
rect 41827 211651 41893 211652
rect 41459 211036 41525 211037
rect 41459 210972 41460 211036
rect 41524 210972 41525 211036
rect 41459 210971 41525 210972
rect 42747 210492 42813 210493
rect 42747 210428 42748 210492
rect 42812 210428 42813 210492
rect 42747 210427 42813 210428
rect 41827 209676 41893 209677
rect 41827 209612 41828 209676
rect 41892 209612 41893 209676
rect 41827 209611 41893 209612
rect 41643 207772 41709 207773
rect 41643 207708 41644 207772
rect 41708 207708 41709 207772
rect 41643 207707 41709 207708
rect 41459 205732 41525 205733
rect 41459 205668 41460 205732
rect 41524 205668 41525 205732
rect 41459 205667 41525 205668
rect 41462 187645 41522 205667
rect 41459 187644 41525 187645
rect 41459 187580 41460 187644
rect 41524 187580 41525 187644
rect 41459 187579 41525 187580
rect 41646 183701 41706 207707
rect 41643 183700 41709 183701
rect 41643 183636 41644 183700
rect 41708 183636 41709 183700
rect 41643 183635 41709 183636
rect 41830 182749 41890 209611
rect 42379 209268 42445 209269
rect 42379 209204 42380 209268
rect 42444 209204 42445 209268
rect 42379 209203 42445 209204
rect 42011 207636 42077 207637
rect 42011 207572 42012 207636
rect 42076 207572 42077 207636
rect 42011 207571 42077 207572
rect 42014 186421 42074 207571
rect 42195 207228 42261 207229
rect 42195 207164 42196 207228
rect 42260 207164 42261 207228
rect 42195 207163 42261 207164
rect 42198 187101 42258 207163
rect 42195 187100 42261 187101
rect 42195 187036 42196 187100
rect 42260 187036 42261 187100
rect 42195 187035 42261 187036
rect 42011 186420 42077 186421
rect 42011 186356 42012 186420
rect 42076 186356 42077 186420
rect 42011 186355 42077 186356
rect 42382 185877 42442 209203
rect 42563 208860 42629 208861
rect 42563 208796 42564 208860
rect 42628 208796 42629 208860
rect 42563 208795 42629 208796
rect 42566 190229 42626 208795
rect 42563 190228 42629 190229
rect 42563 190164 42564 190228
rect 42628 190164 42629 190228
rect 42563 190163 42629 190164
rect 42379 185876 42445 185877
rect 42379 185812 42380 185876
rect 42444 185812 42445 185876
rect 42379 185811 42445 185812
rect 42750 184245 42810 210427
rect 42747 184244 42813 184245
rect 42747 184180 42748 184244
rect 42812 184180 42813 184244
rect 42747 184179 42813 184180
rect 41827 182748 41893 182749
rect 41827 182684 41828 182748
rect 41892 182684 41893 182748
rect 41827 182683 41893 182684
rect 675891 173636 675957 173637
rect 675891 173572 675892 173636
rect 675956 173572 675957 173636
rect 675891 173571 675957 173572
rect 675707 170780 675773 170781
rect 675707 170716 675708 170780
rect 675772 170716 675773 170780
rect 675707 170715 675773 170716
rect 675710 156501 675770 170715
rect 675707 156500 675773 156501
rect 675707 156436 675708 156500
rect 675772 156436 675773 156500
rect 675707 156435 675773 156436
rect 675894 148477 675954 173571
rect 676075 171868 676141 171869
rect 676075 171804 676076 171868
rect 676140 171804 676141 171868
rect 676075 171803 676141 171804
rect 675891 148476 675957 148477
rect 675891 148412 675892 148476
rect 675956 148412 675957 148476
rect 675891 148411 675957 148412
rect 676078 146301 676138 171803
rect 676075 146300 676141 146301
rect 676075 146236 676076 146300
rect 676140 146236 676141 146300
rect 676075 146235 676141 146236
rect 675891 128484 675957 128485
rect 675891 128420 675892 128484
rect 675956 128420 675957 128484
rect 675891 128419 675957 128420
rect 580947 113252 581013 113253
rect 580947 113188 580948 113252
rect 581012 113188 581013 113252
rect 580947 113187 581013 113188
rect 580950 73541 581010 113187
rect 675894 103325 675954 128419
rect 676075 126580 676141 126581
rect 676075 126516 676076 126580
rect 676140 126516 676141 126580
rect 676075 126515 676141 126516
rect 675891 103324 675957 103325
rect 675891 103260 675892 103324
rect 675956 103260 675957 103324
rect 675891 103259 675957 103260
rect 676078 101421 676138 126515
rect 676075 101420 676141 101421
rect 676075 101356 676076 101420
rect 676140 101356 676141 101420
rect 676075 101355 676141 101356
rect 662091 95572 662157 95573
rect 662091 95508 662092 95572
rect 662156 95508 662157 95572
rect 662091 95507 662157 95508
rect 662094 88773 662154 95507
rect 662091 88772 662157 88773
rect 662091 88708 662092 88772
rect 662156 88708 662157 88772
rect 662091 88707 662157 88708
rect 580947 73540 581013 73541
rect 580947 73476 580948 73540
rect 581012 73476 581013 73540
rect 580947 73475 581013 73476
rect 520411 48244 520477 48245
rect 520411 48180 520412 48244
rect 520476 48180 520477 48244
rect 520411 48179 520477 48180
rect 520414 42125 520474 48179
rect 520411 42124 520477 42125
rect 520411 42060 520412 42124
rect 520476 42060 520477 42124
rect 520411 42059 520477 42060
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
<< comment >>
rect 0 1037400 717600 1037600
rect 0 37510 200 1037400
rect 717400 200 717600 1037400
rect 39330 0 717600 200
use caravel_clocking  clocking
timestamp 1637509978
transform 1 0 205746 0 1 5488
box -38 -48 20000 12000
use xres_buf  rstb_level
timestamp 1637509978
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use caravel_logo  caravel_logo_0
timestamp 1636495793
transform 1 0 324236 0 1 5094
box -2520 0 15000 15560
use open_source  open_source_0 hexdigits
timestamp 1635801696
transform 1 0 260430 0 1 2174
box 752 5164 29030 16242
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use copyright_block  copyright_block_0
timestamp 1636248654
transform 1 0 149582 0 1 16298
box -262 -9464 35048 2764
use simple_por  por
timestamp 1637509978
transform 1 0 650146 0 -1 55282
box 0 0 11344 8338
use gpio_defaults_block  gpio_01_defaults\[0\]
timestamp 1637509978
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1637509978
transform -1 0 710203 0 1 121000
box 882 167 34000 13000
use housekeeping  housekeeping
timestamp 1637509978
transform 1 0 606434 0 1 100002
box 0 0 60046 110190
use digital_pll  pll
timestamp 1637509978
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use user_id_programming  user_id_value
timestamp 1637509978
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1637416673
transform 1 0 52034 0 1 53002
box 382 -400 524400 164400
use gpio_defaults_block  gpio_37_defaults
timestamp 1637509978
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1637509978
transform 1 0 7631 0 1 202600
box 882 167 34000 13000
use gpio_defaults_block  gpio_01_defaults\[1\]
timestamp 1637509978
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1637509978
transform -1 0 710203 0 1 166200
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1637509978
transform -1 0 710203 0 1 211200
box 882 167 34000 13000
use gpio_defaults_block  gpio_36_defaults
timestamp 1637509978
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1637509978
transform 1 0 7631 0 1 245800
box 882 167 34000 13000
use mgmt_protect  mgmt_buffers
timestamp 1637509978
transform 1 0 192180 0 1 232036
box -400 -400 220400 32400
use gpio_defaults_block  gpio_234_defaults\[1\]
timestamp 1637509978
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_234_defaults\[0\]
timestamp 1637509978
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1637509978
transform -1 0 710203 0 1 256400
box 882 167 34000 13000
use gpio_defaults_block  gpio_35_defaults
timestamp 1637509978
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1637509978
transform 1 0 7631 0 1 289000
box 882 167 34000 13000
use gpio_defaults_block  gpio_234_defaults\[2\]
timestamp 1637509978
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1637509978
transform -1 0 710203 0 1 301400
box 882 167 34000 13000
use gpio_defaults_block  gpio_32_defaults
timestamp 1637509978
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_33_defaults
timestamp 1637509978
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_34_defaults
timestamp 1637509978
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1637509978
transform 1 0 7631 0 1 418600
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1637509978
transform 1 0 7631 0 1 375400
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1637509978
transform 1 0 7631 0 1 332200
box 882 167 34000 13000
use gpio_defaults_block  gpio_6_defaults
timestamp 1637509978
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_5_defaults
timestamp 1637509978
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_7_defaults
timestamp 1637509978
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1637509978
transform -1 0 710203 0 1 346400
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1637509978
transform -1 0 710203 0 1 391600
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1637509978
transform -1 0 710203 0 1 479800
box 882 167 34000 13000
use gpio_defaults_block  gpio_30_defaults
timestamp 1637509978
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_defaults_block  gpio_31_defaults
timestamp 1637509978
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1637509978
transform 1 0 7631 0 1 589400
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1637509978
transform 1 0 7631 0 1 546200
box 882 167 34000 13000
use gpio_defaults_block  gpio_9_defaults
timestamp 1637509978
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_8_defaults
timestamp 1637509978
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1637509978
transform -1 0 710203 0 1 523800
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1637509978
transform -1 0 710203 0 1 568800
box 882 167 34000 13000
use gpio_defaults_block  gpio_28_defaults
timestamp 1637509978
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_29_defaults
timestamp 1637509978
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1637509978
transform 1 0 7631 0 1 632600
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1637509978
transform 1 0 7631 0 1 675800
box 882 167 34000 13000
use gpio_defaults_block  gpio_11_defaults
timestamp 1637509978
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_10_defaults
timestamp 1637509978
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1637509978
transform -1 0 710203 0 1 614000
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1637509978
transform -1 0 710203 0 1 659000
box 882 167 34000 13000
use gpio_defaults_block  gpio_26_defaults
timestamp 1637509978
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_27_defaults
timestamp 1637509978
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1637509978
transform 1 0 7631 0 1 762200
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1637509978
transform 1 0 7631 0 1 719000
box 882 167 34000 13000
use gpio_defaults_block  gpio_13_defaults
timestamp 1637509978
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_12_defaults
timestamp 1637509978
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1637509978
transform -1 0 710203 0 1 704200
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1637509978
transform -1 0 710203 0 1 749200
box 882 167 34000 13000
use gpio_defaults_block  gpio_25_defaults
timestamp 1637509978
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1637509978
transform 1 0 7631 0 1 805400
box 882 167 34000 13000
use gpio_defaults_block  gpio_24_defaults
timestamp 1637509978
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1637509978
transform 1 0 7631 0 1 931200
box 882 167 34000 13000
use gpio_defaults_block  gpio_14_defaults
timestamp 1637509978
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1637509978
transform -1 0 710203 0 1 927600
box 882 167 34000 13000
use gpio_defaults_block  gpio_22_defaults
timestamp 1637509978
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_23_defaults
timestamp 1637509978
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1637509978
transform 0 1 148600 -1 0 1030077
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1637509978
transform 0 1 97200 -1 0 1030077
box 882 167 34000 13000
use gpio_defaults_block  gpio_21_defaults
timestamp 1637509978
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1637509978
transform 0 1 251400 -1 0 1030077
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1637509978
transform 0 1 200000 -1 0 1030077
box 882 167 34000 13000
use gpio_defaults_block  gpio_19_defaults
timestamp 1637509978
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_20_defaults
timestamp 1637509978
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1637509978
transform 0 1 303000 -1 0 1030077
box 882 167 34000 13000
use gpio_defaults_block  gpio_17_defaults
timestamp 1637509978
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_18_defaults
timestamp 1637509978
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1637509978
transform 0 1 353400 -1 0 1030077
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1637509978
transform 0 1 420800 -1 0 1030077
box 882 167 34000 13000
use gpio_defaults_block  gpio_16_defaults
timestamp 1637509978
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1637509978
transform 0 1 497800 -1 0 1030077
box 882 167 34000 13000
use gpio_defaults_block  gpio_15_defaults
timestamp 1637509978
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1637509978
transform 0 1 549200 -1 0 1030077
box 882 167 34000 13000
use user_project_wrapper  mprj
timestamp 1637147503
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1637509978
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use caravel_power_routing  caravel_power_routing_0
timestamp 1637516397
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 24000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 24000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 24000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 24000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 24000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 24000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 24000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 24000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 24000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 24000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 24000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698512 952840 711002 965360 0 FreeSans 24000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628240 1018512 640760 1031002 0 FreeSans 24000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526440 1018512 538960 1031002 0 FreeSans 24000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475040 1018512 487560 1031002 0 FreeSans 24000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386040 1018512 398560 1031002 0 FreeSans 24000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284240 1018512 296760 1031002 0 FreeSans 24000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 24000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 232640 1018512 245160 1031002 0 FreeSans 24000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181240 1018512 193760 1031002 0 FreeSans 24000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 129840 1018512 142360 1031002 0 FreeSans 24000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78440 1018512 90960 1031002 0 FreeSans 24000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6598 956440 19088 968960 0 FreeSans 24000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 24000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 24000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 24000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 24000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 24000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 24000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 24000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 24000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 24000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 24000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 24000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 24000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 24000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 24000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 24000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 24000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 24000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 24000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 24000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 24000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 24000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144150 18309 0 FreeSans 24000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 24000 0 0 0 vccd
port 45 nsew signal bidirectional
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 24000 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 24000 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 24000 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 24000 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 24000 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 24000 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 24000 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 24000 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 24000 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 24000 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 24000 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 24000 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 24000 0 0 0 vssd
port 58 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 24000 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 24000 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 24000 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 24000 0 0 0 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
