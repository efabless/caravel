magic
tech sky130A
magscale 1 2
timestamp 1636035201
<< locali >>
rect 9873 11067 9907 11305
rect 7297 8891 7331 9061
rect 3065 7735 3099 7905
rect 3433 7803 3467 7905
rect 2789 7191 2823 7293
rect 2697 2839 2731 6409
rect 2789 3179 2823 5729
rect 2881 4471 2915 5185
<< viali >>
rect 1685 11305 1719 11339
rect 2237 11305 2271 11339
rect 2421 11305 2455 11339
rect 4077 11305 4111 11339
rect 4445 11305 4479 11339
rect 4813 11305 4847 11339
rect 5181 11305 5215 11339
rect 7849 11305 7883 11339
rect 9873 11305 9907 11339
rect 2697 11237 2731 11271
rect 9045 11237 9079 11271
rect 9413 11237 9447 11271
rect 1869 11101 1903 11135
rect 2605 11101 2639 11135
rect 2881 11101 2915 11135
rect 3157 11101 3191 11135
rect 3433 11101 3467 11135
rect 3617 11101 3651 11135
rect 3893 11101 3927 11135
rect 4261 11101 4295 11135
rect 4629 11101 4663 11135
rect 4997 11101 5031 11135
rect 5733 11101 5767 11135
rect 6193 11101 6227 11135
rect 6561 11101 6595 11135
rect 6929 11101 6963 11135
rect 7297 11101 7331 11135
rect 7665 11101 7699 11135
rect 8309 11101 8343 11135
rect 8861 11101 8895 11135
rect 9229 11101 9263 11135
rect 5457 11033 5491 11067
rect 5641 11033 5675 11067
rect 9873 11033 9907 11067
rect 1501 10965 1535 10999
rect 2973 10965 3007 10999
rect 3249 10965 3283 10999
rect 3709 10965 3743 10999
rect 5917 10965 5951 10999
rect 6377 10965 6411 10999
rect 6745 10965 6779 10999
rect 7113 10965 7147 10999
rect 7481 10965 7515 10999
rect 8493 10965 8527 10999
rect 1225 10761 1259 10795
rect 2053 10761 2087 10795
rect 2145 10761 2179 10795
rect 8677 10761 8711 10795
rect 9045 10693 9079 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 2329 10625 2363 10659
rect 4250 10625 4284 10659
rect 6285 10625 6319 10659
rect 8125 10625 8159 10659
rect 2421 10557 2455 10591
rect 2697 10557 2731 10591
rect 4537 10557 4571 10591
rect 6653 10557 6687 10591
rect 9137 10557 9171 10591
rect 9229 10557 9263 10591
rect 1501 10489 1535 10523
rect 8585 10489 8619 10523
rect 4169 10421 4203 10455
rect 6009 10421 6043 10455
rect 1777 10217 1811 10251
rect 2145 10217 2179 10251
rect 2697 10217 2731 10251
rect 7389 10217 7423 10251
rect 7573 10217 7607 10251
rect 8769 10217 8803 10251
rect 2421 10149 2455 10183
rect 2973 10149 3007 10183
rect 4261 10149 4295 10183
rect 6929 10149 6963 10183
rect 4629 10081 4663 10115
rect 8401 10081 8435 10115
rect 9321 10081 9355 10115
rect 2053 10013 2087 10047
rect 2329 10013 2363 10047
rect 2605 10013 2639 10047
rect 2881 10013 2915 10047
rect 3157 10013 3191 10047
rect 3433 10013 3467 10047
rect 3893 10013 3927 10047
rect 4169 10013 4203 10047
rect 4445 10013 4479 10047
rect 4997 10013 5031 10047
rect 6469 10013 6503 10047
rect 7481 10013 7515 10047
rect 9137 10013 9171 10047
rect 7021 9945 7055 9979
rect 7205 9945 7239 9979
rect 8033 9945 8067 9979
rect 8217 9945 8251 9979
rect 9229 9945 9263 9979
rect 1869 9877 1903 9911
rect 3249 9877 3283 9911
rect 3709 9877 3743 9911
rect 3985 9877 4019 9911
rect 7941 9877 7975 9911
rect 2421 9673 2455 9707
rect 6653 9673 6687 9707
rect 2329 9605 2363 9639
rect 8033 9605 8067 9639
rect 2605 9537 2639 9571
rect 2697 9537 2731 9571
rect 2789 9537 2823 9571
rect 3341 9537 3375 9571
rect 3617 9537 3651 9571
rect 4077 9537 4111 9571
rect 5549 9537 5583 9571
rect 6193 9537 6227 9571
rect 6745 9537 6779 9571
rect 6929 9537 6963 9571
rect 7389 9537 7423 9571
rect 8217 9537 8251 9571
rect 3709 9469 3743 9503
rect 6009 9469 6043 9503
rect 7481 9469 7515 9503
rect 8585 9469 8619 9503
rect 3157 9401 3191 9435
rect 7941 9401 7975 9435
rect 3433 9333 3467 9367
rect 6285 9333 6319 9367
rect 7113 9333 7147 9367
rect 7205 9333 7239 9367
rect 1777 9129 1811 9163
rect 2973 9129 3007 9163
rect 5365 9129 5399 9163
rect 8585 9129 8619 9163
rect 2697 9061 2731 9095
rect 7297 9061 7331 9095
rect 7665 9061 7699 9095
rect 3617 8993 3651 9027
rect 5733 8993 5767 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 1961 8925 1995 8959
rect 2329 8925 2363 8959
rect 2605 8925 2639 8959
rect 2881 8925 2915 8959
rect 3157 8925 3191 8959
rect 3433 8925 3467 8959
rect 5457 8925 5491 8959
rect 7481 8925 7515 8959
rect 8125 8925 8159 8959
rect 8217 8925 8251 8959
rect 8401 8925 8435 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 3893 8857 3927 8891
rect 7297 8857 7331 8891
rect 8769 8857 8803 8891
rect 1225 8789 1259 8823
rect 1501 8789 1535 8823
rect 2421 8789 2455 8823
rect 3249 8789 3283 8823
rect 7205 8789 7239 8823
rect 9137 8789 9171 8823
rect 9413 8789 9447 8823
rect 4353 8585 4387 8619
rect 4675 8585 4709 8619
rect 5825 8585 5859 8619
rect 6193 8585 6227 8619
rect 9505 8585 9539 8619
rect 2237 8517 2271 8551
rect 2881 8517 2915 8551
rect 1593 8449 1627 8483
rect 1869 8449 1903 8483
rect 2513 8473 2547 8507
rect 5365 8449 5399 8483
rect 6377 8449 6411 8483
rect 6469 8449 6503 8483
rect 9045 8449 9079 8483
rect 2605 8381 2639 8415
rect 4445 8381 4479 8415
rect 7205 8381 7239 8415
rect 7573 8381 7607 8415
rect 1409 8313 1443 8347
rect 2329 8313 2363 8347
rect 7113 8313 7147 8347
rect 1685 8245 1719 8279
rect 5457 8245 5491 8279
rect 1685 8041 1719 8075
rect 3709 8041 3743 8075
rect 6469 8041 6503 8075
rect 8401 8041 8435 8075
rect 8861 8041 8895 8075
rect 9321 8041 9355 8075
rect 1409 7973 1443 8007
rect 2237 7973 2271 8007
rect 4261 7973 4295 8007
rect 8309 7973 8343 8007
rect 3065 7905 3099 7939
rect 1593 7837 1627 7871
rect 1869 7837 1903 7871
rect 2145 7837 2179 7871
rect 2421 7837 2455 7871
rect 2697 7837 2731 7871
rect 2981 7833 3015 7867
rect 3433 7905 3467 7939
rect 4997 7905 5031 7939
rect 6561 7905 6595 7939
rect 6837 7905 6871 7939
rect 9229 7905 9263 7939
rect 4721 7837 4755 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 9505 7837 9539 7871
rect 3433 7769 3467 7803
rect 3801 7769 3835 7803
rect 3985 7769 4019 7803
rect 1961 7701 1995 7735
rect 2513 7701 2547 7735
rect 2789 7701 2823 7735
rect 3065 7701 3099 7735
rect 3341 7701 3375 7735
rect 4445 7701 4479 7735
rect 3249 7497 3283 7531
rect 8493 7497 8527 7531
rect 9321 7497 9355 7531
rect 3065 7429 3099 7463
rect 1501 7361 1535 7395
rect 1777 7361 1811 7395
rect 2053 7361 2087 7395
rect 2329 7361 2363 7395
rect 2697 7361 2731 7395
rect 3433 7361 3467 7395
rect 3893 7361 3927 7395
rect 4077 7361 4111 7395
rect 6561 7361 6595 7395
rect 8033 7361 8067 7395
rect 8769 7361 8803 7395
rect 9505 7361 9539 7395
rect 2789 7293 2823 7327
rect 4353 7293 4387 7327
rect 6193 7293 6227 7327
rect 1593 7225 1627 7259
rect 3801 7225 3835 7259
rect 5825 7225 5859 7259
rect 9229 7225 9263 7259
rect 1317 7157 1351 7191
rect 1869 7157 1903 7191
rect 2145 7157 2179 7191
rect 2513 7157 2547 7191
rect 2789 7157 2823 7191
rect 3617 7157 3651 7191
rect 9045 7157 9079 7191
rect 8125 6953 8159 6987
rect 1685 6817 1719 6851
rect 5917 6817 5951 6851
rect 9321 6817 9355 6851
rect 1593 6749 1627 6783
rect 3617 6749 3651 6783
rect 3985 6749 4019 6783
rect 5457 6749 5491 6783
rect 8033 6749 8067 6783
rect 9137 6749 9171 6783
rect 1317 6681 1351 6715
rect 1961 6681 1995 6715
rect 6193 6681 6227 6715
rect 1409 6613 1443 6647
rect 3433 6613 3467 6647
rect 7481 6613 7515 6647
rect 8493 6613 8527 6647
rect 8769 6613 8803 6647
rect 9229 6613 9263 6647
rect 2697 6409 2731 6443
rect 8677 6409 8711 6443
rect 9137 6409 9171 6443
rect 3433 6341 3467 6375
rect 3617 6341 3651 6375
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 4169 6273 4203 6307
rect 4537 6273 4571 6307
rect 6009 6273 6043 6307
rect 7481 6273 7515 6307
rect 8309 6273 8343 6307
rect 9045 6273 9079 6307
rect 6561 6205 6595 6239
rect 6837 6205 6871 6239
rect 9321 6205 9355 6239
rect 4077 6137 4111 6171
rect 6469 6137 6503 6171
rect 8493 6137 8527 6171
rect 7757 6069 7791 6103
rect 7941 6069 7975 6103
rect 3604 5865 3638 5899
rect 5825 5865 5859 5899
rect 6285 5865 6319 5899
rect 8677 5865 8711 5899
rect 8953 5865 8987 5899
rect 2789 5729 2823 5763
rect 3341 5729 3375 5763
rect 6193 5729 6227 5763
rect 7021 5729 7055 5763
rect 5181 5661 5215 5695
rect 5365 5661 5399 5695
rect 5733 5661 5767 5695
rect 6469 5661 6503 5695
rect 6653 5661 6687 5695
rect 8493 5661 8527 5695
rect 9045 5661 9079 5695
rect 5549 5593 5583 5627
rect 9229 5593 9263 5627
rect 5089 5525 5123 5559
rect 9413 5525 9447 5559
rect 3341 5321 3375 5355
rect 9137 5253 9171 5287
rect 9321 5253 9355 5287
rect 2881 5185 2915 5219
rect 3525 5185 3559 5219
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 6193 5185 6227 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 8677 5185 8711 5219
rect 8861 5185 8895 5219
rect 4261 5117 4295 5151
rect 5733 5117 5767 5151
rect 5825 5117 5859 5151
rect 8493 5049 8527 5083
rect 3617 4981 3651 5015
rect 8125 4981 8159 5015
rect 9045 4981 9079 5015
rect 9505 4981 9539 5015
rect 5549 4777 5583 4811
rect 5825 4777 5859 4811
rect 6285 4777 6319 4811
rect 9505 4777 9539 4811
rect 3433 4709 3467 4743
rect 6193 4709 6227 4743
rect 6653 4709 6687 4743
rect 6929 4709 6963 4743
rect 3525 4641 3559 4675
rect 4077 4641 4111 4675
rect 7205 4641 7239 4675
rect 3709 4573 3743 4607
rect 3801 4573 3835 4607
rect 5733 4573 5767 4607
rect 6469 4573 6503 4607
rect 6837 4573 6871 4607
rect 7113 4573 7147 4607
rect 7573 4573 7607 4607
rect 9045 4573 9079 4607
rect 2881 4437 2915 4471
rect 7573 4233 7607 4267
rect 9321 4233 9355 4267
rect 3709 4097 3743 4131
rect 3985 4097 4019 4131
rect 4353 4097 4387 4131
rect 4813 4097 4847 4131
rect 6285 4097 6319 4131
rect 7205 4097 7239 4131
rect 7481 4097 7515 4131
rect 7757 4097 7791 4131
rect 7849 4097 7883 4131
rect 8309 4097 8343 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 9505 4097 9539 4131
rect 4445 4029 4479 4063
rect 8769 4029 8803 4063
rect 9229 4029 9263 4063
rect 3801 3961 3835 3995
rect 4169 3961 4203 3995
rect 7021 3961 7055 3995
rect 7297 3961 7331 3995
rect 8033 3961 8067 3995
rect 3525 3893 3559 3927
rect 6745 3893 6779 3927
rect 8585 3893 8619 3927
rect 5181 3689 5215 3723
rect 5365 3689 5399 3723
rect 8677 3689 8711 3723
rect 8861 3621 8895 3655
rect 3433 3553 3467 3587
rect 3709 3553 3743 3587
rect 6101 3553 6135 3587
rect 9321 3553 9355 3587
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 7573 3485 7607 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 9137 3417 9171 3451
rect 8033 3349 8067 3383
rect 8125 3349 8159 3383
rect 2789 3145 2823 3179
rect 6377 3145 6411 3179
rect 6469 3145 6503 3179
rect 7389 3145 7423 3179
rect 8309 3145 8343 3179
rect 3893 3009 3927 3043
rect 5365 3009 5399 3043
rect 5917 3009 5951 3043
rect 6653 3009 6687 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 7665 3009 7699 3043
rect 8493 3009 8527 3043
rect 3525 2941 3559 2975
rect 5825 2941 5859 2975
rect 8677 2941 8711 2975
rect 8861 2941 8895 2975
rect 7297 2873 7331 2907
rect 2697 2805 2731 2839
rect 6009 2805 6043 2839
rect 6929 2805 6963 2839
rect 7757 2805 7791 2839
rect 8125 2805 8159 2839
rect 9321 2805 9355 2839
rect 3341 2601 3375 2635
rect 3617 2601 3651 2635
rect 4353 2601 4387 2635
rect 6469 2601 6503 2635
rect 6745 2601 6779 2635
rect 7481 2601 7515 2635
rect 8309 2601 8343 2635
rect 9137 2601 9171 2635
rect 5273 2533 5307 2567
rect 6285 2533 6319 2567
rect 4629 2465 4663 2499
rect 3525 2397 3559 2431
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 4169 2397 4203 2431
rect 5457 2397 5491 2431
rect 5917 2397 5951 2431
rect 6653 2397 6687 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 7665 2397 7699 2431
rect 7941 2397 7975 2431
rect 8493 2397 8527 2431
rect 8769 2397 8803 2431
rect 9045 2397 9079 2431
rect 9321 2397 9355 2431
rect 4721 2329 4755 2363
rect 4905 2329 4939 2363
rect 6101 2329 6135 2363
rect 7021 2329 7055 2363
rect 7389 2329 7423 2363
rect 3893 2261 3927 2295
rect 5089 2261 5123 2295
rect 7757 2261 7791 2295
rect 8585 2261 8619 2295
rect 8861 2261 8895 2295
<< metal1 >>
rect 1854 11908 1860 11960
rect 1912 11948 1918 11960
rect 8110 11948 8116 11960
rect 1912 11920 8116 11948
rect 1912 11908 1918 11920
rect 8110 11908 8116 11920
rect 8168 11908 8174 11960
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 6638 11880 6644 11892
rect 2464 11852 6644 11880
rect 2464 11840 2470 11852
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 3142 11772 3148 11824
rect 3200 11812 3206 11824
rect 4062 11812 4068 11824
rect 3200 11784 4068 11812
rect 3200 11772 3206 11784
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 7374 11704 7380 11756
rect 7432 11744 7438 11756
rect 9490 11744 9496 11756
rect 7432 11716 9496 11744
rect 7432 11704 7438 11716
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 4338 11676 4344 11688
rect 2188 11648 4344 11676
rect 2188 11636 2194 11648
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 6730 11676 6736 11688
rect 6104 11648 6736 11676
rect 2314 11568 2320 11620
rect 2372 11608 2378 11620
rect 3602 11608 3608 11620
rect 2372 11580 3608 11608
rect 2372 11568 2378 11580
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 3694 11568 3700 11620
rect 3752 11608 3758 11620
rect 6104 11608 6132 11648
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 9766 11676 9772 11688
rect 7524 11648 9772 11676
rect 7524 11636 7530 11648
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 3752 11580 6132 11608
rect 3752 11568 3758 11580
rect 6178 11568 6184 11620
rect 6236 11608 6242 11620
rect 7650 11608 7656 11620
rect 6236 11580 7656 11608
rect 6236 11568 6242 11580
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 6822 11540 6828 11552
rect 3016 11512 6828 11540
rect 3016 11500 3022 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 13354 11540 13360 11552
rect 7616 11512 13360 11540
rect 7616 11500 7622 11512
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 5666 11450
rect 5718 11398 5730 11450
rect 5782 11398 5794 11450
rect 5846 11398 5858 11450
rect 5910 11398 5922 11450
rect 5974 11398 8766 11450
rect 8818 11398 8830 11450
rect 8882 11398 8894 11450
rect 8946 11398 8958 11450
rect 9010 11398 9022 11450
rect 9074 11398 9844 11450
rect 920 11376 9844 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2222 11336 2228 11348
rect 2183 11308 2228 11336
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2958 11336 2964 11348
rect 2455 11308 2964 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 4028 11308 4077 11336
rect 4028 11296 4034 11308
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 4614 11336 4620 11348
rect 4479 11308 4620 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 4798 11336 4804 11348
rect 4759 11308 4804 11336
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 5169 11339 5227 11345
rect 5169 11305 5181 11339
rect 5215 11336 5227 11339
rect 7006 11336 7012 11348
rect 5215 11308 7012 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 7742 11336 7748 11348
rect 7340 11308 7748 11336
rect 7340 11296 7346 11308
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 7837 11339 7895 11345
rect 7837 11305 7849 11339
rect 7883 11336 7895 11339
rect 9861 11339 9919 11345
rect 7883 11308 9352 11336
rect 7883 11305 7895 11308
rect 7837 11299 7895 11305
rect 2685 11271 2743 11277
rect 2685 11237 2697 11271
rect 2731 11237 2743 11271
rect 2685 11231 2743 11237
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 2222 11132 2228 11144
rect 1903 11104 2228 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2406 11092 2412 11144
rect 2464 11132 2470 11144
rect 2593 11135 2651 11141
rect 2593 11132 2605 11135
rect 2464 11104 2605 11132
rect 2464 11092 2470 11104
rect 2593 11101 2605 11104
rect 2639 11101 2651 11135
rect 2700 11132 2728 11231
rect 2774 11228 2780 11280
rect 2832 11268 2838 11280
rect 9033 11271 9091 11277
rect 9033 11268 9045 11271
rect 2832 11240 9045 11268
rect 2832 11228 2838 11240
rect 9033 11237 9045 11240
rect 9079 11237 9091 11271
rect 9033 11231 9091 11237
rect 5626 11200 5632 11212
rect 3068 11172 5632 11200
rect 2869 11135 2927 11141
rect 2700 11104 2820 11132
rect 2593 11095 2651 11101
rect 2792 11064 2820 11104
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 2958 11132 2964 11144
rect 2915 11104 2964 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3068 11064 3096 11172
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 6822 11200 6828 11212
rect 5736 11172 6828 11200
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11126 3203 11135
rect 3234 11126 3240 11144
rect 3191 11101 3240 11126
rect 3145 11098 3240 11101
rect 3145 11095 3203 11098
rect 3234 11092 3240 11098
rect 3292 11092 3298 11144
rect 3418 11132 3424 11144
rect 3379 11104 3424 11132
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3602 11132 3608 11144
rect 3563 11104 3608 11132
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 3881 11135 3939 11141
rect 3881 11132 3893 11135
rect 3752 11104 3893 11132
rect 3752 11092 3758 11104
rect 3881 11101 3893 11104
rect 3927 11101 3939 11135
rect 3881 11095 3939 11101
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4249 11135 4307 11141
rect 4249 11132 4261 11135
rect 4120 11104 4261 11132
rect 4120 11092 4126 11104
rect 4249 11101 4261 11104
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4396 11104 4629 11132
rect 4396 11092 4402 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4764 11104 4997 11132
rect 4764 11092 4770 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 5534 11132 5540 11144
rect 4985 11095 5043 11101
rect 5092 11104 5540 11132
rect 5092 11064 5120 11104
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 5736 11141 5764 11172
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 7098 11200 7104 11212
rect 6932 11172 7104 11200
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5994 11092 6000 11144
rect 6052 11132 6058 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 6052 11104 6193 11132
rect 6052 11092 6058 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 6932 11141 6960 11172
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7190 11160 7196 11212
rect 7248 11200 7254 11212
rect 9324 11200 9352 11308
rect 9861 11305 9873 11339
rect 9907 11336 9919 11339
rect 13722 11336 13728 11348
rect 9907 11308 13728 11336
rect 9907 11305 9919 11308
rect 9861 11299 9919 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 9401 11271 9459 11277
rect 9401 11237 9413 11271
rect 9447 11268 9459 11271
rect 13814 11268 13820 11280
rect 9447 11240 13820 11268
rect 9447 11237 9459 11240
rect 9401 11231 9459 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 13446 11200 13452 11212
rect 7248 11172 8156 11200
rect 9324 11172 13452 11200
rect 7248 11160 7254 11172
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 6512 11104 6561 11132
rect 6512 11092 6518 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11101 6975 11135
rect 7282 11132 7288 11144
rect 7243 11104 7288 11132
rect 6917 11095 6975 11101
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 7466 11132 7472 11144
rect 7392 11104 7472 11132
rect 2792 11036 3096 11064
rect 3252 11036 5120 11064
rect 1489 10999 1547 11005
rect 1489 10965 1501 10999
rect 1535 10996 1547 10999
rect 2590 10996 2596 11008
rect 1535 10968 2596 10996
rect 1535 10965 1547 10968
rect 1489 10959 1547 10965
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 2958 10996 2964 11008
rect 2919 10968 2964 10996
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 3252 11005 3280 11036
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 5445 11067 5503 11073
rect 5445 11064 5457 11067
rect 5316 11036 5457 11064
rect 5316 11024 5322 11036
rect 5445 11033 5457 11036
rect 5491 11033 5503 11067
rect 5445 11027 5503 11033
rect 5629 11067 5687 11073
rect 5629 11033 5641 11067
rect 5675 11064 5687 11067
rect 6270 11064 6276 11076
rect 5675 11036 6276 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 3237 10999 3295 11005
rect 3237 10965 3249 10999
rect 3283 10965 3295 10999
rect 3237 10959 3295 10965
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 3697 10999 3755 11005
rect 3697 10996 3709 10999
rect 3384 10968 3709 10996
rect 3384 10956 3390 10968
rect 3697 10965 3709 10968
rect 3743 10965 3755 10999
rect 3697 10959 3755 10965
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 5074 10996 5080 11008
rect 4028 10968 5080 10996
rect 4028 10956 4034 10968
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5166 10956 5172 11008
rect 5224 10996 5230 11008
rect 5644 10996 5672 11027
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 7190 11064 7196 11076
rect 6748 11036 7196 11064
rect 5224 10968 5672 10996
rect 5905 10999 5963 11005
rect 5224 10956 5230 10968
rect 5905 10965 5917 10999
rect 5951 10996 5963 10999
rect 6086 10996 6092 11008
rect 5951 10968 6092 10996
rect 5951 10965 5963 10968
rect 5905 10959 5963 10965
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 6362 10996 6368 11008
rect 6323 10968 6368 10996
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 6748 11005 6776 11036
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 6733 10999 6791 11005
rect 6733 10965 6745 10999
rect 6779 10965 6791 10999
rect 6733 10959 6791 10965
rect 7101 10999 7159 11005
rect 7101 10965 7113 10999
rect 7147 10996 7159 10999
rect 7392 10996 7420 11104
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 7650 11132 7656 11144
rect 7611 11104 7656 11132
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 8128 11064 8156 11172
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 8294 11132 8300 11144
rect 8255 11104 8300 11132
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 8849 11135 8907 11141
rect 8849 11132 8861 11135
rect 8444 11104 8861 11132
rect 8444 11092 8450 11104
rect 8849 11101 8861 11104
rect 8895 11101 8907 11135
rect 9214 11132 9220 11144
rect 9175 11104 9220 11132
rect 8849 11095 8907 11101
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 8128 11036 9873 11064
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 9861 11027 9919 11033
rect 7147 10968 7420 10996
rect 7469 10999 7527 11005
rect 7147 10965 7159 10968
rect 7101 10959 7159 10965
rect 7469 10965 7481 10999
rect 7515 10996 7527 10999
rect 7558 10996 7564 11008
rect 7515 10968 7564 10996
rect 7515 10965 7527 10968
rect 7469 10959 7527 10965
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 8478 10996 8484 11008
rect 8439 10968 8484 10996
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 16666 10996 16672 11008
rect 8628 10968 16672 10996
rect 8628 10956 8634 10968
rect 16666 10956 16672 10968
rect 16724 10956 16730 11008
rect 920 10906 9844 10928
rect 920 10854 4116 10906
rect 4168 10854 4180 10906
rect 4232 10854 4244 10906
rect 4296 10854 4308 10906
rect 4360 10854 4372 10906
rect 4424 10854 7216 10906
rect 7268 10854 7280 10906
rect 7332 10854 7344 10906
rect 7396 10854 7408 10906
rect 7460 10854 7472 10906
rect 7524 10854 9844 10906
rect 920 10832 9844 10854
rect 1210 10792 1216 10804
rect 1171 10764 1216 10792
rect 1210 10752 1216 10764
rect 1268 10752 1274 10804
rect 2038 10792 2044 10804
rect 1999 10764 2044 10792
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 3970 10792 3976 10804
rect 2179 10764 3976 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 5166 10792 5172 10804
rect 4172 10764 5172 10792
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2056 10656 2084 10752
rect 2682 10724 2688 10736
rect 2332 10696 2688 10724
rect 2332 10665 2360 10696
rect 2682 10684 2688 10696
rect 2740 10684 2746 10736
rect 3418 10684 3424 10736
rect 3476 10730 3482 10736
rect 3476 10724 3924 10730
rect 4062 10724 4068 10736
rect 3476 10702 4068 10724
rect 3476 10684 3482 10702
rect 3910 10696 4068 10702
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 1719 10628 2084 10656
rect 2317 10659 2375 10665
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 4172 10656 4200 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 8665 10795 8723 10801
rect 5828 10764 7880 10792
rect 4430 10684 4436 10736
rect 4488 10724 4494 10736
rect 4798 10724 4804 10736
rect 4488 10696 4804 10724
rect 4488 10684 4494 10696
rect 4798 10684 4804 10696
rect 4856 10724 4862 10736
rect 4856 10696 5014 10724
rect 4856 10684 4862 10696
rect 4238 10659 4296 10665
rect 4238 10656 4250 10659
rect 4172 10628 4250 10656
rect 2317 10619 2375 10625
rect 4238 10625 4250 10628
rect 4284 10625 4296 10659
rect 4238 10619 4296 10625
rect 2406 10588 2412 10600
rect 2367 10560 2412 10588
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 2685 10591 2743 10597
rect 2685 10557 2697 10591
rect 2731 10588 2743 10591
rect 4522 10588 4528 10600
rect 2731 10560 4108 10588
rect 4483 10560 4528 10588
rect 2731 10557 2743 10560
rect 2685 10551 2743 10557
rect 1489 10523 1547 10529
rect 1489 10489 1501 10523
rect 1535 10520 1547 10523
rect 4080 10520 4108 10560
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 5828 10588 5856 10764
rect 6914 10684 6920 10736
rect 6972 10724 6978 10736
rect 7852 10724 7880 10764
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 9214 10792 9220 10804
rect 8711 10764 9220 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 6972 10696 7038 10724
rect 7852 10696 9045 10724
rect 6972 10684 6978 10696
rect 9033 10693 9045 10696
rect 9079 10693 9091 10727
rect 9033 10687 9091 10693
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5960 10628 6285 10656
rect 5960 10616 5966 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 8110 10656 8116 10668
rect 8071 10628 8116 10656
rect 6273 10619 6331 10625
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 4672 10560 5856 10588
rect 6288 10560 6653 10588
rect 4672 10548 4678 10560
rect 6288 10520 6316 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8720 10560 9137 10588
rect 8720 10548 8726 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 1535 10492 2268 10520
rect 4080 10492 4384 10520
rect 1535 10489 1547 10492
rect 1489 10483 1547 10489
rect 2240 10452 2268 10492
rect 4062 10452 4068 10464
rect 2240 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4356 10452 4384 10492
rect 6012 10492 6316 10520
rect 8573 10523 8631 10529
rect 6012 10461 6040 10492
rect 8573 10489 8585 10523
rect 8619 10520 8631 10523
rect 9232 10520 9260 10551
rect 9306 10520 9312 10532
rect 8619 10492 9312 10520
rect 8619 10489 8631 10492
rect 8573 10483 8631 10489
rect 9306 10480 9312 10492
rect 9364 10480 9370 10532
rect 5997 10455 6055 10461
rect 5997 10452 6009 10455
rect 4212 10424 4257 10452
rect 4356 10424 6009 10452
rect 4212 10412 4218 10424
rect 5997 10421 6009 10424
rect 6043 10421 6055 10455
rect 5997 10415 6055 10421
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 5666 10362
rect 5718 10310 5730 10362
rect 5782 10310 5794 10362
rect 5846 10310 5858 10362
rect 5910 10310 5922 10362
rect 5974 10310 8766 10362
rect 8818 10310 8830 10362
rect 8882 10310 8894 10362
rect 8946 10310 8958 10362
rect 9010 10310 9022 10362
rect 9074 10310 9844 10362
rect 920 10288 9844 10310
rect 1765 10251 1823 10257
rect 1765 10217 1777 10251
rect 1811 10248 1823 10251
rect 1946 10248 1952 10260
rect 1811 10220 1952 10248
rect 1811 10217 1823 10220
rect 1765 10211 1823 10217
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2130 10248 2136 10260
rect 2091 10220 2136 10248
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 2685 10251 2743 10257
rect 2685 10217 2697 10251
rect 2731 10248 2743 10251
rect 3510 10248 3516 10260
rect 2731 10220 3516 10248
rect 2731 10217 2743 10220
rect 2685 10211 2743 10217
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 7377 10251 7435 10257
rect 7377 10248 7389 10251
rect 4172 10220 7389 10248
rect 1854 10140 1860 10192
rect 1912 10180 1918 10192
rect 2409 10183 2467 10189
rect 2409 10180 2421 10183
rect 1912 10152 2421 10180
rect 1912 10140 1918 10152
rect 2409 10149 2421 10152
rect 2455 10149 2467 10183
rect 2958 10180 2964 10192
rect 2919 10152 2964 10180
rect 2409 10143 2467 10149
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 3970 10112 3976 10124
rect 2746 10084 3976 10112
rect 1946 10004 1952 10056
rect 2004 10044 2010 10056
rect 2041 10047 2099 10053
rect 2041 10044 2053 10047
rect 2004 10016 2053 10044
rect 2004 10004 2010 10016
rect 2041 10013 2053 10016
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2498 10044 2504 10056
rect 2363 10016 2504 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2746 10044 2774 10084
rect 3970 10072 3976 10084
rect 4028 10072 4034 10124
rect 3050 10054 3056 10056
rect 2884 10053 3056 10054
rect 2639 10016 2774 10044
rect 2869 10047 3056 10053
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 2869 10013 2881 10047
rect 2915 10026 3056 10047
rect 2915 10013 2927 10026
rect 2869 10007 2927 10013
rect 3050 10004 3056 10026
rect 3108 10004 3114 10056
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10013 3203 10047
rect 3145 10007 3203 10013
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 1762 9936 1768 9988
rect 1820 9976 1826 9988
rect 1820 9948 2360 9976
rect 3160 9970 3188 10007
rect 1820 9936 1826 9948
rect 1857 9911 1915 9917
rect 1857 9877 1869 9911
rect 1903 9908 1915 9911
rect 2222 9908 2228 9920
rect 1903 9880 2228 9908
rect 1903 9877 1915 9880
rect 1857 9871 1915 9877
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 2332 9908 2360 9948
rect 3068 9942 3188 9970
rect 3436 9976 3464 10007
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 4172 10053 4200 10220
rect 7377 10217 7389 10220
rect 7423 10217 7435 10251
rect 7377 10211 7435 10217
rect 7561 10251 7619 10257
rect 7561 10217 7573 10251
rect 7607 10248 7619 10251
rect 7607 10220 7641 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 4249 10183 4307 10189
rect 4249 10149 4261 10183
rect 4295 10180 4307 10183
rect 4295 10152 4660 10180
rect 4295 10149 4307 10152
rect 4249 10143 4307 10149
rect 4632 10121 4660 10152
rect 5902 10140 5908 10192
rect 5960 10180 5966 10192
rect 5960 10152 6500 10180
rect 5960 10140 5966 10152
rect 4617 10115 4675 10121
rect 4617 10081 4629 10115
rect 4663 10081 4675 10115
rect 6472 10112 6500 10152
rect 6822 10140 6828 10192
rect 6880 10180 6886 10192
rect 6917 10183 6975 10189
rect 6917 10180 6929 10183
rect 6880 10152 6929 10180
rect 6880 10140 6886 10152
rect 6917 10149 6929 10152
rect 6963 10149 6975 10183
rect 6917 10143 6975 10149
rect 7006 10140 7012 10192
rect 7064 10180 7070 10192
rect 7190 10180 7196 10192
rect 7064 10152 7196 10180
rect 7064 10140 7070 10152
rect 7190 10140 7196 10152
rect 7248 10180 7254 10192
rect 7576 10180 7604 10211
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 8352 10220 8769 10248
rect 8352 10208 8358 10220
rect 8757 10217 8769 10220
rect 8803 10217 8815 10251
rect 8757 10211 8815 10217
rect 8018 10180 8024 10192
rect 7248 10152 8024 10180
rect 7248 10140 7254 10152
rect 8018 10140 8024 10152
rect 8076 10140 8082 10192
rect 8389 10115 8447 10121
rect 8389 10112 8401 10115
rect 6472 10084 8401 10112
rect 4617 10075 4675 10081
rect 8389 10081 8401 10084
rect 8435 10081 8447 10115
rect 9306 10112 9312 10124
rect 9267 10084 9312 10112
rect 8389 10075 8447 10081
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 3881 10047 3939 10053
rect 3881 10044 3893 10047
rect 3752 10016 3893 10044
rect 3752 10004 3758 10016
rect 3881 10013 3893 10016
rect 3927 10013 3939 10047
rect 3881 10007 3939 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 4522 10044 4528 10056
rect 4479 10016 4528 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4982 10044 4988 10056
rect 4943 10016 4988 10044
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 3786 9976 3792 9988
rect 3436 9948 3792 9976
rect 3068 9908 3096 9942
rect 3786 9936 3792 9948
rect 3844 9936 3850 9988
rect 5534 9936 5540 9988
rect 5592 9936 5598 9988
rect 3234 9908 3240 9920
rect 2332 9880 3096 9908
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 3697 9911 3755 9917
rect 3697 9908 3709 9911
rect 3660 9880 3709 9908
rect 3660 9868 3666 9880
rect 3697 9877 3709 9880
rect 3743 9877 3755 9911
rect 3697 9871 3755 9877
rect 3973 9911 4031 9917
rect 3973 9877 3985 9911
rect 4019 9908 4031 9911
rect 6472 9908 6500 10007
rect 6546 10004 6552 10056
rect 6604 10044 6610 10056
rect 7466 10044 7472 10056
rect 6604 10016 7328 10044
rect 7427 10016 7472 10044
rect 6604 10004 6610 10016
rect 7006 9976 7012 9988
rect 6967 9948 7012 9976
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 7190 9976 7196 9988
rect 7151 9948 7196 9976
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 7300 9976 7328 10016
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 7576 10016 9137 10044
rect 7576 9976 7604 10016
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 8018 9976 8024 9988
rect 7300 9948 7604 9976
rect 7979 9948 8024 9976
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 8205 9979 8263 9985
rect 8205 9976 8217 9979
rect 8168 9948 8217 9976
rect 8168 9936 8174 9948
rect 8205 9945 8217 9948
rect 8251 9945 8263 9979
rect 9214 9976 9220 9988
rect 9175 9948 9220 9976
rect 8205 9939 8263 9945
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 4019 9880 6500 9908
rect 4019 9877 4031 9880
rect 3973 9871 4031 9877
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 7929 9911 7987 9917
rect 7929 9908 7941 9911
rect 6696 9880 7941 9908
rect 6696 9868 6702 9880
rect 7929 9877 7941 9880
rect 7975 9877 7987 9911
rect 7929 9871 7987 9877
rect 920 9818 9844 9840
rect 920 9766 4116 9818
rect 4168 9766 4180 9818
rect 4232 9766 4244 9818
rect 4296 9766 4308 9818
rect 4360 9766 4372 9818
rect 4424 9766 7216 9818
rect 7268 9766 7280 9818
rect 7332 9766 7344 9818
rect 7396 9766 7408 9818
rect 7460 9766 7472 9818
rect 7524 9766 9844 9818
rect 920 9744 9844 9766
rect 2409 9707 2467 9713
rect 2409 9673 2421 9707
rect 2455 9673 2467 9707
rect 3142 9704 3148 9716
rect 2409 9667 2467 9673
rect 2792 9676 3148 9704
rect 2314 9636 2320 9648
rect 2275 9608 2320 9636
rect 2314 9596 2320 9608
rect 2372 9596 2378 9648
rect 2424 9636 2452 9667
rect 2792 9636 2820 9676
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 3712 9676 5304 9704
rect 3712 9636 3740 9676
rect 2424 9608 2820 9636
rect 2884 9608 3740 9636
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2280 9540 2605 9568
rect 2280 9528 2286 9540
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9568 2835 9571
rect 2884 9568 2912 9608
rect 4430 9596 4436 9648
rect 4488 9596 4494 9648
rect 5276 9642 5304 9676
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 6641 9707 6699 9713
rect 6641 9704 6653 9707
rect 5592 9676 6653 9704
rect 5592 9664 5598 9676
rect 6641 9673 6653 9676
rect 6687 9673 6699 9707
rect 6641 9667 6699 9673
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 8110 9704 8116 9716
rect 7616 9676 8116 9704
rect 7616 9664 7622 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 5276 9636 5488 9642
rect 8021 9639 8079 9645
rect 8021 9636 8033 9639
rect 5276 9614 8033 9636
rect 5460 9608 8033 9614
rect 8021 9605 8033 9608
rect 8067 9605 8079 9639
rect 8021 9599 8079 9605
rect 2823 9540 2912 9568
rect 2823 9537 2835 9540
rect 2777 9531 2835 9537
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2700 9500 2728 9531
rect 2958 9528 2964 9580
rect 3016 9568 3022 9580
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 3016 9540 3341 9568
rect 3016 9528 3022 9540
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3651 9540 3832 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 2096 9472 2728 9500
rect 2096 9460 2102 9472
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3620 9500 3648 9531
rect 3292 9472 3648 9500
rect 3697 9503 3755 9509
rect 3292 9460 3298 9472
rect 3697 9469 3709 9503
rect 3743 9469 3755 9503
rect 3804 9500 3832 9540
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3936 9540 4077 9568
rect 3936 9528 3942 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 4065 9531 4123 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5736 9540 6193 9568
rect 4706 9500 4712 9512
rect 3804 9472 4712 9500
rect 3697 9463 3755 9469
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 3145 9435 3203 9441
rect 2004 9404 2774 9432
rect 2004 9392 2010 9404
rect 2746 9364 2774 9404
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3712 9432 3740 9463
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 3191 9404 3740 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3326 9364 3332 9376
rect 2746 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 4522 9364 4528 9376
rect 3467 9336 4528 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5736 9364 5764 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 5994 9500 6000 9512
rect 5955 9472 6000 9500
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6196 9500 6224 9531
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6733 9571 6791 9577
rect 6733 9568 6745 9571
rect 6328 9540 6745 9568
rect 6328 9528 6334 9540
rect 6733 9537 6745 9540
rect 6779 9537 6791 9571
rect 6914 9568 6920 9580
rect 6875 9540 6920 9568
rect 6733 9531 6791 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9568 7435 9571
rect 7926 9568 7932 9580
rect 7423 9540 7932 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 8202 9568 8208 9580
rect 8163 9540 8208 9568
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 7006 9500 7012 9512
rect 6196 9472 7012 9500
rect 7006 9460 7012 9472
rect 7064 9460 7070 9512
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 8018 9460 8024 9512
rect 8076 9500 8082 9512
rect 8570 9500 8576 9512
rect 8076 9472 8576 9500
rect 8076 9460 8082 9472
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 6730 9392 6736 9444
rect 6788 9432 6794 9444
rect 7929 9435 7987 9441
rect 7929 9432 7941 9435
rect 6788 9404 7941 9432
rect 6788 9392 6794 9404
rect 7929 9401 7941 9404
rect 7975 9401 7987 9435
rect 7929 9395 7987 9401
rect 5132 9336 5764 9364
rect 5132 9324 5138 9336
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6273 9367 6331 9373
rect 6273 9364 6285 9367
rect 6052 9336 6285 9364
rect 6052 9324 6058 9336
rect 6273 9333 6285 9336
rect 6319 9364 6331 9367
rect 6914 9364 6920 9376
rect 6319 9336 6920 9364
rect 6319 9333 6331 9336
rect 6273 9327 6331 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7098 9364 7104 9376
rect 7059 9336 7104 9364
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7193 9367 7251 9373
rect 7193 9333 7205 9367
rect 7239 9364 7251 9367
rect 7650 9364 7656 9376
rect 7239 9336 7656 9364
rect 7239 9333 7251 9336
rect 7193 9327 7251 9333
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 5666 9274
rect 5718 9222 5730 9274
rect 5782 9222 5794 9274
rect 5846 9222 5858 9274
rect 5910 9222 5922 9274
rect 5974 9222 8766 9274
rect 8818 9222 8830 9274
rect 8882 9222 8894 9274
rect 8946 9222 8958 9274
rect 9010 9222 9022 9274
rect 9074 9222 9844 9274
rect 920 9200 9844 9222
rect 1762 9160 1768 9172
rect 1723 9132 1768 9160
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 4430 9160 4436 9172
rect 3620 9132 4436 9160
rect 2314 9052 2320 9104
rect 2372 9052 2378 9104
rect 2685 9095 2743 9101
rect 2685 9061 2697 9095
rect 2731 9092 2743 9095
rect 3620 9092 3648 9132
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 5353 9163 5411 9169
rect 5353 9160 5365 9163
rect 5040 9132 5365 9160
rect 5040 9120 5046 9132
rect 5353 9129 5365 9132
rect 5399 9129 5411 9163
rect 5353 9123 5411 9129
rect 2731 9064 3648 9092
rect 5368 9092 5396 9123
rect 5442 9120 5448 9172
rect 5500 9160 5506 9172
rect 8573 9163 8631 9169
rect 8573 9160 8585 9163
rect 5500 9132 8585 9160
rect 5500 9120 5506 9132
rect 8573 9129 8585 9132
rect 8619 9129 8631 9163
rect 8573 9123 8631 9129
rect 5368 9064 5580 9092
rect 2731 9061 2743 9064
rect 2685 9055 2743 9061
rect 2332 9024 2360 9052
rect 1412 8996 2360 9024
rect 1412 8965 1440 8996
rect 2498 8984 2504 9036
rect 2556 9024 2562 9036
rect 3605 9027 3663 9033
rect 3605 9024 3617 9027
rect 2556 8996 3617 9024
rect 2556 8984 2562 8996
rect 3605 8993 3617 8996
rect 3651 9024 3663 9027
rect 5166 9024 5172 9036
rect 3651 8996 5172 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1946 8956 1952 8968
rect 1907 8928 1952 8956
rect 1673 8919 1731 8925
rect 1688 8888 1716 8919
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 2590 8956 2596 8968
rect 2363 8928 2596 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 3142 8956 3148 8968
rect 3103 8928 3148 8956
rect 2869 8919 2927 8925
rect 2774 8888 2780 8900
rect 1688 8860 2780 8888
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 2884 8888 2912 8919
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 5092 8956 5120 8996
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5552 9024 5580 9064
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 7285 9095 7343 9101
rect 7285 9092 7297 9095
rect 6788 9064 7297 9092
rect 6788 9052 6794 9064
rect 7285 9061 7297 9064
rect 7331 9061 7343 9095
rect 7285 9055 7343 9061
rect 7466 9052 7472 9104
rect 7524 9052 7530 9104
rect 7653 9095 7711 9101
rect 7653 9061 7665 9095
rect 7699 9092 7711 9095
rect 13630 9092 13636 9104
rect 7699 9064 13636 9092
rect 7699 9061 7711 9064
rect 7653 9055 7711 9061
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 5552 8996 5733 9024
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 6086 8984 6092 9036
rect 6144 9024 6150 9036
rect 7484 9024 7512 9052
rect 6144 8996 7512 9024
rect 6144 8984 6150 8996
rect 8570 8984 8576 9036
rect 8628 9024 8634 9036
rect 8628 8996 8984 9024
rect 8628 8984 8634 8996
rect 5442 8956 5448 8968
rect 5092 8928 5448 8956
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 8018 8956 8024 8968
rect 7515 8928 8024 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8956 8171 8959
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 8159 8928 8217 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 3878 8888 3884 8900
rect 2884 8860 3740 8888
rect 3839 8860 3884 8888
rect 1213 8823 1271 8829
rect 1213 8789 1225 8823
rect 1259 8820 1271 8823
rect 1302 8820 1308 8832
rect 1259 8792 1308 8820
rect 1259 8789 1271 8792
rect 1213 8783 1271 8789
rect 1302 8780 1308 8792
rect 1360 8780 1366 8832
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 1489 8823 1547 8829
rect 1489 8820 1501 8823
rect 1452 8792 1501 8820
rect 1452 8780 1458 8792
rect 1489 8789 1501 8792
rect 1535 8789 1547 8823
rect 1489 8783 1547 8789
rect 1946 8780 1952 8832
rect 2004 8820 2010 8832
rect 2409 8823 2467 8829
rect 2409 8820 2421 8823
rect 2004 8792 2421 8820
rect 2004 8780 2010 8792
rect 2409 8789 2421 8792
rect 2455 8789 2467 8823
rect 3234 8820 3240 8832
rect 3195 8792 3240 8820
rect 2409 8783 2467 8789
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 3712 8820 3740 8860
rect 3878 8848 3884 8860
rect 3936 8848 3942 8900
rect 4890 8848 4896 8900
rect 4948 8848 4954 8900
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5224 8860 5948 8888
rect 5224 8848 5230 8860
rect 5810 8820 5816 8832
rect 3712 8792 5816 8820
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 5920 8820 5948 8860
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 7285 8891 7343 8897
rect 6052 8860 6210 8888
rect 6052 8848 6058 8860
rect 7285 8857 7297 8891
rect 7331 8888 7343 8891
rect 8128 8888 8156 8919
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8956 8965 8984 8996
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 8352 8928 8401 8956
rect 8352 8916 8358 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9398 8956 9404 8968
rect 9263 8928 9404 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 7331 8860 8156 8888
rect 7331 8857 7343 8860
rect 7285 8851 7343 8857
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 8757 8891 8815 8897
rect 8757 8888 8769 8891
rect 8628 8860 8769 8888
rect 8628 8848 8634 8860
rect 8757 8857 8769 8860
rect 8803 8857 8815 8891
rect 8757 8851 8815 8857
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 5920 8792 7205 8820
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 9122 8820 9128 8832
rect 9083 8792 9128 8820
rect 7193 8783 7251 8789
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9401 8823 9459 8829
rect 9401 8789 9413 8823
rect 9447 8820 9459 8823
rect 13538 8820 13544 8832
rect 9447 8792 13544 8820
rect 9447 8789 9459 8792
rect 9401 8783 9459 8789
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 920 8730 9844 8752
rect 920 8678 4116 8730
rect 4168 8678 4180 8730
rect 4232 8678 4244 8730
rect 4296 8678 4308 8730
rect 4360 8678 4372 8730
rect 4424 8678 7216 8730
rect 7268 8678 7280 8730
rect 7332 8678 7344 8730
rect 7396 8678 7408 8730
rect 7460 8678 7472 8730
rect 7524 8678 9844 8730
rect 920 8656 9844 8678
rect 1854 8576 1860 8628
rect 1912 8616 1918 8628
rect 3786 8616 3792 8628
rect 1912 8588 3792 8616
rect 1912 8576 1918 8588
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 4706 8625 4712 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 3936 8588 4353 8616
rect 3936 8576 3942 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 4663 8619 4712 8625
rect 4663 8585 4675 8619
rect 4709 8585 4712 8619
rect 4663 8579 4712 8585
rect 4706 8576 4712 8579
rect 4764 8576 4770 8628
rect 5810 8616 5816 8628
rect 5771 8588 5816 8616
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 8202 8616 8208 8628
rect 6227 8588 8208 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 9490 8616 9496 8628
rect 9451 8588 9496 8616
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 2222 8548 2228 8560
rect 2183 8520 2228 8548
rect 2222 8508 2228 8520
rect 2280 8548 2286 8560
rect 2869 8551 2927 8557
rect 2280 8520 2452 8548
rect 2280 8508 2286 8520
rect 1486 8440 1492 8492
rect 1544 8480 1550 8492
rect 1581 8483 1639 8489
rect 1581 8480 1593 8483
rect 1544 8452 1593 8480
rect 1544 8440 1550 8452
rect 1581 8449 1593 8452
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2424 8480 2452 8520
rect 2869 8517 2881 8551
rect 2915 8548 2927 8551
rect 2958 8548 2964 8560
rect 2915 8520 2964 8548
rect 2915 8517 2927 8520
rect 2501 8507 2559 8513
rect 2869 8511 2927 8517
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 3326 8508 3332 8560
rect 3384 8508 3390 8560
rect 7098 8548 7104 8560
rect 4264 8520 7104 8548
rect 2501 8480 2513 8507
rect 1903 8452 2360 8480
rect 2424 8473 2513 8480
rect 2547 8473 2559 8507
rect 2424 8467 2559 8473
rect 2424 8452 2544 8467
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2332 8412 2360 8452
rect 2096 8384 2268 8412
rect 2332 8384 2452 8412
rect 2096 8372 2102 8384
rect 1397 8347 1455 8353
rect 1397 8313 1409 8347
rect 1443 8344 1455 8347
rect 1578 8344 1584 8356
rect 1443 8316 1584 8344
rect 1443 8313 1455 8316
rect 1397 8307 1455 8313
rect 1578 8304 1584 8316
rect 1636 8304 1642 8356
rect 2240 8344 2268 8384
rect 2317 8347 2375 8353
rect 2317 8344 2329 8347
rect 2240 8316 2329 8344
rect 2317 8313 2329 8316
rect 2363 8313 2375 8347
rect 2424 8344 2452 8384
rect 2498 8372 2504 8424
rect 2556 8412 2562 8424
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 2556 8384 2605 8412
rect 2556 8372 2562 8384
rect 2593 8381 2605 8384
rect 2639 8381 2651 8415
rect 4264 8412 4292 8520
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 9214 8548 9220 8560
rect 8694 8520 9220 8548
rect 9214 8508 9220 8520
rect 9272 8508 9278 8560
rect 4338 8440 4344 8492
rect 4396 8480 4402 8492
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 4396 8452 5365 8480
rect 4396 8440 4402 8452
rect 5353 8449 5365 8452
rect 5399 8480 5411 8483
rect 6270 8480 6276 8492
rect 5399 8452 6276 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 2593 8375 2651 8381
rect 2700 8384 4292 8412
rect 4433 8415 4491 8421
rect 2700 8344 2728 8384
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4522 8412 4528 8424
rect 4479 8384 4528 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4522 8372 4528 8384
rect 4580 8412 4586 8424
rect 6380 8412 6408 8443
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 9033 8483 9091 8489
rect 6512 8452 6557 8480
rect 6512 8440 6518 8452
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9306 8480 9312 8492
rect 9079 8452 9312 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 22462 8480 22468 8492
rect 13780 8452 22468 8480
rect 13780 8440 13786 8452
rect 22462 8440 22468 8452
rect 22520 8440 22526 8492
rect 6730 8412 6736 8424
rect 4580 8384 5672 8412
rect 6380 8384 6736 8412
rect 4580 8372 4586 8384
rect 5534 8344 5540 8356
rect 2424 8316 2728 8344
rect 3896 8316 5540 8344
rect 2317 8307 2375 8313
rect 1673 8279 1731 8285
rect 1673 8245 1685 8279
rect 1719 8276 1731 8279
rect 3896 8276 3924 8316
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5644 8344 5672 8384
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 7190 8412 7196 8424
rect 7151 8384 7196 8412
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 8110 8412 8116 8424
rect 7607 8384 8116 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 22186 8412 22192 8424
rect 13872 8384 22192 8412
rect 13872 8372 13878 8384
rect 22186 8372 22192 8384
rect 22244 8372 22250 8424
rect 6546 8344 6552 8356
rect 5644 8316 6552 8344
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 7101 8347 7159 8353
rect 7101 8344 7113 8347
rect 6880 8316 7113 8344
rect 6880 8304 6886 8316
rect 7101 8313 7113 8316
rect 7147 8313 7159 8347
rect 7101 8307 7159 8313
rect 1719 8248 3924 8276
rect 1719 8245 1731 8248
rect 1673 8239 1731 8245
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5350 8276 5356 8288
rect 4948 8248 5356 8276
rect 4948 8236 4954 8248
rect 5350 8236 5356 8248
rect 5408 8276 5414 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5408 8248 5457 8276
rect 5408 8236 5414 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 5445 8239 5503 8245
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 22738 8276 22744 8288
rect 6052 8248 22744 8276
rect 6052 8236 6058 8248
rect 22738 8236 22744 8248
rect 22796 8236 22802 8288
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 5666 8186
rect 5718 8134 5730 8186
rect 5782 8134 5794 8186
rect 5846 8134 5858 8186
rect 5910 8134 5922 8186
rect 5974 8134 8766 8186
rect 8818 8134 8830 8186
rect 8882 8134 8894 8186
rect 8946 8134 8958 8186
rect 9010 8134 9022 8186
rect 9074 8134 9844 8186
rect 920 8112 9844 8134
rect 1670 8072 1676 8084
rect 1631 8044 1676 8072
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 3697 8075 3755 8081
rect 3697 8072 3709 8075
rect 2056 8044 2728 8072
rect 1397 8007 1455 8013
rect 1397 7973 1409 8007
rect 1443 8004 1455 8007
rect 1762 8004 1768 8016
rect 1443 7976 1768 8004
rect 1443 7973 1455 7976
rect 1397 7967 1455 7973
rect 1762 7964 1768 7976
rect 1820 7964 1826 8016
rect 1210 7896 1216 7948
rect 1268 7936 1274 7948
rect 1268 7908 1900 7936
rect 1268 7896 1274 7908
rect 1872 7877 1900 7908
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 1596 7800 1624 7831
rect 2056 7800 2084 8044
rect 2130 7964 2136 8016
rect 2188 8004 2194 8016
rect 2225 8007 2283 8013
rect 2225 8004 2237 8007
rect 2188 7976 2237 8004
rect 2188 7964 2194 7976
rect 2225 7973 2237 7976
rect 2271 7973 2283 8007
rect 2225 7967 2283 7973
rect 2406 7964 2412 8016
rect 2464 7964 2470 8016
rect 2700 8004 2728 8044
rect 2884 8044 3709 8072
rect 2884 8004 2912 8044
rect 3697 8041 3709 8044
rect 3743 8072 3755 8075
rect 5994 8072 6000 8084
rect 3743 8044 6000 8072
rect 3743 8041 3755 8044
rect 3697 8035 3755 8041
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 6454 8072 6460 8084
rect 6415 8044 6460 8072
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 7248 8044 8401 8072
rect 7248 8032 7254 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 8849 8075 8907 8081
rect 8849 8041 8861 8075
rect 8895 8041 8907 8075
rect 8849 8035 8907 8041
rect 4249 8007 4307 8013
rect 4249 8004 4261 8007
rect 2700 7976 2912 8004
rect 2976 7976 4261 8004
rect 2424 7936 2452 7964
rect 2976 7936 3004 7976
rect 4249 7973 4261 7976
rect 4295 8004 4307 8007
rect 4706 8004 4712 8016
rect 4295 7976 4712 8004
rect 4295 7973 4307 7976
rect 4249 7967 4307 7973
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8110 8004 8116 8016
rect 7984 7976 8116 8004
rect 7984 7964 7990 7976
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 8294 8004 8300 8016
rect 8255 7976 8300 8004
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 2332 7908 2452 7936
rect 2884 7908 3004 7936
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2332 7868 2360 7908
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 2332 7840 2421 7868
rect 2133 7831 2191 7837
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7837 2743 7871
rect 2884 7868 2912 7908
rect 3050 7896 3056 7948
rect 3108 7936 3114 7948
rect 3108 7908 3153 7936
rect 3108 7896 3114 7908
rect 3234 7896 3240 7948
rect 3292 7936 3298 7948
rect 3421 7939 3479 7945
rect 3421 7936 3433 7939
rect 3292 7908 3433 7936
rect 3292 7896 3298 7908
rect 3421 7905 3433 7908
rect 3467 7905 3479 7939
rect 3421 7899 3479 7905
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7936 5043 7939
rect 5074 7936 5080 7948
rect 5031 7908 5080 7936
rect 5031 7905 5043 7908
rect 4985 7899 5043 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 5500 7908 6561 7936
rect 5500 7896 5506 7908
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6822 7936 6828 7948
rect 6783 7908 6828 7936
rect 6549 7899 6607 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 8864 7936 8892 8035
rect 9214 8032 9220 8084
rect 9272 8072 9278 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 9272 8044 9321 8072
rect 9272 8032 9278 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 13446 7964 13452 8016
rect 13504 8004 13510 8016
rect 22278 8004 22284 8016
rect 13504 7976 22284 8004
rect 13504 7964 13510 7976
rect 22278 7964 22284 7976
rect 22336 7964 22342 8016
rect 6972 7908 8892 7936
rect 9217 7939 9275 7945
rect 6972 7896 6978 7908
rect 9217 7905 9229 7939
rect 9263 7905 9275 7939
rect 22370 7936 22376 7948
rect 9217 7899 9275 7905
rect 12406 7908 22376 7936
rect 2685 7831 2743 7837
rect 2792 7840 2912 7868
rect 2969 7867 3027 7873
rect 1596 7772 2084 7800
rect 2148 7744 2176 7831
rect 2700 7800 2728 7831
rect 2792 7800 2820 7840
rect 2969 7833 2981 7867
rect 3015 7864 3027 7867
rect 3015 7862 3096 7864
rect 3160 7862 3924 7868
rect 3015 7840 3924 7862
rect 3015 7836 3188 7840
rect 3015 7833 3027 7836
rect 3068 7834 3188 7836
rect 2969 7827 3027 7833
rect 3896 7812 3924 7840
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4709 7871 4767 7877
rect 4709 7868 4721 7871
rect 4120 7840 4721 7868
rect 4120 7828 4126 7840
rect 4709 7837 4721 7840
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 8573 7871 8631 7877
rect 8573 7868 8585 7871
rect 8260 7840 8585 7868
rect 8260 7828 8266 7840
rect 8573 7837 8585 7840
rect 8619 7837 8631 7871
rect 8754 7868 8760 7880
rect 8715 7840 8760 7868
rect 8573 7831 8631 7837
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 9232 7868 9260 7899
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9232 7840 9505 7868
rect 9493 7837 9505 7840
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 3421 7803 3479 7809
rect 3421 7800 3433 7803
rect 2700 7772 2820 7800
rect 3252 7772 3433 7800
rect 3252 7744 3280 7772
rect 3421 7769 3433 7772
rect 3467 7769 3479 7803
rect 3421 7763 3479 7769
rect 3510 7760 3516 7812
rect 3568 7800 3574 7812
rect 3789 7803 3847 7809
rect 3789 7800 3801 7803
rect 3568 7772 3801 7800
rect 3568 7760 3574 7772
rect 3789 7769 3801 7772
rect 3835 7769 3847 7803
rect 3789 7763 3847 7769
rect 3878 7760 3884 7812
rect 3936 7800 3942 7812
rect 3973 7803 4031 7809
rect 3973 7800 3985 7803
rect 3936 7772 3985 7800
rect 3936 7760 3942 7772
rect 3973 7769 3985 7772
rect 4019 7769 4031 7803
rect 3973 7763 4031 7769
rect 4246 7760 4252 7812
rect 4304 7800 4310 7812
rect 5074 7800 5080 7812
rect 4304 7772 5080 7800
rect 4304 7760 4310 7772
rect 1118 7692 1124 7744
rect 1176 7732 1182 7744
rect 1949 7735 2007 7741
rect 1949 7732 1961 7735
rect 1176 7704 1961 7732
rect 1176 7692 1182 7704
rect 1949 7701 1961 7704
rect 1995 7701 2007 7735
rect 1949 7695 2007 7701
rect 2130 7692 2136 7744
rect 2188 7692 2194 7744
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 2774 7732 2780 7744
rect 2735 7704 2780 7732
rect 2774 7692 2780 7704
rect 2832 7692 2838 7744
rect 3050 7732 3056 7744
rect 3011 7704 3056 7732
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 3234 7692 3240 7744
rect 3292 7692 3298 7744
rect 3329 7735 3387 7741
rect 3329 7701 3341 7735
rect 3375 7732 3387 7735
rect 4356 7732 4384 7772
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 5442 7760 5448 7812
rect 5500 7760 5506 7812
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7098 7800 7104 7812
rect 6972 7772 7104 7800
rect 6972 7760 6978 7772
rect 7098 7760 7104 7772
rect 7156 7800 7162 7812
rect 7156 7772 7314 7800
rect 7156 7760 7162 7772
rect 3375 7704 4384 7732
rect 4433 7735 4491 7741
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 4522 7732 4528 7744
rect 4479 7704 4528 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 12406 7732 12434 7908
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 4672 7704 12434 7732
rect 4672 7692 4678 7704
rect 920 7642 9844 7664
rect 920 7590 4116 7642
rect 4168 7590 4180 7642
rect 4232 7590 4244 7642
rect 4296 7590 4308 7642
rect 4360 7590 4372 7642
rect 4424 7590 7216 7642
rect 7268 7590 7280 7642
rect 7332 7590 7344 7642
rect 7396 7590 7408 7642
rect 7460 7590 7472 7642
rect 7524 7590 9844 7642
rect 920 7568 9844 7590
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 2608 7500 3249 7528
rect 2498 7420 2504 7472
rect 2556 7460 2562 7472
rect 2608 7460 2636 7500
rect 3237 7497 3249 7500
rect 3283 7528 3295 7531
rect 3283 7500 7788 7528
rect 3283 7497 3295 7500
rect 3237 7491 3295 7497
rect 3053 7463 3111 7469
rect 3053 7460 3065 7463
rect 2556 7432 2636 7460
rect 2792 7432 3065 7460
rect 2556 7420 2562 7432
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7392 1547 7395
rect 1670 7392 1676 7404
rect 1535 7364 1676 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 1946 7392 1952 7404
rect 1811 7364 1952 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2317 7396 2375 7401
rect 2685 7396 2743 7401
rect 2792 7396 2820 7432
rect 3053 7429 3065 7432
rect 3099 7460 3111 7463
rect 4614 7460 4620 7472
rect 3099 7432 4620 7460
rect 3099 7429 3111 7432
rect 3053 7423 3111 7429
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 5350 7420 5356 7472
rect 5408 7420 5414 7472
rect 7760 7460 7788 7500
rect 8018 7488 8024 7540
rect 8076 7528 8082 7540
rect 8481 7531 8539 7537
rect 8481 7528 8493 7531
rect 8076 7500 8493 7528
rect 8076 7488 8082 7500
rect 8481 7497 8493 7500
rect 8527 7497 8539 7531
rect 9306 7528 9312 7540
rect 9267 7500 9312 7528
rect 8481 7491 8539 7497
rect 2317 7395 2452 7396
rect 2317 7361 2329 7395
rect 2363 7392 2452 7395
rect 2685 7395 2820 7396
rect 2363 7368 2636 7392
rect 2363 7361 2375 7368
rect 2424 7364 2636 7368
rect 2317 7355 2375 7361
rect 1026 7216 1032 7268
rect 1084 7256 1090 7268
rect 1581 7259 1639 7265
rect 1581 7256 1593 7259
rect 1084 7228 1593 7256
rect 1084 7216 1090 7228
rect 1581 7225 1593 7228
rect 1627 7225 1639 7259
rect 2056 7256 2084 7355
rect 2608 7324 2636 7364
rect 2685 7361 2697 7395
rect 2731 7368 2820 7395
rect 2731 7361 2743 7368
rect 2685 7355 2743 7361
rect 3234 7352 3240 7404
rect 3292 7352 3298 7404
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 3881 7395 3939 7401
rect 3881 7392 3893 7395
rect 3568 7364 3893 7392
rect 3568 7352 3574 7364
rect 3881 7361 3893 7364
rect 3927 7361 3939 7395
rect 3881 7355 3939 7361
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 4028 7364 4077 7392
rect 4028 7352 4034 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6512 7364 6561 7392
rect 6512 7352 6518 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 7668 7392 7696 7446
rect 7760 7432 8294 7460
rect 7834 7392 7840 7404
rect 7668 7364 7840 7392
rect 6549 7355 6607 7361
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 2777 7327 2835 7333
rect 2777 7324 2789 7327
rect 2608 7296 2789 7324
rect 2777 7293 2789 7296
rect 2823 7293 2835 7327
rect 3252 7324 3280 7352
rect 4341 7327 4399 7333
rect 3252 7296 4016 7324
rect 2777 7287 2835 7293
rect 3786 7256 3792 7268
rect 2056 7228 3792 7256
rect 1581 7219 1639 7225
rect 3786 7216 3792 7228
rect 3844 7216 3850 7268
rect 1210 7148 1216 7200
rect 1268 7188 1274 7200
rect 1305 7191 1363 7197
rect 1305 7188 1317 7191
rect 1268 7160 1317 7188
rect 1268 7148 1274 7160
rect 1305 7157 1317 7160
rect 1351 7157 1363 7191
rect 1305 7151 1363 7157
rect 1394 7148 1400 7200
rect 1452 7188 1458 7200
rect 1670 7188 1676 7200
rect 1452 7160 1676 7188
rect 1452 7148 1458 7160
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 2038 7188 2044 7200
rect 1903 7160 2044 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 2188 7160 2233 7188
rect 2188 7148 2194 7160
rect 2406 7148 2412 7200
rect 2464 7188 2470 7200
rect 2501 7191 2559 7197
rect 2501 7188 2513 7191
rect 2464 7160 2513 7188
rect 2464 7148 2470 7160
rect 2501 7157 2513 7160
rect 2547 7157 2559 7191
rect 2501 7151 2559 7157
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 3605 7191 3663 7197
rect 3605 7188 3617 7191
rect 2823 7160 3617 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 3605 7157 3617 7160
rect 3651 7188 3663 7191
rect 3878 7188 3884 7200
rect 3651 7160 3884 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 3988 7188 4016 7296
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 5534 7324 5540 7336
rect 4387 7296 5540 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 6822 7324 6828 7336
rect 6227 7296 6828 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 5813 7259 5871 7265
rect 5813 7256 5825 7259
rect 5500 7228 5825 7256
rect 5500 7216 5506 7228
rect 5813 7225 5825 7228
rect 5859 7225 5871 7259
rect 5813 7219 5871 7225
rect 8036 7188 8064 7355
rect 8266 7324 8294 7432
rect 8496 7392 8524 7491
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8496 7364 8769 7392
rect 8757 7361 8769 7364
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 9122 7352 9128 7404
rect 9180 7392 9186 7404
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 9180 7364 9505 7392
rect 9180 7352 9186 7364
rect 9493 7361 9505 7364
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 8266 7296 12434 7324
rect 8202 7216 8208 7268
rect 8260 7256 8266 7268
rect 9217 7259 9275 7265
rect 9217 7256 9229 7259
rect 8260 7228 9229 7256
rect 8260 7216 8266 7228
rect 9217 7225 9229 7228
rect 9263 7225 9275 7259
rect 9217 7219 9275 7225
rect 3988 7160 8064 7188
rect 9033 7191 9091 7197
rect 9033 7157 9045 7191
rect 9079 7188 9091 7191
rect 9582 7188 9588 7200
rect 9079 7160 9588 7188
rect 9079 7157 9091 7160
rect 9033 7151 9091 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 5666 7098
rect 5718 7046 5730 7098
rect 5782 7046 5794 7098
rect 5846 7046 5858 7098
rect 5910 7046 5922 7098
rect 5974 7046 8766 7098
rect 8818 7046 8830 7098
rect 8882 7046 8894 7098
rect 8946 7046 8958 7098
rect 9010 7046 9022 7098
rect 9074 7046 9844 7098
rect 920 7024 9844 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 3234 6984 3240 6996
rect 1636 6956 3240 6984
rect 1636 6944 1642 6956
rect 3234 6944 3240 6956
rect 3292 6944 3298 6996
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 3936 6956 5580 6984
rect 3936 6944 3942 6956
rect 5552 6916 5580 6956
rect 7098 6944 7104 6996
rect 7156 6984 7162 6996
rect 7742 6984 7748 6996
rect 7156 6956 7748 6984
rect 7156 6944 7162 6956
rect 7742 6944 7748 6956
rect 7800 6984 7806 6996
rect 8113 6987 8171 6993
rect 8113 6984 8125 6987
rect 7800 6956 8125 6984
rect 7800 6944 7806 6956
rect 8113 6953 8125 6956
rect 8159 6953 8171 6987
rect 12406 6984 12434 7296
rect 13814 7080 13820 7132
rect 13872 7120 13878 7132
rect 19794 7120 19800 7132
rect 13872 7092 19800 7120
rect 13872 7080 13878 7092
rect 19794 7080 19800 7092
rect 19852 7080 19858 7132
rect 13630 6984 13636 6996
rect 12406 6956 13636 6984
rect 8113 6947 8171 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 9582 6916 9588 6928
rect 5552 6888 9588 6916
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 3878 6848 3884 6860
rect 1719 6820 3884 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 5905 6851 5963 6857
rect 5905 6817 5917 6851
rect 5951 6848 5963 6851
rect 6178 6848 6184 6860
rect 5951 6820 6184 6848
rect 5951 6817 5963 6820
rect 5905 6811 5963 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6454 6808 6460 6860
rect 6512 6848 6518 6860
rect 9306 6848 9312 6860
rect 6512 6820 9168 6848
rect 9267 6820 9312 6848
rect 6512 6808 6518 6820
rect 9140 6792 9168 6820
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6749 1639 6783
rect 1581 6743 1639 6749
rect 1305 6715 1363 6721
rect 1305 6681 1317 6715
rect 1351 6712 1363 6715
rect 1596 6712 1624 6743
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3605 6783 3663 6789
rect 3605 6780 3617 6783
rect 3292 6752 3617 6780
rect 3292 6740 3298 6752
rect 3605 6749 3617 6752
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3844 6752 3985 6780
rect 3844 6740 3850 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 3973 6743 4031 6749
rect 5184 6752 5457 6780
rect 1351 6684 1624 6712
rect 1351 6681 1363 6684
rect 1305 6675 1363 6681
rect 1394 6644 1400 6656
rect 1355 6616 1400 6644
rect 1394 6604 1400 6616
rect 1452 6604 1458 6656
rect 1596 6644 1624 6684
rect 1854 6672 1860 6724
rect 1912 6712 1918 6724
rect 1949 6715 2007 6721
rect 1949 6712 1961 6715
rect 1912 6684 1961 6712
rect 1912 6672 1918 6684
rect 1949 6681 1961 6684
rect 1995 6681 2007 6715
rect 1949 6675 2007 6681
rect 2590 6644 2596 6656
rect 1596 6616 2596 6644
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 3160 6644 3188 6698
rect 5074 6672 5080 6724
rect 5132 6672 5138 6724
rect 3234 6644 3240 6656
rect 3160 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6644 3479 6647
rect 3786 6644 3792 6656
rect 3467 6616 3792 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 5184 6644 5212 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 8294 6780 8300 6792
rect 8076 6752 8300 6780
rect 8076 6740 8082 6752
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 8846 6780 8852 6792
rect 8444 6752 8852 6780
rect 8444 6740 8450 6752
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 9122 6780 9128 6792
rect 9035 6752 9128 6780
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 6181 6715 6239 6721
rect 6181 6681 6193 6715
rect 6227 6712 6239 6715
rect 22094 6712 22100 6724
rect 6227 6684 22100 6712
rect 6227 6681 6239 6684
rect 6181 6675 6239 6681
rect 22094 6672 22100 6684
rect 22152 6672 22158 6724
rect 3936 6616 5212 6644
rect 3936 6604 3942 6616
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 7469 6647 7527 6653
rect 7469 6644 7481 6647
rect 5316 6616 7481 6644
rect 5316 6604 5322 6616
rect 7469 6613 7481 6616
rect 7515 6613 7527 6647
rect 7469 6607 7527 6613
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 8481 6647 8539 6653
rect 8481 6644 8493 6647
rect 8076 6616 8493 6644
rect 8076 6604 8082 6616
rect 8481 6613 8493 6616
rect 8527 6613 8539 6647
rect 8481 6607 8539 6613
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8720 6616 8769 6644
rect 8720 6604 8726 6616
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9217 6647 9275 6653
rect 9217 6644 9229 6647
rect 8904 6616 9229 6644
rect 8904 6604 8910 6616
rect 9217 6613 9229 6616
rect 9263 6613 9275 6647
rect 9217 6607 9275 6613
rect 920 6554 9844 6576
rect 920 6502 4116 6554
rect 4168 6502 4180 6554
rect 4232 6502 4244 6554
rect 4296 6502 4308 6554
rect 4360 6502 4372 6554
rect 4424 6502 7216 6554
rect 7268 6502 7280 6554
rect 7332 6502 7344 6554
rect 7396 6502 7408 6554
rect 7460 6502 7472 6554
rect 7524 6502 9844 6554
rect 920 6480 9844 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2188 6412 2697 6440
rect 2188 6400 2194 6412
rect 2685 6409 2697 6412
rect 2731 6409 2743 6443
rect 5258 6440 5264 6452
rect 2685 6403 2743 6409
rect 3436 6412 5264 6440
rect 1302 6332 1308 6384
rect 1360 6372 1366 6384
rect 2866 6372 2872 6384
rect 1360 6344 2872 6372
rect 1360 6332 1366 6344
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 3436 6381 3464 6412
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 8665 6443 8723 6449
rect 8665 6440 8677 6443
rect 8444 6412 8677 6440
rect 8444 6400 8450 6412
rect 8665 6409 8677 6412
rect 8711 6409 8723 6443
rect 8665 6403 8723 6409
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 9180 6412 9225 6440
rect 9180 6400 9186 6412
rect 3421 6375 3479 6381
rect 3421 6341 3433 6375
rect 3467 6341 3479 6375
rect 3421 6335 3479 6341
rect 3605 6375 3663 6381
rect 3605 6341 3617 6375
rect 3651 6372 3663 6375
rect 3970 6372 3976 6384
rect 3651 6344 3976 6372
rect 3651 6341 3663 6344
rect 3605 6335 3663 6341
rect 3970 6332 3976 6344
rect 4028 6332 4034 6384
rect 6270 6372 6276 6384
rect 5658 6344 6276 6372
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 7708 6344 9352 6372
rect 7708 6332 7714 6344
rect 1210 6264 1216 6316
rect 1268 6304 1274 6316
rect 3142 6304 3148 6316
rect 1268 6276 3148 6304
rect 1268 6264 1274 6276
rect 3142 6264 3148 6276
rect 3200 6304 3206 6316
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3200 6276 3709 6304
rect 3200 6264 3206 6276
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 3927 6276 4108 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 4080 6236 4108 6276
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 4522 6304 4528 6316
rect 4212 6276 4257 6304
rect 4483 6276 4528 6304
rect 4212 6264 4218 6276
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 5994 6304 6000 6316
rect 5955 6276 6000 6304
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 6288 6276 7481 6304
rect 4890 6236 4896 6248
rect 3292 6208 4896 6236
rect 3292 6196 3298 6208
rect 4890 6196 4896 6208
rect 4948 6196 4954 6248
rect 1394 6128 1400 6180
rect 1452 6168 1458 6180
rect 4065 6171 4123 6177
rect 1452 6140 4016 6168
rect 1452 6128 1458 6140
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 3878 6100 3884 6112
rect 3660 6072 3884 6100
rect 3660 6060 3666 6072
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 3988 6100 4016 6140
rect 4065 6137 4077 6171
rect 4111 6168 4123 6171
rect 4154 6168 4160 6180
rect 4111 6140 4160 6168
rect 4111 6137 4123 6140
rect 4065 6131 4123 6137
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 6288 6100 6316 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 8202 6304 8208 6316
rect 7515 6276 8208 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 8343 6276 8616 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 6546 6236 6552 6248
rect 6507 6208 6552 6236
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6788 6208 6837 6236
rect 6788 6196 6794 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 7006 6196 7012 6248
rect 7064 6236 7070 6248
rect 8588 6236 8616 6276
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 9033 6307 9091 6313
rect 9033 6304 9045 6307
rect 8720 6276 9045 6304
rect 8720 6264 8726 6276
rect 9033 6273 9045 6276
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 9214 6236 9220 6248
rect 7064 6208 8432 6236
rect 8588 6208 9220 6236
rect 7064 6196 7070 6208
rect 6457 6171 6515 6177
rect 6457 6137 6469 6171
rect 6503 6168 6515 6171
rect 8294 6168 8300 6180
rect 6503 6140 8300 6168
rect 6503 6137 6515 6140
rect 6457 6131 6515 6137
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 7742 6100 7748 6112
rect 3988 6072 6316 6100
rect 7703 6072 7748 6100
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 7926 6100 7932 6112
rect 7887 6072 7932 6100
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8404 6100 8432 6208
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9324 6245 9352 6344
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6205 9367 6239
rect 9309 6199 9367 6205
rect 8481 6171 8539 6177
rect 8481 6137 8493 6171
rect 8527 6168 8539 6171
rect 13814 6168 13820 6180
rect 8527 6140 13820 6168
rect 8527 6137 8539 6140
rect 8481 6131 8539 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 9306 6100 9312 6112
rect 8404 6072 9312 6100
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 3036 6010 9844 6032
rect 3036 5958 5666 6010
rect 5718 5958 5730 6010
rect 5782 5958 5794 6010
rect 5846 5958 5858 6010
rect 5910 5958 5922 6010
rect 5974 5958 8766 6010
rect 8818 5958 8830 6010
rect 8882 5958 8894 6010
rect 8946 5958 8958 6010
rect 9010 5958 9022 6010
rect 9074 5958 9844 6010
rect 3036 5936 9844 5958
rect 3592 5899 3650 5905
rect 3592 5865 3604 5899
rect 3638 5896 3650 5899
rect 3786 5896 3792 5908
rect 3638 5868 3792 5896
rect 3638 5865 3650 5868
rect 3592 5859 3650 5865
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 4948 5868 5825 5896
rect 4948 5856 4954 5868
rect 4908 5828 4936 5856
rect 4724 5800 4936 5828
rect 1762 5720 1768 5772
rect 1820 5760 1826 5772
rect 2777 5763 2835 5769
rect 2777 5760 2789 5763
rect 1820 5732 2789 5760
rect 1820 5720 1826 5732
rect 2777 5729 2789 5732
rect 2823 5729 2835 5763
rect 2777 5723 2835 5729
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5760 3387 5763
rect 3970 5760 3976 5772
rect 3375 5732 3976 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 3050 5692 3056 5704
rect 1728 5664 3056 5692
rect 1728 5652 1734 5664
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 4724 5678 4752 5800
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5368 5760 5396 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 6270 5896 6276 5908
rect 6231 5868 6276 5896
rect 5813 5859 5871 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 8662 5896 8668 5908
rect 8623 5868 8668 5896
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 8941 5899 8999 5905
rect 8941 5865 8953 5899
rect 8987 5896 8999 5899
rect 9398 5896 9404 5908
rect 8987 5868 9404 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 5442 5788 5448 5840
rect 5500 5828 5506 5840
rect 5500 5800 6408 5828
rect 5500 5788 5506 5800
rect 6178 5760 6184 5772
rect 5316 5732 5396 5760
rect 6139 5732 6184 5760
rect 5316 5720 5322 5732
rect 5166 5692 5172 5704
rect 5127 5664 5172 5692
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5368 5701 5396 5732
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 6380 5760 6408 5800
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 8260 5800 8984 5828
rect 8260 5788 8266 5800
rect 7009 5763 7067 5769
rect 7009 5760 7021 5763
rect 6380 5732 7021 5760
rect 7009 5729 7021 5732
rect 7055 5729 7067 5763
rect 7009 5723 7067 5729
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5661 5411 5695
rect 5718 5692 5724 5704
rect 5679 5664 5724 5692
rect 5353 5655 5411 5661
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 6454 5692 6460 5704
rect 6415 5664 6460 5692
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6638 5692 6644 5704
rect 6599 5664 6644 5692
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 8478 5692 8484 5704
rect 8439 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8956 5692 8984 5800
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8956 5664 9045 5692
rect 9033 5661 9045 5664
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 1486 5584 1492 5636
rect 1544 5624 1550 5636
rect 1544 5596 2636 5624
rect 1544 5584 1550 5596
rect 2608 5352 2636 5596
rect 4982 5584 4988 5636
rect 5040 5624 5046 5636
rect 5537 5627 5595 5633
rect 5040 5596 5488 5624
rect 5040 5584 5046 5596
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 3752 5528 5089 5556
rect 3752 5516 3758 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5460 5556 5488 5596
rect 5537 5593 5549 5627
rect 5583 5624 5595 5627
rect 6362 5624 6368 5636
rect 5583 5596 6368 5624
rect 5583 5593 5595 5596
rect 5537 5587 5595 5593
rect 6362 5584 6368 5596
rect 6420 5584 6426 5636
rect 7558 5584 7564 5636
rect 7616 5584 7622 5636
rect 8938 5584 8944 5636
rect 8996 5624 9002 5636
rect 9217 5627 9275 5633
rect 9217 5624 9229 5627
rect 8996 5596 9229 5624
rect 8996 5584 9002 5596
rect 9217 5593 9229 5596
rect 9263 5593 9275 5627
rect 9217 5587 9275 5593
rect 9401 5559 9459 5565
rect 9401 5556 9413 5559
rect 5460 5528 9413 5556
rect 5077 5519 5135 5525
rect 9401 5525 9413 5528
rect 9447 5525 9459 5559
rect 9401 5519 9459 5525
rect 3036 5466 9844 5488
rect 3036 5414 4116 5466
rect 4168 5414 4180 5466
rect 4232 5414 4244 5466
rect 4296 5414 4308 5466
rect 4360 5414 4372 5466
rect 4424 5414 7216 5466
rect 7268 5414 7280 5466
rect 7332 5414 7344 5466
rect 7396 5414 7408 5466
rect 7460 5414 7472 5466
rect 7524 5414 9844 5466
rect 3036 5392 9844 5414
rect 3329 5355 3387 5361
rect 3329 5352 3341 5355
rect 2608 5324 3341 5352
rect 3329 5321 3341 5324
rect 3375 5321 3387 5355
rect 6178 5352 6184 5364
rect 3329 5315 3387 5321
rect 3896 5324 6184 5352
rect 3896 5284 3924 5324
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 8662 5352 8668 5364
rect 7892 5324 8668 5352
rect 7892 5312 7898 5324
rect 8662 5312 8668 5324
rect 8720 5352 8726 5364
rect 8938 5352 8944 5364
rect 8720 5324 8944 5352
rect 8720 5312 8726 5324
rect 8938 5312 8944 5324
rect 8996 5352 9002 5364
rect 8996 5324 9352 5352
rect 8996 5312 9002 5324
rect 3804 5256 3924 5284
rect 3804 5225 3832 5256
rect 5258 5244 5264 5296
rect 5316 5244 5322 5296
rect 7098 5244 7104 5296
rect 7156 5244 7162 5296
rect 8386 5244 8392 5296
rect 8444 5284 8450 5296
rect 9324 5293 9352 5324
rect 9125 5287 9183 5293
rect 9125 5284 9137 5287
rect 8444 5256 9137 5284
rect 8444 5244 8450 5256
rect 9125 5253 9137 5256
rect 9171 5253 9183 5287
rect 9125 5247 9183 5253
rect 9309 5287 9367 5293
rect 9309 5253 9321 5287
rect 9355 5253 9367 5287
rect 9309 5247 9367 5253
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 2915 5188 3525 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 3513 5185 3525 5188
rect 3559 5185 3571 5219
rect 3513 5179 3571 5185
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5185 3847 5219
rect 3970 5216 3976 5228
rect 3931 5188 3976 5216
rect 3789 5179 3847 5185
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 5736 5188 6193 5216
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 5534 5148 5540 5160
rect 4295 5120 5540 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 5736 5157 5764 5188
rect 6181 5185 6193 5188
rect 6227 5185 6239 5219
rect 7650 5216 7656 5228
rect 7611 5188 7656 5216
rect 6181 5179 6239 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 8294 5216 8300 5228
rect 8255 5188 8300 5216
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 8628 5188 8677 5216
rect 8628 5176 8634 5188
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5216 8907 5219
rect 9324 5216 9352 5247
rect 8895 5188 9352 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 5684 5120 5733 5148
rect 5684 5108 5690 5120
rect 5721 5117 5733 5120
rect 5767 5117 5779 5151
rect 5721 5111 5779 5117
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6730 5148 6736 5160
rect 5859 5120 6736 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 5258 5040 5264 5092
rect 5316 5080 5322 5092
rect 5902 5080 5908 5092
rect 5316 5052 5908 5080
rect 5316 5040 5322 5052
rect 5902 5040 5908 5052
rect 5960 5040 5966 5092
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 13722 5080 13728 5092
rect 8527 5052 13728 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 13722 5040 13728 5052
rect 13780 5040 13786 5092
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 4982 5012 4988 5024
rect 3651 4984 4988 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7892 4984 8125 5012
rect 7892 4972 7898 4984
rect 8113 4981 8125 4984
rect 8159 4981 8171 5015
rect 8113 4975 8171 4981
rect 9033 5015 9091 5021
rect 9033 4981 9045 5015
rect 9079 5012 9091 5015
rect 9398 5012 9404 5024
rect 9079 4984 9404 5012
rect 9079 4981 9091 4984
rect 9033 4975 9091 4981
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 9548 4984 9593 5012
rect 9548 4972 9554 4984
rect 3036 4922 9844 4944
rect 3036 4870 5666 4922
rect 5718 4870 5730 4922
rect 5782 4870 5794 4922
rect 5846 4870 5858 4922
rect 5910 4870 5922 4922
rect 5974 4870 8766 4922
rect 8818 4870 8830 4922
rect 8882 4870 8894 4922
rect 8946 4870 8958 4922
rect 9010 4870 9022 4922
rect 9074 4870 9844 4922
rect 3036 4848 9844 4870
rect 5258 4808 5264 4820
rect 3896 4780 5264 4808
rect 3326 4700 3332 4752
rect 3384 4740 3390 4752
rect 3421 4743 3479 4749
rect 3421 4740 3433 4743
rect 3384 4712 3433 4740
rect 3384 4700 3390 4712
rect 3421 4709 3433 4712
rect 3467 4740 3479 4743
rect 3896 4740 3924 4780
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 3467 4712 3924 4740
rect 3467 4709 3479 4712
rect 3421 4703 3479 4709
rect 3528 4681 3556 4712
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 5828 4740 5856 4771
rect 5994 4768 6000 4820
rect 6052 4808 6058 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 6052 4780 6285 4808
rect 6052 4768 6058 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 6273 4771 6331 4777
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 9272 4780 9505 4808
rect 9272 4768 9278 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 5224 4712 5856 4740
rect 6181 4743 6239 4749
rect 5224 4700 5230 4712
rect 6181 4709 6193 4743
rect 6227 4740 6239 4743
rect 6454 4740 6460 4752
rect 6227 4712 6460 4740
rect 6227 4709 6239 4712
rect 6181 4703 6239 4709
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 6641 4743 6699 4749
rect 6641 4709 6653 4743
rect 6687 4709 6699 4743
rect 6641 4703 6699 4709
rect 6917 4743 6975 4749
rect 6917 4709 6929 4743
rect 6963 4740 6975 4743
rect 6963 4712 7236 4740
rect 6963 4709 6975 4712
rect 6917 4703 6975 4709
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 4065 4675 4123 4681
rect 3559 4644 3593 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 5074 4672 5080 4684
rect 4111 4644 5080 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 5074 4632 5080 4644
rect 5132 4632 5138 4684
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3697 4607 3755 4613
rect 3697 4604 3709 4607
rect 3292 4576 3709 4604
rect 3292 4564 3298 4576
rect 3697 4573 3709 4576
rect 3743 4573 3755 4607
rect 3697 4567 3755 4573
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4573 3847 4607
rect 5184 4590 5212 4700
rect 5534 4632 5540 4684
rect 5592 4632 5598 4684
rect 6656 4672 6684 4703
rect 7208 4681 7236 4712
rect 7193 4675 7251 4681
rect 6656 4644 7144 4672
rect 3789 4567 3847 4573
rect 2682 4496 2688 4548
rect 2740 4536 2746 4548
rect 2740 4496 2774 4536
rect 3418 4496 3424 4548
rect 3476 4536 3482 4548
rect 3804 4536 3832 4567
rect 3970 4536 3976 4548
rect 3476 4508 3976 4536
rect 3476 4496 3482 4508
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 5552 4536 5580 4632
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5684 4576 5733 4604
rect 5684 4564 5690 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 6362 4564 6368 4616
rect 6420 4604 6426 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6420 4576 6469 4604
rect 6420 4564 6426 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7116 4613 7144 4644
rect 7193 4641 7205 4675
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6788 4576 6837 4604
rect 6788 4564 6794 4576
rect 6825 4573 6837 4576
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7101 4567 7159 4573
rect 7208 4576 7573 4604
rect 7208 4536 7236 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 8570 4564 8576 4616
rect 8628 4604 8634 4616
rect 9033 4607 9091 4613
rect 9033 4604 9045 4607
rect 8628 4576 9045 4604
rect 8628 4564 8634 4576
rect 9033 4573 9045 4576
rect 9079 4573 9091 4607
rect 9033 4567 9091 4573
rect 5552 4508 7236 4536
rect 8294 4496 8300 4548
rect 8352 4496 8358 4548
rect 2746 4264 2774 4496
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 6546 4468 6552 4480
rect 2915 4440 6552 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 6546 4428 6552 4440
rect 6604 4428 6610 4480
rect 3036 4378 9844 4400
rect 3036 4326 4116 4378
rect 4168 4326 4180 4378
rect 4232 4326 4244 4378
rect 4296 4326 4308 4378
rect 4360 4326 4372 4378
rect 4424 4326 7216 4378
rect 7268 4326 7280 4378
rect 7332 4326 7344 4378
rect 7396 4326 7408 4378
rect 7460 4326 7472 4378
rect 7524 4326 9844 4378
rect 3036 4304 9844 4326
rect 6086 4264 6092 4276
rect 2746 4236 6092 4264
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7156 4236 7573 4264
rect 7156 4224 7162 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 7561 4227 7619 4233
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 9309 4267 9367 4273
rect 9309 4264 9321 4267
rect 7708 4236 9321 4264
rect 7708 4224 7714 4236
rect 9309 4233 9321 4236
rect 9355 4233 9367 4267
rect 9309 4227 9367 4233
rect 3234 4156 3240 4208
rect 3292 4196 3298 4208
rect 3878 4196 3884 4208
rect 3292 4168 3884 4196
rect 3292 4156 3298 4168
rect 3878 4156 3884 4168
rect 3936 4156 3942 4208
rect 6546 4196 6552 4208
rect 3988 4168 4476 4196
rect 5934 4168 6552 4196
rect 3510 4088 3516 4140
rect 3568 4128 3574 4140
rect 3988 4137 4016 4168
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3568 4100 3709 4128
rect 3568 4088 3574 4100
rect 3697 4097 3709 4100
rect 3743 4128 3755 4131
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3743 4100 3985 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4448 4128 4476 4168
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 8570 4196 8576 4208
rect 7392 4168 8576 4196
rect 4798 4128 4804 4140
rect 4448 4100 4706 4128
rect 4759 4100 4804 4128
rect 4341 4091 4399 4097
rect 4356 4060 4384 4091
rect 3804 4032 4384 4060
rect 4433 4063 4491 4069
rect 3804 4001 3832 4032
rect 4433 4029 4445 4063
rect 4479 4029 4491 4063
rect 4678 4060 4706 4100
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 6273 4131 6331 4137
rect 6273 4097 6285 4131
rect 6319 4128 6331 4131
rect 6454 4128 6460 4140
rect 6319 4100 6460 4128
rect 6319 4097 6331 4100
rect 6273 4091 6331 4097
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 7190 4128 7196 4140
rect 7151 4100 7196 4128
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 5442 4060 5448 4072
rect 4678 4032 5448 4060
rect 4433 4023 4491 4029
rect 3789 3995 3847 4001
rect 3789 3961 3801 3995
rect 3835 3961 3847 3995
rect 3789 3955 3847 3961
rect 4157 3995 4215 4001
rect 4157 3961 4169 3995
rect 4203 3992 4215 3995
rect 4448 3992 4476 4023
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 6730 4060 6736 4072
rect 6420 4032 6736 4060
rect 6420 4020 6426 4032
rect 6730 4020 6736 4032
rect 6788 4020 6794 4072
rect 7392 4060 7420 4168
rect 8570 4156 8576 4168
rect 8628 4156 8634 4208
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 7650 4128 7656 4140
rect 7515 4100 7656 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 7024 4032 7420 4060
rect 7760 4060 7788 4091
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 7892 4100 7937 4128
rect 7892 4088 7898 4100
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8260 4100 8309 4128
rect 8260 4088 8266 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 8849 4131 8907 4137
rect 8849 4128 8861 4131
rect 8444 4100 8861 4128
rect 8444 4088 8450 4100
rect 8849 4097 8861 4100
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 9306 4128 9312 4140
rect 9079 4100 9312 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9456 4100 9505 4128
rect 9456 4088 9462 4100
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 7760 4032 8769 4060
rect 7024 4001 7052 4032
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 9180 4032 9229 4060
rect 9180 4020 9186 4032
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 4203 3964 4476 3992
rect 7009 3995 7067 4001
rect 4203 3961 4215 3964
rect 4157 3955 4215 3961
rect 7009 3961 7021 3995
rect 7055 3961 7067 3995
rect 7009 3955 7067 3961
rect 7285 3995 7343 4001
rect 7285 3961 7297 3995
rect 7331 3992 7343 3995
rect 8021 3995 8079 4001
rect 7331 3964 7696 3992
rect 7331 3961 7343 3964
rect 7285 3955 7343 3961
rect 3510 3924 3516 3936
rect 3471 3896 3516 3924
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3602 3884 3608 3936
rect 3660 3924 3666 3936
rect 4706 3924 4712 3936
rect 3660 3896 4712 3924
rect 3660 3884 3666 3896
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 6730 3924 6736 3936
rect 6691 3896 6736 3924
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7668 3924 7696 3964
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 13538 3992 13544 4004
rect 8067 3964 13544 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 13538 3952 13544 3964
rect 13596 3952 13602 4004
rect 8294 3924 8300 3936
rect 7668 3896 8300 3924
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8573 3927 8631 3933
rect 8573 3893 8585 3927
rect 8619 3924 8631 3927
rect 8662 3924 8668 3936
rect 8619 3896 8668 3924
rect 8619 3893 8631 3896
rect 8573 3887 8631 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 3036 3834 9844 3856
rect 3036 3782 5666 3834
rect 5718 3782 5730 3834
rect 5782 3782 5794 3834
rect 5846 3782 5858 3834
rect 5910 3782 5922 3834
rect 5974 3782 8766 3834
rect 8818 3782 8830 3834
rect 8882 3782 8894 3834
rect 8946 3782 8958 3834
rect 9010 3782 9022 3834
rect 9074 3782 9844 3834
rect 3036 3760 9844 3782
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 2924 3692 5028 3720
rect 2924 3680 2930 3692
rect 3418 3584 3424 3596
rect 3379 3556 3424 3584
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 3694 3584 3700 3596
rect 3655 3556 3700 3584
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 4890 3544 4896 3596
rect 4948 3544 4954 3596
rect 4908 3516 4936 3544
rect 4830 3488 4936 3516
rect 5000 3448 5028 3692
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5169 3723 5227 3729
rect 5169 3720 5181 3723
rect 5132 3692 5181 3720
rect 5132 3680 5138 3692
rect 5169 3689 5181 3692
rect 5215 3689 5227 3723
rect 5169 3683 5227 3689
rect 5353 3723 5411 3729
rect 5353 3689 5365 3723
rect 5399 3720 5411 3723
rect 6638 3720 6644 3732
rect 5399 3692 6644 3720
rect 5399 3689 5411 3692
rect 5353 3683 5411 3689
rect 5184 3584 5212 3683
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 8386 3720 8392 3732
rect 6788 3692 8392 3720
rect 6788 3680 6794 3692
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 8662 3720 8668 3732
rect 8623 3692 8668 3720
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 7190 3612 7196 3664
rect 7248 3652 7254 3664
rect 7248 3624 7604 3652
rect 7248 3612 7254 3624
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 5184 3556 6101 3584
rect 6089 3553 6101 3556
rect 6135 3553 6147 3587
rect 6089 3547 6147 3553
rect 6362 3544 6368 3596
rect 6420 3584 6426 3596
rect 6638 3584 6644 3596
rect 6420 3556 6644 3584
rect 6420 3544 6426 3556
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 7576 3584 7604 3624
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 8849 3655 8907 3661
rect 8849 3652 8861 3655
rect 7708 3624 8861 3652
rect 7708 3612 7714 3624
rect 8849 3621 8861 3624
rect 8895 3621 8907 3655
rect 8849 3615 8907 3621
rect 9309 3587 9367 3593
rect 9309 3584 9321 3587
rect 7576 3556 9321 3584
rect 9309 3553 9321 3556
rect 9355 3553 9367 3587
rect 9309 3547 9367 3553
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 5994 3516 6000 3528
rect 5767 3488 6000 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 5626 3448 5632 3460
rect 5000 3420 5632 3448
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 7576 3448 7604 3479
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 7800 3488 7972 3516
rect 7800 3476 7806 3488
rect 7834 3448 7840 3460
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 6730 3380 6736 3392
rect 3108 3352 6736 3380
rect 3108 3340 3114 3352
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 7208 3380 7236 3434
rect 7576 3420 7840 3448
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 7944 3448 7972 3488
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8260 3488 8309 3516
rect 8260 3476 8266 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8435 3488 8953 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 8404 3448 8432 3479
rect 7944 3420 8064 3448
rect 7926 3380 7932 3392
rect 7208 3352 7932 3380
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8036 3389 8064 3420
rect 8312 3420 8432 3448
rect 8312 3392 8340 3420
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 9125 3451 9183 3457
rect 9125 3448 9137 3451
rect 8720 3420 9137 3448
rect 8720 3408 8726 3420
rect 9125 3417 9137 3420
rect 9171 3417 9183 3451
rect 9125 3411 9183 3417
rect 8021 3383 8079 3389
rect 8021 3349 8033 3383
rect 8067 3349 8079 3383
rect 8021 3343 8079 3349
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8168 3352 8213 3380
rect 8168 3340 8174 3352
rect 8294 3340 8300 3392
rect 8352 3340 8358 3392
rect 3036 3290 9844 3312
rect 3036 3238 4116 3290
rect 4168 3238 4180 3290
rect 4232 3238 4244 3290
rect 4296 3238 4308 3290
rect 4360 3238 4372 3290
rect 4424 3238 7216 3290
rect 7268 3238 7280 3290
rect 7332 3238 7344 3290
rect 7396 3238 7408 3290
rect 7460 3238 7472 3290
rect 7524 3238 9844 3290
rect 3036 3216 9844 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 2823 3148 5488 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 4212 3080 4278 3108
rect 4212 3068 4218 3080
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3752 3012 3893 3040
rect 3752 3000 3758 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 5350 3040 5356 3052
rect 5311 3012 5356 3040
rect 3881 3003 3939 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5460 3040 5488 3148
rect 6086 3136 6092 3188
rect 6144 3176 6150 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 6144 3148 6377 3176
rect 6144 3136 6150 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 6457 3179 6515 3185
rect 6457 3145 6469 3179
rect 6503 3145 6515 3179
rect 6457 3139 6515 3145
rect 6472 3108 6500 3139
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 7377 3179 7435 3185
rect 7377 3176 7389 3179
rect 6880 3148 7389 3176
rect 6880 3136 6886 3148
rect 7377 3145 7389 3148
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8478 3176 8484 3188
rect 8343 3148 8484 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 6472 3080 7604 3108
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5460 3012 5917 3040
rect 5905 3009 5917 3012
rect 5951 3040 5963 3043
rect 6178 3040 6184 3052
rect 5951 3012 6184 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6638 3040 6644 3052
rect 6599 3012 6644 3040
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7576 3049 7604 3080
rect 7926 3068 7932 3120
rect 7984 3108 7990 3120
rect 8570 3108 8576 3120
rect 7984 3080 8576 3108
rect 7984 3068 7990 3080
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 8386 3040 8392 3052
rect 7699 3012 8392 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3040 8539 3043
rect 9490 3040 9496 3052
rect 8527 3012 9496 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 3384 2944 3525 2972
rect 3384 2932 3390 2944
rect 3513 2941 3525 2944
rect 3559 2941 3571 2975
rect 3513 2935 3571 2941
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 6270 2972 6276 2984
rect 5859 2944 6276 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 6380 2944 8677 2972
rect 6380 2904 6408 2944
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2972 8907 2975
rect 9122 2972 9128 2984
rect 8895 2944 9128 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 4816 2876 6408 2904
rect 2685 2839 2743 2845
rect 2685 2805 2697 2839
rect 2731 2836 2743 2839
rect 4816 2836 4844 2876
rect 7006 2864 7012 2916
rect 7064 2864 7070 2916
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 8478 2904 8484 2916
rect 7331 2876 8484 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 2731 2808 4844 2836
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5997 2839 6055 2845
rect 5997 2836 6009 2839
rect 5224 2808 6009 2836
rect 5224 2796 5230 2808
rect 5997 2805 6009 2808
rect 6043 2836 6055 2839
rect 6822 2836 6828 2848
rect 6043 2808 6828 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6822 2796 6828 2808
rect 6880 2836 6886 2848
rect 6917 2839 6975 2845
rect 6917 2836 6929 2839
rect 6880 2808 6929 2836
rect 6880 2796 6886 2808
rect 6917 2805 6929 2808
rect 6963 2805 6975 2839
rect 7024 2836 7052 2864
rect 7745 2839 7803 2845
rect 7745 2836 7757 2839
rect 7024 2808 7757 2836
rect 6917 2799 6975 2805
rect 7745 2805 7757 2808
rect 7791 2805 7803 2839
rect 8110 2836 8116 2848
rect 8071 2808 8116 2836
rect 7745 2799 7803 2805
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 9306 2836 9312 2848
rect 9267 2808 9312 2836
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 3036 2746 9844 2768
rect 3036 2694 5666 2746
rect 5718 2694 5730 2746
rect 5782 2694 5794 2746
rect 5846 2694 5858 2746
rect 5910 2694 5922 2746
rect 5974 2694 8766 2746
rect 8818 2694 8830 2746
rect 8882 2694 8894 2746
rect 8946 2694 8958 2746
rect 9010 2694 9022 2746
rect 9074 2694 9844 2746
rect 3036 2672 9844 2694
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 4154 2632 4160 2644
rect 3651 2604 4160 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2601 4399 2635
rect 4341 2595 4399 2601
rect 4356 2564 4384 2595
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 5592 2604 6469 2632
rect 5592 2592 5598 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6604 2604 6745 2632
rect 6604 2592 6610 2604
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 6733 2595 6791 2601
rect 7469 2635 7527 2641
rect 7469 2601 7481 2635
rect 7515 2632 7527 2635
rect 7558 2632 7564 2644
rect 7515 2604 7564 2632
rect 7515 2601 7527 2604
rect 7469 2595 7527 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8110 2592 8116 2644
rect 8168 2632 8174 2644
rect 8297 2635 8355 2641
rect 8168 2604 8248 2632
rect 8168 2592 8174 2604
rect 5166 2564 5172 2576
rect 4356 2536 5172 2564
rect 5166 2524 5172 2536
rect 5224 2524 5230 2576
rect 5261 2567 5319 2573
rect 5261 2533 5273 2567
rect 5307 2533 5319 2567
rect 5261 2527 5319 2533
rect 6273 2567 6331 2573
rect 6273 2533 6285 2567
rect 6319 2564 6331 2567
rect 8220 2564 8248 2604
rect 8297 2601 8309 2635
rect 8343 2632 8355 2635
rect 8570 2632 8576 2644
rect 8343 2604 8576 2632
rect 8343 2601 8355 2604
rect 8297 2595 8355 2601
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 9122 2632 9128 2644
rect 9083 2604 9128 2632
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 6319 2536 8156 2564
rect 8220 2536 9352 2564
rect 6319 2533 6331 2536
rect 6273 2527 6331 2533
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 3804 2468 4629 2496
rect 3510 2428 3516 2440
rect 3471 2400 3516 2428
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 3804 2437 3832 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2397 3847 2431
rect 4062 2428 4068 2440
rect 4023 2400 4068 2428
rect 3789 2391 3847 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2397 4215 2431
rect 4157 2391 4215 2397
rect 2314 2320 2320 2372
rect 2372 2360 2378 2372
rect 4172 2360 4200 2391
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 5276 2428 5304 2527
rect 6086 2456 6092 2508
rect 6144 2496 6150 2508
rect 6144 2468 6776 2496
rect 6144 2456 6150 2468
rect 5442 2428 5448 2440
rect 4396 2400 5304 2428
rect 5403 2400 5448 2428
rect 4396 2388 4402 2400
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 6178 2428 6184 2440
rect 5951 2400 6184 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 6638 2428 6644 2440
rect 6599 2400 6644 2428
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 6748 2428 6776 2468
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 8018 2496 8024 2508
rect 6880 2468 7236 2496
rect 6880 2456 6886 2468
rect 7208 2437 7236 2468
rect 7760 2468 8024 2496
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6748 2400 6929 2428
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2424 7711 2431
rect 7760 2424 7788 2468
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 7699 2397 7788 2424
rect 7653 2396 7788 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 8128 2428 8156 2536
rect 8478 2428 8484 2440
rect 7975 2400 8156 2428
rect 8439 2400 8484 2428
rect 7975 2397 7987 2400
rect 7653 2391 7711 2396
rect 7929 2391 7987 2397
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2397 8815 2431
rect 9030 2428 9036 2440
rect 8991 2400 9036 2428
rect 8757 2391 8815 2397
rect 4709 2363 4767 2369
rect 4709 2360 4721 2363
rect 2372 2332 4721 2360
rect 2372 2320 2378 2332
rect 4709 2329 4721 2332
rect 4755 2329 4767 2363
rect 4709 2323 4767 2329
rect 4893 2363 4951 2369
rect 4893 2329 4905 2363
rect 4939 2360 4951 2363
rect 5166 2360 5172 2372
rect 4939 2332 5172 2360
rect 4939 2329 4951 2332
rect 4893 2323 4951 2329
rect 5166 2320 5172 2332
rect 5224 2360 5230 2372
rect 6089 2363 6147 2369
rect 6089 2360 6101 2363
rect 5224 2332 6101 2360
rect 5224 2320 5230 2332
rect 6089 2329 6101 2332
rect 6135 2329 6147 2363
rect 6089 2323 6147 2329
rect 6730 2320 6736 2372
rect 6788 2360 6794 2372
rect 7009 2363 7067 2369
rect 7009 2360 7021 2363
rect 6788 2332 7021 2360
rect 6788 2320 6794 2332
rect 7009 2329 7021 2332
rect 7055 2329 7067 2363
rect 7009 2323 7067 2329
rect 7377 2363 7435 2369
rect 7377 2329 7389 2363
rect 7423 2360 7435 2363
rect 8772 2360 8800 2391
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 9324 2437 9352 2536
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 7423 2332 8800 2360
rect 7423 2329 7435 2332
rect 7377 2323 7435 2329
rect 3878 2292 3884 2304
rect 3839 2264 3884 2292
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 5077 2295 5135 2301
rect 5077 2261 5089 2295
rect 5123 2292 5135 2295
rect 6270 2292 6276 2304
rect 5123 2264 6276 2292
rect 5123 2261 5135 2264
rect 5077 2255 5135 2261
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 7745 2295 7803 2301
rect 7745 2292 7757 2295
rect 6512 2264 7757 2292
rect 6512 2252 6518 2264
rect 7745 2261 7757 2264
rect 7791 2261 7803 2295
rect 7745 2255 7803 2261
rect 7834 2252 7840 2304
rect 7892 2292 7898 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 7892 2264 8585 2292
rect 7892 2252 7898 2264
rect 8573 2261 8585 2264
rect 8619 2261 8631 2295
rect 8846 2292 8852 2304
rect 8807 2264 8852 2292
rect 8573 2255 8631 2261
rect 8846 2252 8852 2264
rect 8904 2252 8910 2304
rect 3036 2202 9844 2224
rect 3036 2150 4116 2202
rect 4168 2150 4180 2202
rect 4232 2150 4244 2202
rect 4296 2150 4308 2202
rect 4360 2150 4372 2202
rect 4424 2150 7216 2202
rect 7268 2150 7280 2202
rect 7332 2150 7344 2202
rect 7396 2150 7408 2202
rect 7460 2150 7472 2202
rect 7524 2150 9844 2202
rect 3036 2128 9844 2150
rect 3878 2048 3884 2100
rect 3936 2088 3942 2100
rect 5994 2088 6000 2100
rect 3936 2060 6000 2088
rect 3936 2048 3942 2060
rect 5994 2048 6000 2060
rect 6052 2048 6058 2100
rect 6270 2048 6276 2100
rect 6328 2088 6334 2100
rect 9030 2088 9036 2100
rect 6328 2060 9036 2088
rect 6328 2048 6334 2060
rect 9030 2048 9036 2060
rect 9088 2048 9094 2100
rect 5350 1980 5356 2032
rect 5408 2020 5414 2032
rect 8846 2020 8852 2032
rect 5408 1992 8852 2020
rect 5408 1980 5414 1992
rect 8846 1980 8852 1992
rect 8904 1980 8910 2032
<< via1 >>
rect 1860 11908 1912 11960
rect 8116 11908 8168 11960
rect 2412 11840 2464 11892
rect 6644 11840 6696 11892
rect 3148 11772 3200 11824
rect 4068 11772 4120 11824
rect 7380 11704 7432 11756
rect 9496 11704 9548 11756
rect 2136 11636 2188 11688
rect 4344 11636 4396 11688
rect 2320 11568 2372 11620
rect 3608 11568 3660 11620
rect 3700 11568 3752 11620
rect 6736 11636 6788 11688
rect 7472 11636 7524 11688
rect 9772 11636 9824 11688
rect 6184 11568 6236 11620
rect 7656 11568 7708 11620
rect 2964 11500 3016 11552
rect 6828 11500 6880 11552
rect 7564 11500 7616 11552
rect 13360 11500 13412 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 5666 11398 5718 11450
rect 5730 11398 5782 11450
rect 5794 11398 5846 11450
rect 5858 11398 5910 11450
rect 5922 11398 5974 11450
rect 8766 11398 8818 11450
rect 8830 11398 8882 11450
rect 8894 11398 8946 11450
rect 8958 11398 9010 11450
rect 9022 11398 9074 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2228 11339 2280 11348
rect 2228 11305 2237 11339
rect 2237 11305 2271 11339
rect 2271 11305 2280 11339
rect 2228 11296 2280 11305
rect 2964 11296 3016 11348
rect 3976 11296 4028 11348
rect 4620 11296 4672 11348
rect 4804 11339 4856 11348
rect 4804 11305 4813 11339
rect 4813 11305 4847 11339
rect 4847 11305 4856 11339
rect 4804 11296 4856 11305
rect 7012 11296 7064 11348
rect 7288 11296 7340 11348
rect 7748 11296 7800 11348
rect 2228 11092 2280 11144
rect 2412 11092 2464 11144
rect 2780 11228 2832 11280
rect 2964 11092 3016 11144
rect 5632 11160 5684 11212
rect 3240 11092 3292 11144
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 3700 11092 3752 11144
rect 4068 11092 4120 11144
rect 4344 11092 4396 11144
rect 4712 11092 4764 11144
rect 5540 11092 5592 11144
rect 6828 11160 6880 11212
rect 6000 11092 6052 11144
rect 6460 11092 6512 11144
rect 7104 11160 7156 11212
rect 7196 11160 7248 11212
rect 13728 11296 13780 11348
rect 13820 11228 13872 11280
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 2596 10956 2648 11008
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 5264 11024 5316 11076
rect 3332 10956 3384 11008
rect 3976 10956 4028 11008
rect 5080 10956 5132 11008
rect 5172 10956 5224 11008
rect 6276 11024 6328 11076
rect 6092 10956 6144 11008
rect 6368 10999 6420 11008
rect 6368 10965 6377 10999
rect 6377 10965 6411 10999
rect 6411 10965 6420 10999
rect 6368 10956 6420 10965
rect 7196 11024 7248 11076
rect 7472 11092 7524 11144
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 13452 11160 13504 11212
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 8392 11092 8444 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 7564 10956 7616 11008
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 8576 10956 8628 11008
rect 16672 10956 16724 11008
rect 4116 10854 4168 10906
rect 4180 10854 4232 10906
rect 4244 10854 4296 10906
rect 4308 10854 4360 10906
rect 4372 10854 4424 10906
rect 7216 10854 7268 10906
rect 7280 10854 7332 10906
rect 7344 10854 7396 10906
rect 7408 10854 7460 10906
rect 7472 10854 7524 10906
rect 1216 10795 1268 10804
rect 1216 10761 1225 10795
rect 1225 10761 1259 10795
rect 1259 10761 1268 10795
rect 1216 10752 1268 10761
rect 2044 10795 2096 10804
rect 2044 10761 2053 10795
rect 2053 10761 2087 10795
rect 2087 10761 2096 10795
rect 2044 10752 2096 10761
rect 3976 10752 4028 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 2688 10684 2740 10736
rect 3424 10684 3476 10736
rect 4068 10684 4120 10736
rect 5172 10752 5224 10804
rect 4436 10684 4488 10736
rect 4804 10684 4856 10736
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 4528 10591 4580 10600
rect 4528 10557 4537 10591
rect 4537 10557 4571 10591
rect 4571 10557 4580 10591
rect 4528 10548 4580 10557
rect 4620 10548 4672 10600
rect 6920 10684 6972 10736
rect 9220 10752 9272 10804
rect 5908 10616 5960 10668
rect 8116 10659 8168 10668
rect 8116 10625 8125 10659
rect 8125 10625 8159 10659
rect 8159 10625 8168 10659
rect 8116 10616 8168 10625
rect 8668 10548 8720 10600
rect 4068 10412 4120 10464
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 9312 10480 9364 10532
rect 4160 10412 4212 10421
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 5666 10310 5718 10362
rect 5730 10310 5782 10362
rect 5794 10310 5846 10362
rect 5858 10310 5910 10362
rect 5922 10310 5974 10362
rect 8766 10310 8818 10362
rect 8830 10310 8882 10362
rect 8894 10310 8946 10362
rect 8958 10310 9010 10362
rect 9022 10310 9074 10362
rect 1952 10208 2004 10260
rect 2136 10251 2188 10260
rect 2136 10217 2145 10251
rect 2145 10217 2179 10251
rect 2179 10217 2188 10251
rect 2136 10208 2188 10217
rect 3516 10208 3568 10260
rect 1860 10140 1912 10192
rect 2964 10183 3016 10192
rect 2964 10149 2973 10183
rect 2973 10149 3007 10183
rect 3007 10149 3016 10183
rect 2964 10140 3016 10149
rect 1952 10004 2004 10056
rect 2504 10004 2556 10056
rect 3976 10072 4028 10124
rect 3056 10004 3108 10056
rect 1768 9936 1820 9988
rect 2228 9868 2280 9920
rect 3700 10004 3752 10056
rect 5908 10140 5960 10192
rect 6828 10140 6880 10192
rect 7012 10140 7064 10192
rect 7196 10140 7248 10192
rect 8300 10208 8352 10260
rect 8024 10140 8076 10192
rect 9312 10115 9364 10124
rect 9312 10081 9321 10115
rect 9321 10081 9355 10115
rect 9355 10081 9364 10115
rect 9312 10072 9364 10081
rect 4528 10004 4580 10056
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 3792 9936 3844 9988
rect 5540 9936 5592 9988
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 3608 9868 3660 9920
rect 6552 10004 6604 10056
rect 7472 10047 7524 10056
rect 7012 9979 7064 9988
rect 7012 9945 7021 9979
rect 7021 9945 7055 9979
rect 7055 9945 7064 9979
rect 7012 9936 7064 9945
rect 7196 9979 7248 9988
rect 7196 9945 7205 9979
rect 7205 9945 7239 9979
rect 7239 9945 7248 9979
rect 7196 9936 7248 9945
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 8024 9979 8076 9988
rect 8024 9945 8033 9979
rect 8033 9945 8067 9979
rect 8067 9945 8076 9979
rect 8024 9936 8076 9945
rect 8116 9936 8168 9988
rect 9220 9979 9272 9988
rect 9220 9945 9229 9979
rect 9229 9945 9263 9979
rect 9263 9945 9272 9979
rect 9220 9936 9272 9945
rect 6644 9868 6696 9920
rect 4116 9766 4168 9818
rect 4180 9766 4232 9818
rect 4244 9766 4296 9818
rect 4308 9766 4360 9818
rect 4372 9766 4424 9818
rect 7216 9766 7268 9818
rect 7280 9766 7332 9818
rect 7344 9766 7396 9818
rect 7408 9766 7460 9818
rect 7472 9766 7524 9818
rect 2320 9639 2372 9648
rect 2320 9605 2329 9639
rect 2329 9605 2363 9639
rect 2363 9605 2372 9639
rect 2320 9596 2372 9605
rect 3148 9664 3200 9716
rect 2228 9528 2280 9580
rect 4436 9596 4488 9648
rect 5540 9664 5592 9716
rect 7564 9664 7616 9716
rect 8116 9664 8168 9716
rect 2044 9460 2096 9512
rect 2964 9528 3016 9580
rect 3240 9460 3292 9512
rect 3884 9528 3936 9580
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 1952 9392 2004 9444
rect 4712 9460 4764 9512
rect 3332 9324 3384 9376
rect 4528 9324 4580 9376
rect 5080 9324 5132 9376
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 6276 9528 6328 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7932 9528 7984 9580
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 7012 9460 7064 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 8024 9460 8076 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 6736 9392 6788 9444
rect 6000 9324 6052 9376
rect 6920 9324 6972 9376
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 7656 9324 7708 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 5666 9222 5718 9274
rect 5730 9222 5782 9274
rect 5794 9222 5846 9274
rect 5858 9222 5910 9274
rect 5922 9222 5974 9274
rect 8766 9222 8818 9274
rect 8830 9222 8882 9274
rect 8894 9222 8946 9274
rect 8958 9222 9010 9274
rect 9022 9222 9074 9274
rect 1768 9163 1820 9172
rect 1768 9129 1777 9163
rect 1777 9129 1811 9163
rect 1811 9129 1820 9163
rect 1768 9120 1820 9129
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 2320 9052 2372 9104
rect 4436 9120 4488 9172
rect 4988 9120 5040 9172
rect 5448 9120 5500 9172
rect 2504 8984 2556 9036
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 3148 8959 3200 8968
rect 2780 8848 2832 8900
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 5172 8984 5224 9036
rect 6736 9052 6788 9104
rect 7472 9052 7524 9104
rect 13636 9052 13688 9104
rect 6092 8984 6144 9036
rect 8576 8984 8628 9036
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 8024 8916 8076 8968
rect 3884 8891 3936 8900
rect 1308 8780 1360 8832
rect 1400 8780 1452 8832
rect 1952 8780 2004 8832
rect 3240 8823 3292 8832
rect 3240 8789 3249 8823
rect 3249 8789 3283 8823
rect 3283 8789 3292 8823
rect 3240 8780 3292 8789
rect 3884 8857 3893 8891
rect 3893 8857 3927 8891
rect 3927 8857 3936 8891
rect 3884 8848 3936 8857
rect 4896 8848 4948 8900
rect 5172 8848 5224 8900
rect 5816 8780 5868 8832
rect 6000 8848 6052 8900
rect 8300 8916 8352 8968
rect 9404 8916 9456 8968
rect 8576 8848 8628 8900
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 13544 8780 13596 8832
rect 4116 8678 4168 8730
rect 4180 8678 4232 8730
rect 4244 8678 4296 8730
rect 4308 8678 4360 8730
rect 4372 8678 4424 8730
rect 7216 8678 7268 8730
rect 7280 8678 7332 8730
rect 7344 8678 7396 8730
rect 7408 8678 7460 8730
rect 7472 8678 7524 8730
rect 1860 8576 1912 8628
rect 3792 8576 3844 8628
rect 3884 8576 3936 8628
rect 4712 8576 4764 8628
rect 5816 8619 5868 8628
rect 5816 8585 5825 8619
rect 5825 8585 5859 8619
rect 5859 8585 5868 8619
rect 5816 8576 5868 8585
rect 8208 8576 8260 8628
rect 9496 8619 9548 8628
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 2228 8551 2280 8560
rect 2228 8517 2237 8551
rect 2237 8517 2271 8551
rect 2271 8517 2280 8551
rect 2228 8508 2280 8517
rect 1492 8440 1544 8492
rect 2964 8508 3016 8560
rect 3332 8508 3384 8560
rect 2044 8372 2096 8424
rect 1584 8304 1636 8356
rect 2504 8372 2556 8424
rect 7104 8508 7156 8560
rect 9220 8508 9272 8560
rect 4344 8440 4396 8492
rect 6276 8440 6328 8492
rect 4528 8372 4580 8424
rect 6460 8483 6512 8492
rect 6460 8449 6469 8483
rect 6469 8449 6503 8483
rect 6503 8449 6512 8483
rect 6460 8440 6512 8449
rect 9312 8440 9364 8492
rect 13728 8440 13780 8492
rect 22468 8440 22520 8492
rect 5540 8304 5592 8356
rect 6736 8372 6788 8424
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 8116 8372 8168 8424
rect 13820 8372 13872 8424
rect 22192 8372 22244 8424
rect 6552 8304 6604 8356
rect 6828 8304 6880 8356
rect 4896 8236 4948 8288
rect 5356 8236 5408 8288
rect 6000 8236 6052 8288
rect 22744 8236 22796 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 5666 8134 5718 8186
rect 5730 8134 5782 8186
rect 5794 8134 5846 8186
rect 5858 8134 5910 8186
rect 5922 8134 5974 8186
rect 8766 8134 8818 8186
rect 8830 8134 8882 8186
rect 8894 8134 8946 8186
rect 8958 8134 9010 8186
rect 9022 8134 9074 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 1768 7964 1820 8016
rect 1216 7896 1268 7948
rect 2136 7964 2188 8016
rect 2412 7964 2464 8016
rect 6000 8032 6052 8084
rect 6460 8075 6512 8084
rect 6460 8041 6469 8075
rect 6469 8041 6503 8075
rect 6503 8041 6512 8075
rect 6460 8032 6512 8041
rect 7196 8032 7248 8084
rect 4712 7964 4764 8016
rect 7932 7964 7984 8016
rect 8116 7964 8168 8016
rect 8300 8007 8352 8016
rect 8300 7973 8309 8007
rect 8309 7973 8343 8007
rect 8343 7973 8352 8007
rect 8300 7964 8352 7973
rect 3056 7939 3108 7948
rect 3056 7905 3065 7939
rect 3065 7905 3099 7939
rect 3099 7905 3108 7939
rect 3056 7896 3108 7905
rect 3240 7896 3292 7948
rect 5080 7896 5132 7948
rect 5448 7896 5500 7948
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 6920 7896 6972 7948
rect 9220 8032 9272 8084
rect 13452 7964 13504 8016
rect 22284 7964 22336 8016
rect 4068 7828 4120 7880
rect 8208 7828 8260 7880
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 3516 7760 3568 7812
rect 3884 7760 3936 7812
rect 4252 7760 4304 7812
rect 1124 7692 1176 7744
rect 2136 7692 2188 7744
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 2780 7692 2832 7701
rect 3056 7735 3108 7744
rect 3056 7701 3065 7735
rect 3065 7701 3099 7735
rect 3099 7701 3108 7735
rect 3056 7692 3108 7701
rect 3240 7692 3292 7744
rect 5080 7760 5132 7812
rect 5448 7760 5500 7812
rect 6920 7760 6972 7812
rect 7104 7760 7156 7812
rect 4528 7692 4580 7744
rect 4620 7692 4672 7744
rect 22376 7896 22428 7948
rect 4116 7590 4168 7642
rect 4180 7590 4232 7642
rect 4244 7590 4296 7642
rect 4308 7590 4360 7642
rect 4372 7590 4424 7642
rect 7216 7590 7268 7642
rect 7280 7590 7332 7642
rect 7344 7590 7396 7642
rect 7408 7590 7460 7642
rect 7472 7590 7524 7642
rect 2504 7420 2556 7472
rect 1676 7352 1728 7404
rect 1952 7352 2004 7404
rect 4620 7420 4672 7472
rect 5356 7420 5408 7472
rect 8024 7488 8076 7540
rect 9312 7531 9364 7540
rect 1032 7216 1084 7268
rect 3240 7352 3292 7404
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 3516 7352 3568 7404
rect 3976 7352 4028 7404
rect 6460 7352 6512 7404
rect 7840 7352 7892 7404
rect 3792 7259 3844 7268
rect 3792 7225 3801 7259
rect 3801 7225 3835 7259
rect 3835 7225 3844 7259
rect 3792 7216 3844 7225
rect 1216 7148 1268 7200
rect 1400 7148 1452 7200
rect 1676 7148 1728 7200
rect 2044 7148 2096 7200
rect 2136 7191 2188 7200
rect 2136 7157 2145 7191
rect 2145 7157 2179 7191
rect 2179 7157 2188 7191
rect 2136 7148 2188 7157
rect 2412 7148 2464 7200
rect 3884 7148 3936 7200
rect 5540 7284 5592 7336
rect 6828 7284 6880 7336
rect 5448 7216 5500 7268
rect 9312 7497 9321 7531
rect 9321 7497 9355 7531
rect 9355 7497 9364 7531
rect 9312 7488 9364 7497
rect 9128 7352 9180 7404
rect 8208 7216 8260 7268
rect 9588 7148 9640 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 5666 7046 5718 7098
rect 5730 7046 5782 7098
rect 5794 7046 5846 7098
rect 5858 7046 5910 7098
rect 5922 7046 5974 7098
rect 8766 7046 8818 7098
rect 8830 7046 8882 7098
rect 8894 7046 8946 7098
rect 8958 7046 9010 7098
rect 9022 7046 9074 7098
rect 1584 6944 1636 6996
rect 3240 6944 3292 6996
rect 3884 6944 3936 6996
rect 7104 6944 7156 6996
rect 7748 6944 7800 6996
rect 13820 7080 13872 7132
rect 19800 7080 19852 7132
rect 13636 6944 13688 6996
rect 9588 6876 9640 6928
rect 3884 6808 3936 6860
rect 6184 6808 6236 6860
rect 6460 6808 6512 6860
rect 9312 6851 9364 6860
rect 9312 6817 9321 6851
rect 9321 6817 9355 6851
rect 9355 6817 9364 6851
rect 9312 6808 9364 6817
rect 3240 6740 3292 6792
rect 3792 6740 3844 6792
rect 1400 6647 1452 6656
rect 1400 6613 1409 6647
rect 1409 6613 1443 6647
rect 1443 6613 1452 6647
rect 1400 6604 1452 6613
rect 1860 6672 1912 6724
rect 2596 6604 2648 6656
rect 5080 6672 5132 6724
rect 3240 6604 3292 6656
rect 3792 6604 3844 6656
rect 3884 6604 3936 6656
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8300 6740 8352 6792
rect 8392 6740 8444 6792
rect 8852 6740 8904 6792
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 22100 6672 22152 6724
rect 5264 6604 5316 6656
rect 8024 6604 8076 6656
rect 8668 6604 8720 6656
rect 8852 6604 8904 6656
rect 4116 6502 4168 6554
rect 4180 6502 4232 6554
rect 4244 6502 4296 6554
rect 4308 6502 4360 6554
rect 4372 6502 4424 6554
rect 7216 6502 7268 6554
rect 7280 6502 7332 6554
rect 7344 6502 7396 6554
rect 7408 6502 7460 6554
rect 7472 6502 7524 6554
rect 2136 6400 2188 6452
rect 1308 6332 1360 6384
rect 2872 6332 2924 6384
rect 5264 6400 5316 6452
rect 8392 6400 8444 6452
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 3976 6332 4028 6384
rect 6276 6332 6328 6384
rect 7656 6332 7708 6384
rect 1216 6264 1268 6316
rect 3148 6264 3200 6316
rect 3240 6196 3292 6248
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4528 6307 4580 6316
rect 4160 6264 4212 6273
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 6000 6307 6052 6316
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 4896 6196 4948 6248
rect 1400 6128 1452 6180
rect 3608 6060 3660 6112
rect 3884 6060 3936 6112
rect 4160 6128 4212 6180
rect 8208 6264 8260 6316
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 6736 6196 6788 6248
rect 7012 6196 7064 6248
rect 8668 6264 8720 6316
rect 8300 6128 8352 6180
rect 7748 6103 7800 6112
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 7932 6060 7984 6069
rect 9220 6196 9272 6248
rect 13820 6128 13872 6180
rect 9312 6060 9364 6112
rect 5666 5958 5718 6010
rect 5730 5958 5782 6010
rect 5794 5958 5846 6010
rect 5858 5958 5910 6010
rect 5922 5958 5974 6010
rect 8766 5958 8818 6010
rect 8830 5958 8882 6010
rect 8894 5958 8946 6010
rect 8958 5958 9010 6010
rect 9022 5958 9074 6010
rect 3792 5856 3844 5908
rect 4896 5856 4948 5908
rect 1768 5720 1820 5772
rect 3976 5720 4028 5772
rect 1676 5652 1728 5704
rect 3056 5652 3108 5704
rect 5264 5720 5316 5772
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 8668 5899 8720 5908
rect 8668 5865 8677 5899
rect 8677 5865 8711 5899
rect 8711 5865 8720 5899
rect 8668 5856 8720 5865
rect 9404 5856 9456 5908
rect 5448 5788 5500 5840
rect 6184 5763 6236 5772
rect 5172 5695 5224 5704
rect 5172 5661 5181 5695
rect 5181 5661 5215 5695
rect 5215 5661 5224 5695
rect 5172 5652 5224 5661
rect 6184 5729 6193 5763
rect 6193 5729 6227 5763
rect 6227 5729 6236 5763
rect 6184 5720 6236 5729
rect 8208 5788 8260 5840
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 1492 5584 1544 5636
rect 4988 5584 5040 5636
rect 3700 5516 3752 5568
rect 6368 5584 6420 5636
rect 7564 5584 7616 5636
rect 8944 5584 8996 5636
rect 4116 5414 4168 5466
rect 4180 5414 4232 5466
rect 4244 5414 4296 5466
rect 4308 5414 4360 5466
rect 4372 5414 4424 5466
rect 7216 5414 7268 5466
rect 7280 5414 7332 5466
rect 7344 5414 7396 5466
rect 7408 5414 7460 5466
rect 7472 5414 7524 5466
rect 6184 5312 6236 5364
rect 7840 5312 7892 5364
rect 8668 5312 8720 5364
rect 8944 5312 8996 5364
rect 5264 5244 5316 5296
rect 7104 5244 7156 5296
rect 8392 5244 8444 5296
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 5540 5108 5592 5160
rect 5632 5108 5684 5160
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 8576 5176 8628 5228
rect 6736 5108 6788 5160
rect 5264 5040 5316 5092
rect 5908 5040 5960 5092
rect 13728 5040 13780 5092
rect 4988 4972 5040 5024
rect 7840 4972 7892 5024
rect 9404 4972 9456 5024
rect 9496 5015 9548 5024
rect 9496 4981 9505 5015
rect 9505 4981 9539 5015
rect 9539 4981 9548 5015
rect 9496 4972 9548 4981
rect 5666 4870 5718 4922
rect 5730 4870 5782 4922
rect 5794 4870 5846 4922
rect 5858 4870 5910 4922
rect 5922 4870 5974 4922
rect 8766 4870 8818 4922
rect 8830 4870 8882 4922
rect 8894 4870 8946 4922
rect 8958 4870 9010 4922
rect 9022 4870 9074 4922
rect 3332 4700 3384 4752
rect 5264 4768 5316 4820
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 5172 4700 5224 4752
rect 6000 4768 6052 4820
rect 9220 4768 9272 4820
rect 6460 4700 6512 4752
rect 5080 4632 5132 4684
rect 3240 4564 3292 4616
rect 5540 4632 5592 4684
rect 2688 4496 2740 4548
rect 3424 4496 3476 4548
rect 3976 4496 4028 4548
rect 5632 4564 5684 4616
rect 6368 4564 6420 4616
rect 6736 4564 6788 4616
rect 8576 4564 8628 4616
rect 8300 4496 8352 4548
rect 6552 4428 6604 4480
rect 4116 4326 4168 4378
rect 4180 4326 4232 4378
rect 4244 4326 4296 4378
rect 4308 4326 4360 4378
rect 4372 4326 4424 4378
rect 7216 4326 7268 4378
rect 7280 4326 7332 4378
rect 7344 4326 7396 4378
rect 7408 4326 7460 4378
rect 7472 4326 7524 4378
rect 6092 4224 6144 4276
rect 7104 4224 7156 4276
rect 7656 4224 7708 4276
rect 3240 4156 3292 4208
rect 3884 4156 3936 4208
rect 3516 4088 3568 4140
rect 6552 4156 6604 4208
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 6460 4088 6512 4140
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 5448 4020 5500 4072
rect 6368 4020 6420 4072
rect 6736 4020 6788 4072
rect 8576 4156 8628 4208
rect 7656 4088 7708 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 8208 4088 8260 4140
rect 8392 4088 8444 4140
rect 9312 4088 9364 4140
rect 9404 4088 9456 4140
rect 9128 4020 9180 4072
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 3608 3884 3660 3936
rect 4712 3884 4764 3936
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 13544 3952 13596 4004
rect 8300 3884 8352 3936
rect 8668 3884 8720 3936
rect 5666 3782 5718 3834
rect 5730 3782 5782 3834
rect 5794 3782 5846 3834
rect 5858 3782 5910 3834
rect 5922 3782 5974 3834
rect 8766 3782 8818 3834
rect 8830 3782 8882 3834
rect 8894 3782 8946 3834
rect 8958 3782 9010 3834
rect 9022 3782 9074 3834
rect 2872 3680 2924 3732
rect 3424 3587 3476 3596
rect 3424 3553 3433 3587
rect 3433 3553 3467 3587
rect 3467 3553 3476 3587
rect 3424 3544 3476 3553
rect 3700 3587 3752 3596
rect 3700 3553 3709 3587
rect 3709 3553 3743 3587
rect 3743 3553 3752 3587
rect 3700 3544 3752 3553
rect 4896 3544 4948 3596
rect 5080 3680 5132 3732
rect 6644 3680 6696 3732
rect 6736 3680 6788 3732
rect 8392 3680 8444 3732
rect 8668 3723 8720 3732
rect 8668 3689 8677 3723
rect 8677 3689 8711 3723
rect 8711 3689 8720 3723
rect 8668 3680 8720 3689
rect 7196 3612 7248 3664
rect 6368 3544 6420 3596
rect 6644 3544 6696 3596
rect 7656 3612 7708 3664
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 6000 3476 6052 3528
rect 5632 3408 5684 3460
rect 7748 3476 7800 3528
rect 3056 3340 3108 3392
rect 6736 3340 6788 3392
rect 7840 3408 7892 3460
rect 8208 3476 8260 3528
rect 7932 3340 7984 3392
rect 8668 3408 8720 3460
rect 8116 3383 8168 3392
rect 8116 3349 8125 3383
rect 8125 3349 8159 3383
rect 8159 3349 8168 3383
rect 8116 3340 8168 3349
rect 8300 3340 8352 3392
rect 4116 3238 4168 3290
rect 4180 3238 4232 3290
rect 4244 3238 4296 3290
rect 4308 3238 4360 3290
rect 4372 3238 4424 3290
rect 7216 3238 7268 3290
rect 7280 3238 7332 3290
rect 7344 3238 7396 3290
rect 7408 3238 7460 3290
rect 7472 3238 7524 3290
rect 4160 3068 4212 3120
rect 3700 3000 3752 3052
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 6092 3136 6144 3188
rect 6828 3136 6880 3188
rect 8484 3136 8536 3188
rect 6184 3000 6236 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 6736 3000 6788 3052
rect 7932 3068 7984 3120
rect 8576 3068 8628 3120
rect 8392 3000 8444 3052
rect 9496 3000 9548 3052
rect 3332 2932 3384 2984
rect 6276 2932 6328 2984
rect 9128 2932 9180 2984
rect 7012 2864 7064 2916
rect 8484 2864 8536 2916
rect 5172 2796 5224 2848
rect 6828 2796 6880 2848
rect 8116 2839 8168 2848
rect 8116 2805 8125 2839
rect 8125 2805 8159 2839
rect 8159 2805 8168 2839
rect 8116 2796 8168 2805
rect 9312 2839 9364 2848
rect 9312 2805 9321 2839
rect 9321 2805 9355 2839
rect 9355 2805 9364 2839
rect 9312 2796 9364 2805
rect 5666 2694 5718 2746
rect 5730 2694 5782 2746
rect 5794 2694 5846 2746
rect 5858 2694 5910 2746
rect 5922 2694 5974 2746
rect 8766 2694 8818 2746
rect 8830 2694 8882 2746
rect 8894 2694 8946 2746
rect 8958 2694 9010 2746
rect 9022 2694 9074 2746
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 4160 2592 4212 2644
rect 5540 2592 5592 2644
rect 6552 2592 6604 2644
rect 7564 2592 7616 2644
rect 8116 2592 8168 2644
rect 5172 2524 5224 2576
rect 8576 2592 8628 2644
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 2320 2320 2372 2372
rect 4344 2388 4396 2440
rect 6092 2456 6144 2508
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6184 2388 6236 2440
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 6828 2456 6880 2508
rect 8024 2456 8076 2508
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 9036 2431 9088 2440
rect 5172 2320 5224 2372
rect 6736 2320 6788 2372
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 3884 2295 3936 2304
rect 3884 2261 3893 2295
rect 3893 2261 3927 2295
rect 3927 2261 3936 2295
rect 3884 2252 3936 2261
rect 6276 2252 6328 2304
rect 6460 2252 6512 2304
rect 7840 2252 7892 2304
rect 8852 2295 8904 2304
rect 8852 2261 8861 2295
rect 8861 2261 8895 2295
rect 8895 2261 8904 2295
rect 8852 2252 8904 2261
rect 4116 2150 4168 2202
rect 4180 2150 4232 2202
rect 4244 2150 4296 2202
rect 4308 2150 4360 2202
rect 4372 2150 4424 2202
rect 7216 2150 7268 2202
rect 7280 2150 7332 2202
rect 7344 2150 7396 2202
rect 7408 2150 7460 2202
rect 7472 2150 7524 2202
rect 3884 2048 3936 2100
rect 6000 2048 6052 2100
rect 6276 2048 6328 2100
rect 9036 2048 9088 2100
rect 5356 1980 5408 2032
rect 8852 1980 8904 2032
<< metal2 >>
rect 2042 13832 2098 13841
rect 2042 13767 2098 13776
rect 1950 12472 2006 12481
rect 1950 12407 2006 12416
rect 1860 11960 1912 11966
rect 1860 11902 1912 11908
rect 1674 11656 1730 11665
rect 1674 11591 1730 11600
rect 1688 11354 1716 11591
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1214 11112 1270 11121
rect 1214 11047 1270 11056
rect 1228 10810 1256 11047
rect 1216 10804 1268 10810
rect 1216 10746 1268 10752
rect 1398 10704 1454 10713
rect 1398 10639 1400 10648
rect 1452 10639 1454 10648
rect 1400 10610 1452 10616
rect 1872 10198 1900 11902
rect 1964 10266 1992 12407
rect 2056 10810 2084 13767
rect 16670 13560 16726 13569
rect 16670 13495 16726 13504
rect 3974 13152 4030 13161
rect 3974 13087 4030 13096
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2226 11792 2282 11801
rect 2226 11727 2282 11736
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2148 10266 2176 11630
rect 2240 11354 2268 11727
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2240 11150 2268 11290
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 1860 10192 1912 10198
rect 1860 10134 1912 10140
rect 1964 10062 1992 10202
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1780 9178 1808 9930
rect 2240 9926 2268 9957
rect 2228 9920 2280 9926
rect 2332 9874 2360 11562
rect 2424 11150 2452 11834
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2976 11354 3004 11494
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2780 11280 2832 11286
rect 2686 11248 2742 11257
rect 2780 11222 2832 11228
rect 2686 11183 2742 11192
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2596 11008 2648 11014
rect 2700 10996 2728 11183
rect 2648 10968 2728 10996
rect 2596 10950 2648 10956
rect 2700 10742 2728 10968
rect 2688 10736 2740 10742
rect 2792 10713 2820 11222
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2976 11014 3004 11086
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 3054 10840 3110 10849
rect 3054 10775 3110 10784
rect 2688 10678 2740 10684
rect 2778 10704 2834 10713
rect 2778 10639 2834 10648
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2280 9868 2360 9874
rect 2228 9862 2360 9868
rect 2240 9846 2360 9862
rect 2240 9586 2268 9846
rect 2318 9752 2374 9761
rect 2318 9687 2374 9696
rect 2332 9654 2360 9687
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2134 9480 2190 9489
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1964 8974 1992 9386
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1308 8832 1360 8838
rect 1308 8774 1360 8780
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1952 8832 2004 8838
rect 2056 8820 2084 9454
rect 2134 9415 2190 9424
rect 2004 8792 2084 8820
rect 1952 8774 2004 8780
rect 1216 7948 1268 7954
rect 1216 7890 1268 7896
rect 1124 7744 1176 7750
rect 1228 7721 1256 7890
rect 1124 7686 1176 7692
rect 1214 7712 1270 7721
rect 1032 7268 1084 7274
rect 1032 7210 1084 7216
rect 1044 5953 1072 7210
rect 1136 6769 1164 7686
rect 1214 7647 1270 7656
rect 1216 7200 1268 7206
rect 1216 7142 1268 7148
rect 1122 6760 1178 6769
rect 1122 6695 1178 6704
rect 1228 6322 1256 7142
rect 1320 6390 1348 8774
rect 1412 7206 1440 8774
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1308 6384 1360 6390
rect 1308 6326 1360 6332
rect 1216 6316 1268 6322
rect 1216 6258 1268 6264
rect 1412 6186 1440 6598
rect 1400 6180 1452 6186
rect 1400 6122 1452 6128
rect 1030 5944 1086 5953
rect 1030 5879 1086 5888
rect 1504 5642 1532 8434
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 7002 1624 8298
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1688 7857 1716 8026
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 1674 7848 1730 7857
rect 1674 7783 1730 7792
rect 1674 7576 1730 7585
rect 1674 7511 1730 7520
rect 1688 7410 1716 7511
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1688 5710 1716 7142
rect 1780 5778 1808 7958
rect 1872 7449 1900 8570
rect 1964 7732 1992 8774
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2056 7834 2084 8366
rect 2148 8022 2176 9415
rect 2332 9110 2360 9590
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2424 9024 2452 10542
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2964 10192 3016 10198
rect 2502 10160 2558 10169
rect 2502 10095 2558 10104
rect 2870 10160 2926 10169
rect 2964 10134 3016 10140
rect 2870 10095 2926 10104
rect 2516 10062 2544 10095
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2884 9625 2912 10095
rect 2976 9674 3004 10134
rect 3068 10062 3096 10775
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3160 9722 3188 11766
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3422 11520 3478 11529
rect 3422 11455 3478 11464
rect 3436 11150 3464 11455
rect 3514 11384 3570 11393
rect 3514 11319 3570 11328
rect 3240 11144 3292 11150
rect 3424 11144 3476 11150
rect 3292 11104 3372 11132
rect 3240 11086 3292 11092
rect 3344 11014 3372 11104
rect 3424 11086 3476 11092
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3238 10024 3294 10033
rect 3238 9959 3294 9968
rect 3252 9926 3280 9959
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3148 9716 3200 9722
rect 2976 9646 3096 9674
rect 3148 9658 3200 9664
rect 2870 9616 2926 9625
rect 2870 9551 2926 9560
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2976 9178 3004 9522
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2504 9036 2556 9042
rect 2424 8996 2504 9024
rect 2504 8978 2556 8984
rect 2318 8936 2374 8945
rect 2318 8871 2374 8880
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2240 8401 2268 8502
rect 2226 8392 2282 8401
rect 2226 8327 2282 8336
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2332 7868 2360 8871
rect 2516 8430 2544 8978
rect 2596 8968 2648 8974
rect 2594 8936 2596 8945
rect 2648 8936 2650 8945
rect 2594 8871 2650 8880
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2792 8537 2820 8842
rect 2964 8560 3016 8566
rect 2778 8528 2834 8537
rect 2964 8502 3016 8508
rect 2778 8463 2834 8472
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 2412 8016 2464 8022
rect 2410 7984 2412 7993
rect 2976 8004 3004 8502
rect 2464 7984 2466 7993
rect 2410 7919 2466 7928
rect 2792 7976 3004 8004
rect 2792 7936 2820 7976
rect 3068 7954 3096 9646
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 8968 3200 8974
rect 3252 8956 3280 9454
rect 3344 9382 3372 10950
rect 3422 10840 3478 10849
rect 3422 10775 3478 10784
rect 3436 10742 3464 10775
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 9217 3372 9318
rect 3330 9208 3386 9217
rect 3330 9143 3386 9152
rect 3436 9092 3464 10678
rect 3528 10266 3556 11319
rect 3620 11150 3648 11562
rect 3712 11150 3740 11562
rect 3988 11354 4016 13087
rect 4618 12880 4674 12889
rect 4618 12815 4674 12824
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4080 11150 4108 11766
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4526 11656 4582 11665
rect 4356 11150 4384 11630
rect 4526 11591 4582 11600
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10810 4016 10950
rect 4116 10908 4424 10928
rect 4116 10906 4122 10908
rect 4178 10906 4202 10908
rect 4258 10906 4282 10908
rect 4338 10906 4362 10908
rect 4418 10906 4424 10908
rect 4178 10854 4180 10906
rect 4360 10854 4362 10906
rect 4116 10852 4122 10854
rect 4178 10852 4202 10854
rect 4258 10852 4282 10854
rect 4338 10852 4362 10854
rect 4418 10852 4424 10854
rect 4116 10832 4424 10852
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4068 10736 4120 10742
rect 4436 10736 4488 10742
rect 4120 10696 4436 10724
rect 4068 10678 4120 10684
rect 4436 10678 4488 10684
rect 4540 10606 4568 11591
rect 4632 11354 4660 12815
rect 4802 12200 4858 12209
rect 4802 12135 4858 12144
rect 4710 11384 4766 11393
rect 4620 11348 4672 11354
rect 4816 11354 4844 12135
rect 8116 11960 8168 11966
rect 8116 11902 8168 11908
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 5354 11520 5410 11529
rect 5354 11455 5410 11464
rect 4710 11319 4766 11328
rect 4804 11348 4856 11354
rect 4620 11290 4672 11296
rect 4724 11150 4752 11319
rect 4804 11290 4856 11296
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5092 10849 5120 10950
rect 5078 10840 5134 10849
rect 5184 10810 5212 10950
rect 5078 10775 5134 10784
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 4804 10736 4856 10742
rect 4856 10696 4936 10724
rect 4804 10678 4856 10684
rect 4528 10600 4580 10606
rect 4066 10568 4122 10577
rect 4620 10600 4672 10606
rect 4528 10542 4580 10548
rect 4618 10568 4620 10577
rect 4672 10568 4674 10577
rect 4066 10503 4122 10512
rect 4618 10503 4674 10512
rect 4080 10470 4108 10503
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4172 10305 4200 10406
rect 4158 10296 4214 10305
rect 3516 10260 3568 10266
rect 4158 10231 4214 10240
rect 4802 10296 4858 10305
rect 4802 10231 4858 10240
rect 3516 10202 3568 10208
rect 3974 10160 4030 10169
rect 3974 10095 3976 10104
rect 4028 10095 4030 10104
rect 3976 10066 4028 10072
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3200 8928 3280 8956
rect 3344 9064 3464 9092
rect 3148 8910 3200 8916
rect 3056 7948 3108 7954
rect 2792 7908 2912 7936
rect 2884 7868 2912 7908
rect 3056 7890 3108 7896
rect 2332 7840 2452 7868
rect 2884 7840 3004 7868
rect 2056 7806 2268 7834
rect 2240 7800 2268 7806
rect 2240 7772 2352 7800
rect 2136 7744 2188 7750
rect 1964 7704 2084 7732
rect 1858 7440 1914 7449
rect 1858 7375 1914 7384
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 6497 1900 6666
rect 1964 6633 1992 7346
rect 2056 7313 2084 7704
rect 2324 7732 2352 7772
rect 2188 7704 2268 7732
rect 2324 7704 2360 7732
rect 2136 7686 2188 7692
rect 2134 7440 2190 7449
rect 2134 7375 2190 7384
rect 2042 7304 2098 7313
rect 2042 7239 2098 7248
rect 2148 7206 2176 7375
rect 2240 7313 2268 7704
rect 2226 7304 2282 7313
rect 2226 7239 2282 7248
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 1950 6624 2006 6633
rect 1950 6559 2006 6568
rect 1858 6488 1914 6497
rect 1858 6423 1914 6432
rect 2056 6361 2084 7142
rect 2134 7032 2190 7041
rect 2134 6967 2190 6976
rect 2148 6458 2176 6967
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2042 6352 2098 6361
rect 2042 6287 2098 6296
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1492 5636 1544 5642
rect 1492 5578 1544 5584
rect 2332 2378 2360 7704
rect 2424 7206 2452 7840
rect 2504 7744 2556 7750
rect 2780 7744 2832 7750
rect 2556 7704 2728 7732
rect 2504 7686 2556 7692
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2516 7313 2544 7414
rect 2700 7313 2728 7704
rect 2780 7686 2832 7692
rect 2502 7304 2558 7313
rect 2502 7239 2558 7248
rect 2686 7304 2742 7313
rect 2686 7239 2742 7248
rect 2412 7200 2464 7206
rect 2792 7188 2820 7686
rect 2412 7142 2464 7148
rect 2508 7160 2820 7188
rect 2508 6984 2536 7160
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 2508 6956 2544 6984
rect 2516 5137 2544 6956
rect 2976 6905 3004 7840
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 2962 6896 3018 6905
rect 2962 6831 3018 6840
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2608 5273 2636 6598
rect 2872 6384 2924 6390
rect 3068 6361 3096 7686
rect 3160 7290 3188 8910
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 7954 3280 8774
rect 3344 8566 3372 9064
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3436 8129 3464 8910
rect 3514 8528 3570 8537
rect 3514 8463 3570 8472
rect 3422 8120 3478 8129
rect 3422 8055 3478 8064
rect 3422 7984 3478 7993
rect 3240 7948 3292 7954
rect 3422 7919 3478 7928
rect 3240 7890 3292 7896
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7410 3280 7686
rect 3436 7585 3464 7919
rect 3528 7818 3556 8463
rect 3516 7812 3568 7818
rect 3516 7754 3568 7760
rect 3422 7576 3478 7585
rect 3422 7511 3478 7520
rect 3436 7410 3464 7511
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3160 7262 3464 7290
rect 3330 7168 3386 7177
rect 3330 7103 3386 7112
rect 3146 7032 3202 7041
rect 3146 6967 3202 6976
rect 3240 6996 3292 7002
rect 3160 6497 3188 6967
rect 3240 6938 3292 6944
rect 3252 6798 3280 6938
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3146 6488 3202 6497
rect 3146 6423 3202 6432
rect 2872 6326 2924 6332
rect 3054 6352 3110 6361
rect 2594 5264 2650 5273
rect 2594 5199 2650 5208
rect 2502 5128 2558 5137
rect 2502 5063 2558 5072
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2700 4457 2728 4490
rect 2686 4448 2742 4457
rect 2686 4383 2742 4392
rect 2884 3738 2912 6326
rect 3054 6287 3110 6296
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3056 5704 3108 5710
rect 3160 5681 3188 6258
rect 3252 6254 3280 6598
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3344 5817 3372 7103
rect 3330 5808 3386 5817
rect 3330 5743 3386 5752
rect 3056 5646 3108 5652
rect 3146 5672 3202 5681
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 3068 3398 3096 5646
rect 3146 5607 3202 5616
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4214 3280 4558
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3344 3482 3372 4694
rect 3436 4672 3464 7262
rect 3528 6633 3556 7346
rect 3514 6624 3570 6633
rect 3514 6559 3570 6568
rect 3528 5930 3556 6559
rect 3620 6118 3648 9862
rect 3608 6112 3660 6118
rect 3712 6089 3740 9998
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 3804 9353 3832 9930
rect 4116 9820 4424 9840
rect 4116 9818 4122 9820
rect 4178 9818 4202 9820
rect 4258 9818 4282 9820
rect 4338 9818 4362 9820
rect 4418 9818 4424 9820
rect 4178 9766 4180 9818
rect 4360 9766 4362 9818
rect 4116 9764 4122 9766
rect 4178 9764 4202 9766
rect 4258 9764 4282 9766
rect 4338 9764 4362 9766
rect 4418 9764 4424 9766
rect 4116 9744 4424 9764
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3790 9344 3846 9353
rect 3790 9279 3846 9288
rect 3896 8906 3924 9522
rect 4448 9178 4476 9590
rect 4540 9382 4568 9998
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4526 9208 4582 9217
rect 4436 9172 4488 9178
rect 4526 9143 4582 9152
rect 4436 9114 4488 9120
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3896 8634 3924 8842
rect 4116 8732 4424 8752
rect 4116 8730 4122 8732
rect 4178 8730 4202 8732
rect 4258 8730 4282 8732
rect 4338 8730 4362 8732
rect 4418 8730 4424 8732
rect 4178 8678 4180 8730
rect 4360 8678 4362 8730
rect 4116 8676 4122 8678
rect 4178 8676 4202 8678
rect 4258 8676 4282 8678
rect 4338 8676 4362 8678
rect 4418 8676 4424 8678
rect 4116 8656 4424 8676
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3804 8514 3832 8570
rect 3804 8498 4384 8514
rect 3804 8492 4396 8498
rect 3804 8486 4344 8492
rect 4344 8434 4396 8440
rect 4540 8430 4568 9143
rect 4724 8634 4752 9454
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4526 8256 4582 8265
rect 4526 8191 4582 8200
rect 3804 8044 4292 8072
rect 3804 7721 3832 8044
rect 4068 7880 4120 7886
rect 3988 7840 4068 7868
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3790 7712 3846 7721
rect 3790 7647 3846 7656
rect 3896 7449 3924 7754
rect 3882 7440 3938 7449
rect 3988 7410 4016 7840
rect 4068 7822 4120 7828
rect 4264 7818 4292 8044
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4540 7750 4568 8191
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4116 7644 4424 7664
rect 4116 7642 4122 7644
rect 4178 7642 4202 7644
rect 4258 7642 4282 7644
rect 4338 7642 4362 7644
rect 4418 7642 4424 7644
rect 4178 7590 4180 7642
rect 4360 7590 4362 7642
rect 4116 7588 4122 7590
rect 4178 7588 4202 7590
rect 4258 7588 4282 7590
rect 4338 7588 4362 7590
rect 4418 7588 4424 7590
rect 4116 7568 4424 7588
rect 3882 7375 3938 7384
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3790 7304 3846 7313
rect 3790 7239 3792 7248
rect 3844 7239 3846 7248
rect 3792 7210 3844 7216
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3896 7002 3924 7142
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3988 6882 4016 7346
rect 4540 7324 4568 7686
rect 4632 7478 4660 7686
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4540 7296 4660 7324
rect 3896 6866 4016 6882
rect 3884 6860 4016 6866
rect 3936 6854 4016 6860
rect 3884 6802 3936 6808
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3804 6662 3832 6734
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3608 6054 3660 6060
rect 3698 6080 3754 6089
rect 3698 6015 3754 6024
rect 3528 5902 3648 5930
rect 3804 5914 3832 6598
rect 3896 6118 3924 6598
rect 3988 6390 4016 6854
rect 4526 6896 4582 6905
rect 4526 6831 4582 6840
rect 4116 6556 4424 6576
rect 4116 6554 4122 6556
rect 4178 6554 4202 6556
rect 4258 6554 4282 6556
rect 4338 6554 4362 6556
rect 4418 6554 4424 6556
rect 4178 6502 4180 6554
rect 4360 6502 4362 6554
rect 4116 6500 4122 6502
rect 4178 6500 4202 6502
rect 4258 6500 4282 6502
rect 4338 6500 4362 6502
rect 4418 6500 4424 6502
rect 4116 6480 4424 6500
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 4158 6352 4214 6361
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3436 4644 3556 4672
rect 3424 4548 3476 4554
rect 3424 4490 3476 4496
rect 3436 3602 3464 4490
rect 3528 4146 3556 4644
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3620 3942 3648 5902
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3988 5778 4016 6326
rect 4158 6287 4160 6296
rect 4212 6287 4214 6296
rect 4434 6352 4490 6361
rect 4540 6322 4568 6831
rect 4434 6287 4490 6296
rect 4528 6316 4580 6322
rect 4160 6258 4212 6264
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4172 6089 4200 6122
rect 4158 6080 4214 6089
rect 4158 6015 4214 6024
rect 4448 5953 4476 6287
rect 4528 6258 4580 6264
rect 4434 5944 4490 5953
rect 4434 5879 4490 5888
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3344 3454 3464 3482
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3344 2650 3372 2926
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 2320 2372 2372 2378
rect 2320 2314 2372 2320
rect 3436 513 3464 3454
rect 3528 2446 3556 3878
rect 3712 3602 3740 5510
rect 3988 5234 4016 5714
rect 4116 5468 4424 5488
rect 4116 5466 4122 5468
rect 4178 5466 4202 5468
rect 4258 5466 4282 5468
rect 4338 5466 4362 5468
rect 4418 5466 4424 5468
rect 4178 5414 4180 5466
rect 4360 5414 4362 5466
rect 4116 5412 4122 5414
rect 4178 5412 4202 5414
rect 4258 5412 4282 5414
rect 4338 5412 4362 5414
rect 4418 5412 4424 5414
rect 4116 5392 4424 5412
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3988 4554 4016 5170
rect 4632 4729 4660 7296
rect 4618 4720 4674 4729
rect 4618 4655 4674 4664
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 4116 4380 4424 4400
rect 4116 4378 4122 4380
rect 4178 4378 4202 4380
rect 4258 4378 4282 4380
rect 4338 4378 4362 4380
rect 4418 4378 4424 4380
rect 4178 4326 4180 4378
rect 4360 4326 4362 4378
rect 4116 4324 4122 4326
rect 4178 4324 4202 4326
rect 4258 4324 4282 4326
rect 4338 4324 4362 4326
rect 4418 4324 4424 4326
rect 4116 4304 4424 4324
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3896 3720 3924 4150
rect 4724 4049 4752 7958
rect 4816 7041 4844 10231
rect 4908 8906 4936 10696
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9178 5028 9998
rect 5078 9480 5134 9489
rect 5078 9415 5134 9424
rect 5092 9382 5120 9415
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5184 9042 5212 10746
rect 5276 9674 5304 11018
rect 5368 9738 5396 11455
rect 5666 11452 5974 11472
rect 5666 11450 5672 11452
rect 5728 11450 5752 11452
rect 5808 11450 5832 11452
rect 5888 11450 5912 11452
rect 5968 11450 5974 11452
rect 5728 11398 5730 11450
rect 5910 11398 5912 11450
rect 5666 11396 5672 11398
rect 5728 11396 5752 11398
rect 5808 11396 5832 11398
rect 5888 11396 5912 11398
rect 5968 11396 5974 11398
rect 5666 11376 5974 11396
rect 5632 11212 5684 11218
rect 5684 11172 5948 11200
rect 5632 11154 5684 11160
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10690 5580 11086
rect 5460 10662 5580 10690
rect 5920 10674 5948 11172
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5908 10668 5960 10674
rect 5460 10010 5488 10662
rect 5908 10610 5960 10616
rect 5666 10364 5974 10384
rect 5666 10362 5672 10364
rect 5728 10362 5752 10364
rect 5808 10362 5832 10364
rect 5888 10362 5912 10364
rect 5968 10362 5974 10364
rect 5728 10310 5730 10362
rect 5910 10310 5912 10362
rect 5666 10308 5672 10310
rect 5728 10308 5752 10310
rect 5808 10308 5832 10310
rect 5888 10308 5912 10310
rect 5968 10308 5974 10310
rect 5666 10288 5974 10308
rect 5908 10192 5960 10198
rect 5906 10160 5908 10169
rect 5960 10160 5962 10169
rect 5906 10095 5962 10104
rect 5460 9994 5580 10010
rect 5460 9988 5592 9994
rect 5460 9982 5540 9988
rect 5540 9930 5592 9936
rect 5368 9722 5580 9738
rect 5368 9716 5592 9722
rect 5368 9710 5540 9716
rect 5276 9646 5394 9674
rect 5540 9658 5592 9664
rect 5366 9602 5394 9646
rect 5446 9616 5502 9625
rect 5366 9574 5396 9602
rect 5368 9500 5396 9574
rect 5446 9551 5502 9560
rect 5540 9580 5592 9586
rect 5276 9472 5396 9500
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 4908 8809 4936 8842
rect 4894 8800 4950 8809
rect 4894 8735 4950 8744
rect 4908 8294 4936 8735
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4802 7032 4858 7041
rect 4802 6967 4858 6976
rect 4816 4146 4844 6967
rect 4908 6254 4936 8230
rect 4986 8120 5042 8129
rect 4986 8055 5042 8064
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4908 5914 4936 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5000 5642 5028 8055
rect 5184 7970 5212 8842
rect 5092 7954 5212 7970
rect 5080 7948 5212 7954
rect 5132 7942 5212 7948
rect 5080 7890 5132 7896
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5092 7721 5120 7754
rect 5078 7712 5134 7721
rect 5078 7647 5134 7656
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5092 5114 5120 6666
rect 5184 6066 5212 7942
rect 5276 6662 5304 9472
rect 5460 9178 5488 9551
rect 5540 9522 5592 9528
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 7800 5396 8230
rect 5460 7954 5488 8910
rect 5552 8362 5580 9522
rect 6012 9518 6040 11086
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6104 10577 6132 10950
rect 6090 10568 6146 10577
rect 6090 10503 6146 10512
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5666 9276 5974 9296
rect 5666 9274 5672 9276
rect 5728 9274 5752 9276
rect 5808 9274 5832 9276
rect 5888 9274 5912 9276
rect 5968 9274 5974 9276
rect 5728 9222 5730 9274
rect 5910 9222 5912 9274
rect 5666 9220 5672 9222
rect 5728 9220 5752 9222
rect 5808 9220 5832 9222
rect 5888 9220 5912 9222
rect 5968 9220 5974 9222
rect 5666 9200 5974 9220
rect 6012 8906 6040 9318
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5816 8832 5868 8838
rect 6012 8809 6040 8842
rect 5816 8774 5868 8780
rect 5998 8800 6054 8809
rect 5828 8634 5856 8774
rect 5998 8735 6054 8744
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5666 8188 5974 8208
rect 5666 8186 5672 8188
rect 5728 8186 5752 8188
rect 5808 8186 5832 8188
rect 5888 8186 5912 8188
rect 5968 8186 5974 8188
rect 5728 8134 5730 8186
rect 5910 8134 5912 8186
rect 5666 8132 5672 8134
rect 5728 8132 5752 8134
rect 5808 8132 5832 8134
rect 5888 8132 5912 8134
rect 5968 8132 5974 8134
rect 5666 8112 5974 8132
rect 6012 8090 6040 8230
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5448 7812 5500 7818
rect 5368 7772 5448 7800
rect 5368 7478 5396 7772
rect 5448 7754 5500 7760
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5460 6905 5488 7210
rect 5446 6896 5502 6905
rect 5446 6831 5502 6840
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 6458 5304 6598
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5184 6038 5488 6066
rect 5460 5846 5488 6038
rect 5448 5840 5500 5846
rect 5170 5808 5226 5817
rect 5354 5808 5410 5817
rect 5170 5743 5226 5752
rect 5264 5772 5316 5778
rect 5184 5710 5212 5743
rect 5448 5782 5500 5788
rect 5354 5743 5410 5752
rect 5264 5714 5316 5720
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5276 5302 5304 5714
rect 5264 5296 5316 5302
rect 5000 5086 5120 5114
rect 5184 5256 5264 5284
rect 5000 5030 5028 5086
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5184 4758 5212 5256
rect 5264 5238 5316 5244
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5276 4826 5304 5034
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4710 4040 4766 4049
rect 4710 3975 4766 3984
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 3896 3692 4016 3720
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3712 3058 3740 3538
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3896 2106 3924 2246
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 3422 504 3478 513
rect 3422 439 3478 448
rect 3988 241 4016 3692
rect 4116 3292 4424 3312
rect 4116 3290 4122 3292
rect 4178 3290 4202 3292
rect 4258 3290 4282 3292
rect 4338 3290 4362 3292
rect 4418 3290 4424 3292
rect 4178 3238 4180 3290
rect 4360 3238 4362 3290
rect 4116 3236 4122 3238
rect 4178 3236 4202 3238
rect 4258 3236 4282 3238
rect 4338 3236 4362 3238
rect 4418 3236 4424 3238
rect 4116 3216 4424 3236
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4172 2650 4200 3062
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4068 2440 4120 2446
rect 4344 2440 4396 2446
rect 4120 2400 4344 2428
rect 4068 2382 4120 2388
rect 4344 2382 4396 2388
rect 4116 2204 4424 2224
rect 4116 2202 4122 2204
rect 4178 2202 4202 2204
rect 4258 2202 4282 2204
rect 4338 2202 4362 2204
rect 4418 2202 4424 2204
rect 4178 2150 4180 2202
rect 4360 2150 4362 2202
rect 4116 2148 4122 2150
rect 4178 2148 4202 2150
rect 4258 2148 4282 2150
rect 4338 2148 4362 2150
rect 4418 2148 4424 2150
rect 4116 2128 4424 2148
rect 4724 1465 4752 3878
rect 5092 3738 5120 4626
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4896 3596 4948 3602
rect 5184 3584 5212 4694
rect 5368 4570 5396 5743
rect 5552 5250 5580 7278
rect 5666 7100 5974 7120
rect 5666 7098 5672 7100
rect 5728 7098 5752 7100
rect 5808 7098 5832 7100
rect 5888 7098 5912 7100
rect 5968 7098 5974 7100
rect 5728 7046 5730 7098
rect 5910 7046 5912 7098
rect 5666 7044 5672 7046
rect 5728 7044 5752 7046
rect 5808 7044 5832 7046
rect 5888 7044 5912 7046
rect 5968 7044 5974 7046
rect 5666 7024 5974 7044
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5666 6012 5974 6032
rect 5666 6010 5672 6012
rect 5728 6010 5752 6012
rect 5808 6010 5832 6012
rect 5888 6010 5912 6012
rect 5968 6010 5974 6012
rect 5728 5958 5730 6010
rect 5910 5958 5912 6010
rect 5666 5956 5672 5958
rect 5728 5956 5752 5958
rect 5808 5956 5832 5958
rect 5888 5956 5912 5958
rect 5968 5956 5974 5958
rect 5666 5936 5974 5956
rect 5906 5808 5962 5817
rect 5906 5743 5962 5752
rect 5724 5704 5776 5710
rect 5722 5672 5724 5681
rect 5776 5672 5778 5681
rect 5722 5607 5778 5616
rect 5552 5222 5672 5250
rect 5644 5166 5672 5222
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5552 4826 5580 5102
rect 5920 5098 5948 5743
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5666 4924 5974 4944
rect 5666 4922 5672 4924
rect 5728 4922 5752 4924
rect 5808 4922 5832 4924
rect 5888 4922 5912 4924
rect 5968 4922 5974 4924
rect 5728 4870 5730 4922
rect 5910 4870 5912 4922
rect 5666 4868 5672 4870
rect 5728 4868 5752 4870
rect 5808 4868 5832 4870
rect 5888 4868 5912 4870
rect 5968 4868 5974 4870
rect 5666 4848 5974 4868
rect 6012 4826 6040 6258
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5552 4690 5580 4762
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5632 4616 5684 4622
rect 5368 4564 5632 4570
rect 5368 4558 5684 4564
rect 5368 4542 5672 4558
rect 6104 4282 6132 8978
rect 6196 6866 6224 11562
rect 6274 11384 6330 11393
rect 6274 11319 6330 11328
rect 6288 11082 6316 11319
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6380 10169 6408 10950
rect 6366 10160 6422 10169
rect 6366 10095 6422 10104
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 8498 6316 9522
rect 6472 8650 6500 11086
rect 6550 10840 6606 10849
rect 6550 10775 6606 10784
rect 6564 10062 6592 10775
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6656 9926 6684 11834
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6748 9450 6776 11630
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11370 6868 11494
rect 6840 11342 6960 11370
rect 7024 11354 7328 11370
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6840 10198 6868 11154
rect 6932 10742 6960 11342
rect 7012 11348 7340 11354
rect 7064 11342 7288 11348
rect 7012 11290 7064 11296
rect 7288 11290 7340 11296
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6828 10192 6880 10198
rect 7012 10192 7064 10198
rect 6828 10134 6880 10140
rect 6932 10152 7012 10180
rect 6932 9586 6960 10152
rect 7012 10134 7064 10140
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6932 9382 6960 9522
rect 7024 9518 7052 9930
rect 7116 9674 7144 11154
rect 7208 11082 7236 11154
rect 7288 11144 7340 11150
rect 7392 11132 7420 11698
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7484 11150 7512 11630
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7340 11104 7420 11132
rect 7472 11144 7524 11150
rect 7288 11086 7340 11092
rect 7472 11086 7524 11092
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7576 11014 7604 11494
rect 7668 11150 7696 11562
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 11008 7616 11014
rect 7760 10985 7788 11290
rect 7564 10950 7616 10956
rect 7746 10976 7802 10985
rect 7216 10908 7524 10928
rect 7746 10911 7802 10920
rect 7216 10906 7222 10908
rect 7278 10906 7302 10908
rect 7358 10906 7382 10908
rect 7438 10906 7462 10908
rect 7518 10906 7524 10908
rect 7278 10854 7280 10906
rect 7460 10854 7462 10906
rect 7216 10852 7222 10854
rect 7278 10852 7302 10854
rect 7358 10852 7382 10854
rect 7438 10852 7462 10854
rect 7518 10852 7524 10854
rect 7216 10832 7524 10852
rect 8128 10674 8156 11902
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 8766 11452 9074 11472
rect 8766 11450 8772 11452
rect 8828 11450 8852 11452
rect 8908 11450 8932 11452
rect 8988 11450 9012 11452
rect 9068 11450 9074 11452
rect 8828 11398 8830 11450
rect 9010 11398 9012 11450
rect 8766 11396 8772 11398
rect 8828 11396 8852 11398
rect 8908 11396 8932 11398
rect 8988 11396 9012 11398
rect 9068 11396 9074 11398
rect 8390 11384 8446 11393
rect 8766 11376 9074 11396
rect 8390 11319 8446 11328
rect 8404 11150 8432 11319
rect 8574 11248 8630 11257
rect 8574 11183 8630 11192
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8206 10704 8262 10713
rect 8116 10668 8168 10674
rect 8206 10639 8262 10648
rect 8116 10610 8168 10616
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 7208 9994 7236 10134
rect 7472 10056 7524 10062
rect 7524 10016 7604 10044
rect 7472 9998 7524 10004
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7216 9820 7524 9840
rect 7216 9818 7222 9820
rect 7278 9818 7302 9820
rect 7358 9818 7382 9820
rect 7438 9818 7462 9820
rect 7518 9818 7524 9820
rect 7278 9766 7280 9818
rect 7460 9766 7462 9818
rect 7216 9764 7222 9766
rect 7278 9764 7302 9766
rect 7358 9764 7382 9766
rect 7438 9764 7462 9766
rect 7518 9764 7524 9766
rect 7216 9744 7524 9764
rect 7576 9722 7604 10016
rect 8036 9994 8064 10134
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 7564 9716 7616 9722
rect 7116 9646 7236 9674
rect 7564 9658 7616 9664
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6736 9104 6788 9110
rect 6380 8622 6500 8650
rect 6656 9064 6736 9092
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6288 5914 6316 6326
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6380 5794 6408 8622
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6472 8090 6500 8434
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6472 7410 6500 8026
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6472 6361 6500 6802
rect 6458 6352 6514 6361
rect 6458 6287 6514 6296
rect 6564 6254 6592 8298
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6288 5766 6408 5794
rect 6196 5370 6224 5714
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 4948 3556 5212 3584
rect 4896 3538 4948 3544
rect 5184 2854 5212 3556
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5184 2582 5212 2790
rect 5172 2576 5224 2582
rect 5172 2518 5224 2524
rect 5184 2378 5212 2518
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 5368 2038 5396 2994
rect 5460 2446 5488 4014
rect 5666 3836 5974 3856
rect 5666 3834 5672 3836
rect 5728 3834 5752 3836
rect 5808 3834 5832 3836
rect 5888 3834 5912 3836
rect 5968 3834 5974 3836
rect 5728 3782 5730 3834
rect 5910 3782 5912 3834
rect 5666 3780 5672 3782
rect 5728 3780 5752 3782
rect 5808 3780 5832 3782
rect 5888 3780 5912 3782
rect 5968 3780 5974 3782
rect 5666 3760 5974 3780
rect 5540 3528 5592 3534
rect 6000 3528 6052 3534
rect 5540 3470 5592 3476
rect 5630 3496 5686 3505
rect 5552 2650 5580 3470
rect 6000 3470 6052 3476
rect 5630 3431 5632 3440
rect 5684 3431 5686 3440
rect 5632 3402 5684 3408
rect 5666 2748 5974 2768
rect 5666 2746 5672 2748
rect 5728 2746 5752 2748
rect 5808 2746 5832 2748
rect 5888 2746 5912 2748
rect 5968 2746 5974 2748
rect 5728 2694 5730 2746
rect 5910 2694 5912 2746
rect 5666 2692 5672 2694
rect 5728 2692 5752 2694
rect 5808 2692 5832 2694
rect 5888 2692 5912 2694
rect 5968 2692 5974 2694
rect 5666 2672 5974 2692
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 6012 2106 6040 3470
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6104 2514 6132 3130
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 6196 2446 6224 2994
rect 6288 2990 6316 5766
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6380 4622 6408 5578
rect 6472 4758 6500 5646
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6564 4486 6592 6190
rect 6656 5817 6684 9064
rect 6736 9046 6788 9052
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 6254 6776 8366
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6840 7954 6868 8298
rect 6932 7954 6960 9318
rect 7116 8566 7144 9318
rect 7208 8820 7236 9646
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 9110 7512 9454
rect 7472 9104 7524 9110
rect 7576 9081 7604 9658
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7472 9046 7524 9052
rect 7562 9072 7618 9081
rect 7562 9007 7618 9016
rect 7208 8792 7604 8820
rect 7216 8732 7524 8752
rect 7216 8730 7222 8732
rect 7278 8730 7302 8732
rect 7358 8730 7382 8732
rect 7438 8730 7462 8732
rect 7518 8730 7524 8732
rect 7278 8678 7280 8730
rect 7460 8678 7462 8730
rect 7216 8676 7222 8678
rect 7278 8676 7302 8678
rect 7358 8676 7382 8678
rect 7438 8676 7462 8678
rect 7518 8676 7524 8678
rect 7216 8656 7524 8676
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7208 8090 7236 8366
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6932 7818 6960 7890
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 6918 7712 6974 7721
rect 6918 7647 6974 7656
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6642 5808 6698 5817
rect 6642 5743 6698 5752
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6380 3602 6408 4014
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6276 2984 6328 2990
rect 6274 2952 6276 2961
rect 6328 2952 6330 2961
rect 6274 2887 6330 2896
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6472 2310 6500 4082
rect 6564 2650 6592 4150
rect 6656 3738 6684 5646
rect 6748 5166 6776 6190
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6748 4622 6776 5102
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6748 4078 6776 4558
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3738 6776 3878
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6656 3058 6684 3538
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3058 6776 3334
rect 6840 3194 6868 7278
rect 6932 5681 6960 7647
rect 7116 7002 7144 7754
rect 7216 7644 7524 7664
rect 7216 7642 7222 7644
rect 7278 7642 7302 7644
rect 7358 7642 7382 7644
rect 7438 7642 7462 7644
rect 7518 7642 7524 7644
rect 7278 7590 7280 7642
rect 7460 7590 7462 7642
rect 7216 7588 7222 7590
rect 7278 7588 7302 7590
rect 7358 7588 7382 7590
rect 7438 7588 7462 7590
rect 7518 7588 7524 7590
rect 7216 7568 7524 7588
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7216 6556 7524 6576
rect 7216 6554 7222 6556
rect 7278 6554 7302 6556
rect 7358 6554 7382 6556
rect 7438 6554 7462 6556
rect 7518 6554 7524 6556
rect 7278 6502 7280 6554
rect 7460 6502 7462 6554
rect 7216 6500 7222 6502
rect 7278 6500 7302 6502
rect 7358 6500 7382 6502
rect 7438 6500 7462 6502
rect 7518 6500 7524 6502
rect 7216 6480 7524 6500
rect 7012 6248 7064 6254
rect 7010 6216 7012 6225
rect 7064 6216 7066 6225
rect 7010 6151 7066 6160
rect 7576 5760 7604 8792
rect 7668 6390 7696 9318
rect 7944 8022 7972 9522
rect 8036 9518 8064 9930
rect 8128 9722 8156 9930
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8220 9586 8248 10639
rect 8312 10266 8340 11086
rect 8588 11014 8616 11183
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8496 9625 8524 10950
rect 9232 10810 9260 11086
rect 9402 10840 9458 10849
rect 9220 10804 9272 10810
rect 9402 10775 9458 10784
rect 9220 10746 9272 10752
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8482 9616 8538 9625
rect 8208 9580 8260 9586
rect 8482 9551 8538 9560
rect 8208 9522 8260 9528
rect 8024 9512 8076 9518
rect 8576 9512 8628 9518
rect 8024 9454 8076 9460
rect 8482 9480 8538 9489
rect 8576 9454 8628 9460
rect 8482 9415 8538 9424
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 8036 7546 8064 8910
rect 8312 8786 8340 8910
rect 8128 8758 8340 8786
rect 8128 8430 8156 8758
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8128 7562 8156 7958
rect 8220 7886 8248 8570
rect 8312 8022 8340 8758
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8024 7540 8076 7546
rect 8128 7534 8248 7562
rect 8024 7482 8076 7488
rect 7840 7404 7892 7410
rect 7892 7364 8156 7392
rect 7840 7346 7892 7352
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7760 6118 7788 6938
rect 8024 6792 8076 6798
rect 8022 6760 8024 6769
rect 8076 6760 8078 6769
rect 8022 6695 8078 6704
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7748 6112 7800 6118
rect 7932 6112 7984 6118
rect 7800 6072 7880 6100
rect 7748 6054 7800 6060
rect 7576 5732 7788 5760
rect 6918 5672 6974 5681
rect 6918 5607 6974 5616
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7216 5468 7524 5488
rect 7216 5466 7222 5468
rect 7278 5466 7302 5468
rect 7358 5466 7382 5468
rect 7438 5466 7462 5468
rect 7518 5466 7524 5468
rect 7278 5414 7280 5466
rect 7460 5414 7462 5466
rect 7216 5412 7222 5414
rect 7278 5412 7302 5414
rect 7358 5412 7382 5414
rect 7438 5412 7462 5414
rect 7518 5412 7524 5414
rect 7216 5392 7524 5412
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 7116 4282 7144 5238
rect 7216 4380 7524 4400
rect 7216 4378 7222 4380
rect 7278 4378 7302 4380
rect 7358 4378 7382 4380
rect 7438 4378 7462 4380
rect 7518 4378 7524 4380
rect 7278 4326 7280 4378
rect 7460 4326 7462 4378
rect 7216 4324 7222 4326
rect 7278 4324 7302 4326
rect 7358 4324 7382 4326
rect 7438 4324 7462 4326
rect 7518 4324 7524 4326
rect 7216 4304 7524 4324
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7208 3670 7236 4082
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7216 3292 7524 3312
rect 7216 3290 7222 3292
rect 7278 3290 7302 3292
rect 7358 3290 7382 3292
rect 7438 3290 7462 3292
rect 7518 3290 7524 3292
rect 7278 3238 7280 3290
rect 7460 3238 7462 3290
rect 7216 3236 7222 3238
rect 7278 3236 7302 3238
rect 7358 3236 7382 3238
rect 7438 3236 7462 3238
rect 7518 3236 7524 3238
rect 7216 3216 7524 3236
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6656 2446 6684 2994
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6748 2378 6776 2994
rect 6826 2952 6882 2961
rect 6882 2922 7052 2938
rect 6882 2916 7064 2922
rect 6882 2910 7012 2916
rect 6826 2887 6882 2896
rect 7012 2858 7064 2864
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 2514 6868 2790
rect 7576 2650 7604 5578
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7668 4282 7696 5170
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7668 3670 7696 4082
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7760 3534 7788 5732
rect 7852 5370 7880 6072
rect 7932 6054 7984 6060
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4146 7880 4966
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7944 3641 7972 6054
rect 7930 3632 7986 3641
rect 7930 3567 7986 3576
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 7852 2310 7880 3402
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 3126 7972 3334
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 8036 2514 8064 6598
rect 8128 3398 8156 7364
rect 8220 7274 8248 7534
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8496 7018 8524 9415
rect 8588 9042 8616 9454
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8588 7857 8616 8842
rect 8574 7848 8630 7857
rect 8574 7783 8630 7792
rect 8496 6990 8616 7018
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8208 6316 8260 6322
rect 8312 6304 8340 6734
rect 8404 6458 8432 6734
rect 8588 6474 8616 6990
rect 8680 6662 8708 10542
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 8766 10364 9074 10384
rect 8766 10362 8772 10364
rect 8828 10362 8852 10364
rect 8908 10362 8932 10364
rect 8988 10362 9012 10364
rect 9068 10362 9074 10364
rect 8828 10310 8830 10362
rect 9010 10310 9012 10362
rect 8766 10308 8772 10310
rect 8828 10308 8852 10310
rect 8908 10308 8932 10310
rect 8988 10308 9012 10310
rect 9068 10308 9074 10310
rect 8766 10288 9074 10308
rect 9324 10130 9352 10474
rect 9416 10441 9444 10775
rect 9402 10432 9458 10441
rect 9402 10367 9458 10376
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9218 10024 9274 10033
rect 9218 9959 9220 9968
rect 9272 9959 9274 9968
rect 9220 9930 9272 9936
rect 8766 9276 9074 9296
rect 8766 9274 8772 9276
rect 8828 9274 8852 9276
rect 8908 9274 8932 9276
rect 8988 9274 9012 9276
rect 9068 9274 9074 9276
rect 8828 9222 8830 9274
rect 9010 9222 9012 9274
rect 8766 9220 8772 9222
rect 8828 9220 8852 9222
rect 8908 9220 8932 9222
rect 8988 9220 9012 9222
rect 9068 9220 9074 9222
rect 8766 9200 9074 9220
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8766 8188 9074 8208
rect 8766 8186 8772 8188
rect 8828 8186 8852 8188
rect 8908 8186 8932 8188
rect 8988 8186 9012 8188
rect 9068 8186 9074 8188
rect 8828 8134 8830 8186
rect 9010 8134 9012 8186
rect 8766 8132 8772 8134
rect 8828 8132 8852 8134
rect 8908 8132 8932 8134
rect 8988 8132 9012 8134
rect 9068 8132 9074 8134
rect 8766 8112 9074 8132
rect 8760 7880 8812 7886
rect 8758 7848 8760 7857
rect 8812 7848 8814 7857
rect 8758 7783 8814 7792
rect 9140 7410 9168 8774
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9232 8090 9260 8502
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9324 7546 9352 8434
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8766 7100 9074 7120
rect 8766 7098 8772 7100
rect 8828 7098 8852 7100
rect 8908 7098 8932 7100
rect 8988 7098 9012 7100
rect 9068 7098 9074 7100
rect 8828 7046 8830 7098
rect 9010 7046 9012 7098
rect 8766 7044 8772 7046
rect 8828 7044 8852 7046
rect 8908 7044 8932 7046
rect 8988 7044 9012 7046
rect 9068 7044 9074 7046
rect 8766 7024 9074 7044
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8864 6662 8892 6734
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8392 6452 8444 6458
rect 8588 6446 9076 6474
rect 9140 6458 9168 6734
rect 8392 6394 8444 6400
rect 8668 6316 8720 6322
rect 8312 6276 8432 6304
rect 8208 6258 8260 6264
rect 8220 5846 8248 6258
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8312 5234 8340 6122
rect 8404 5302 8432 6276
rect 8668 6258 8720 6264
rect 8680 5914 8708 6258
rect 9048 6202 9076 6446
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9220 6248 9272 6254
rect 9048 6174 9168 6202
rect 9220 6190 9272 6196
rect 8766 6012 9074 6032
rect 8766 6010 8772 6012
rect 8828 6010 8852 6012
rect 8908 6010 8932 6012
rect 8988 6010 9012 6012
rect 9068 6010 9074 6012
rect 8828 5958 8830 6010
rect 9010 5958 9012 6010
rect 8766 5956 8772 5958
rect 8828 5956 8852 5958
rect 8908 5956 8932 5958
rect 8988 5956 9012 5958
rect 9068 5956 9074 5958
rect 8766 5936 9074 5956
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8206 5128 8262 5137
rect 8206 5063 8262 5072
rect 8220 4146 8248 5063
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8312 3942 8340 4490
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8404 3738 8432 4082
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8206 3632 8262 3641
rect 8206 3567 8262 3576
rect 8220 3534 8248 3567
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8298 3496 8354 3505
rect 8298 3431 8354 3440
rect 8312 3398 8340 3431
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8404 3058 8432 3674
rect 8496 3194 8524 5646
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 8956 5370 8984 5578
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8588 5137 8616 5170
rect 8574 5128 8630 5137
rect 8574 5063 8630 5072
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8588 4214 8616 4558
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8680 3942 8708 5306
rect 8766 4924 9074 4944
rect 8766 4922 8772 4924
rect 8828 4922 8852 4924
rect 8908 4922 8932 4924
rect 8988 4922 9012 4924
rect 9068 4922 9074 4924
rect 8828 4870 8830 4922
rect 9010 4870 9012 4922
rect 8766 4868 8772 4870
rect 8828 4868 8852 4870
rect 8908 4868 8932 4870
rect 8988 4868 9012 4870
rect 9068 4868 9074 4870
rect 8766 4848 9074 4868
rect 9140 4078 9168 6174
rect 9232 4826 9260 6190
rect 9324 6118 9352 6802
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9324 4146 9352 6054
rect 9416 5914 9444 8910
rect 9508 8634 9536 11698
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9508 8106 9536 8570
rect 9784 8265 9812 11630
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13266 10432 13322 10441
rect 13266 10367 13322 10376
rect 9770 8256 9826 8265
rect 9770 8191 9826 8200
rect 9508 8078 9628 8106
rect 9600 7206 9628 8078
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9416 4146 9444 4966
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8680 3738 8708 3878
rect 8766 3836 9074 3856
rect 8766 3834 8772 3836
rect 8828 3834 8852 3836
rect 8908 3834 8932 3836
rect 8988 3834 9012 3836
rect 9068 3834 9074 3836
rect 8828 3782 8830 3834
rect 9010 3782 9012 3834
rect 8766 3780 8772 3782
rect 8828 3780 8852 3782
rect 8908 3780 8932 3782
rect 8988 3780 9012 3782
rect 9068 3780 9074 3782
rect 8766 3760 9074 3780
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8680 3466 8708 3674
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8128 2650 8156 2790
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8496 2446 8524 2858
rect 8588 2650 8616 3062
rect 9508 3058 9536 4966
rect 9600 4593 9628 6870
rect 9586 4584 9642 4593
rect 9586 4519 9642 4528
rect 13280 3369 13308 10367
rect 13372 7721 13400 11494
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 8129 13492 11154
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13450 8120 13506 8129
rect 13450 8055 13506 8064
rect 13452 8016 13504 8022
rect 13450 7984 13452 7993
rect 13504 7984 13506 7993
rect 13450 7919 13506 7928
rect 13358 7712 13414 7721
rect 13358 7647 13414 7656
rect 13450 7440 13506 7449
rect 13450 7375 13506 7384
rect 13464 3777 13492 7375
rect 13556 7041 13584 8774
rect 13648 7313 13676 9046
rect 13740 8945 13768 11290
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13832 9353 13860 11222
rect 16684 11014 16712 13495
rect 22098 11248 22154 11257
rect 22098 11183 22154 11192
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13726 8936 13782 8945
rect 13726 8871 13782 8880
rect 13726 8528 13782 8537
rect 13726 8463 13728 8472
rect 13780 8463 13782 8472
rect 13728 8434 13780 8440
rect 13820 8424 13872 8430
rect 13818 8392 13820 8401
rect 13872 8392 13874 8401
rect 13818 8327 13874 8336
rect 13634 7304 13690 7313
rect 13634 7239 13690 7248
rect 13818 7168 13874 7177
rect 13818 7103 13820 7112
rect 13872 7103 13874 7112
rect 19800 7132 19852 7138
rect 13820 7074 13872 7080
rect 19800 7074 19852 7080
rect 13542 7032 13598 7041
rect 13542 6967 13598 6976
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13542 6624 13598 6633
rect 13542 6559 13598 6568
rect 13556 4010 13584 6559
rect 13648 5001 13676 6938
rect 13726 6352 13782 6361
rect 13726 6287 13782 6296
rect 13740 5098 13768 6287
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13832 6089 13860 6122
rect 13818 6080 13874 6089
rect 13818 6015 13874 6024
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13634 4992 13690 5001
rect 13634 4927 13690 4936
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13450 3768 13506 3777
rect 13450 3703 13506 3712
rect 13266 3360 13322 3369
rect 13266 3295 13322 3304
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 8766 2748 9074 2768
rect 8766 2746 8772 2748
rect 8828 2746 8852 2748
rect 8908 2746 8932 2748
rect 8988 2746 9012 2748
rect 9068 2746 9074 2748
rect 8828 2694 8830 2746
rect 9010 2694 9012 2746
rect 8766 2692 8772 2694
rect 8828 2692 8852 2694
rect 8908 2692 8932 2694
rect 8988 2692 9012 2694
rect 9068 2692 9074 2694
rect 8766 2672 9074 2692
rect 9140 2650 9168 2926
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 6288 2106 6316 2246
rect 7216 2204 7524 2224
rect 7216 2202 7222 2204
rect 7278 2202 7302 2204
rect 7358 2202 7382 2204
rect 7438 2202 7462 2204
rect 7518 2202 7524 2204
rect 7278 2150 7280 2202
rect 7460 2150 7462 2202
rect 7216 2148 7222 2150
rect 7278 2148 7302 2150
rect 7358 2148 7382 2150
rect 7438 2148 7462 2150
rect 7518 2148 7524 2150
rect 7216 2128 7524 2148
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 8864 2038 8892 2246
rect 9048 2106 9076 2382
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 5356 2032 5408 2038
rect 5356 1974 5408 1980
rect 8852 2032 8904 2038
rect 8852 1974 8904 1980
rect 4710 1456 4766 1465
rect 4710 1391 4766 1400
rect 9324 785 9352 2790
rect 19812 1193 19840 7074
rect 22112 6730 22140 11183
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22204 2825 22232 8366
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22190 2816 22246 2825
rect 22190 2751 22246 2760
rect 22296 2417 22324 7958
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22282 2408 22338 2417
rect 22282 2343 22338 2352
rect 22388 1737 22416 7890
rect 22480 3097 22508 8434
rect 22744 8288 22796 8294
rect 22744 8230 22796 8236
rect 22466 3088 22522 3097
rect 22466 3023 22522 3032
rect 22756 2145 22784 8230
rect 22742 2136 22798 2145
rect 22742 2071 22798 2080
rect 22374 1728 22430 1737
rect 22374 1663 22430 1672
rect 19798 1184 19854 1193
rect 19798 1119 19854 1128
rect 9310 776 9366 785
rect 9310 711 9366 720
rect 3974 232 4030 241
rect 3974 167 4030 176
<< via2 >>
rect 2042 13776 2098 13832
rect 1950 12416 2006 12472
rect 1674 11600 1730 11656
rect 1214 11056 1270 11112
rect 1398 10668 1454 10704
rect 1398 10648 1400 10668
rect 1400 10648 1452 10668
rect 1452 10648 1454 10668
rect 16670 13504 16726 13560
rect 3974 13096 4030 13152
rect 2226 11736 2282 11792
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2686 11192 2742 11248
rect 3054 10784 3110 10840
rect 2778 10648 2834 10704
rect 2318 9696 2374 9752
rect 2134 9424 2190 9480
rect 1214 7656 1270 7712
rect 1122 6704 1178 6760
rect 1030 5888 1086 5944
rect 1674 7792 1730 7848
rect 1674 7520 1730 7576
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2502 10104 2558 10160
rect 2870 10104 2926 10160
rect 3422 11464 3478 11520
rect 3514 11328 3570 11384
rect 3238 9968 3294 10024
rect 2870 9560 2926 9616
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2318 8880 2374 8936
rect 2226 8336 2282 8392
rect 2594 8916 2596 8936
rect 2596 8916 2648 8936
rect 2648 8916 2650 8936
rect 2594 8880 2650 8916
rect 2778 8472 2834 8528
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2410 7964 2412 7984
rect 2412 7964 2464 7984
rect 2464 7964 2466 7984
rect 2410 7928 2466 7964
rect 3422 10784 3478 10840
rect 3330 9152 3386 9208
rect 4618 12824 4674 12880
rect 4526 11600 4582 11656
rect 4122 10906 4178 10908
rect 4202 10906 4258 10908
rect 4282 10906 4338 10908
rect 4362 10906 4418 10908
rect 4122 10854 4168 10906
rect 4168 10854 4178 10906
rect 4202 10854 4232 10906
rect 4232 10854 4244 10906
rect 4244 10854 4258 10906
rect 4282 10854 4296 10906
rect 4296 10854 4308 10906
rect 4308 10854 4338 10906
rect 4362 10854 4372 10906
rect 4372 10854 4418 10906
rect 4122 10852 4178 10854
rect 4202 10852 4258 10854
rect 4282 10852 4338 10854
rect 4362 10852 4418 10854
rect 4802 12144 4858 12200
rect 4710 11328 4766 11384
rect 5354 11464 5410 11520
rect 5078 10784 5134 10840
rect 4066 10512 4122 10568
rect 4618 10548 4620 10568
rect 4620 10548 4672 10568
rect 4672 10548 4674 10568
rect 4618 10512 4674 10548
rect 4158 10240 4214 10296
rect 4802 10240 4858 10296
rect 3974 10124 4030 10160
rect 3974 10104 3976 10124
rect 3976 10104 4028 10124
rect 4028 10104 4030 10124
rect 1858 7384 1914 7440
rect 2134 7384 2190 7440
rect 2042 7248 2098 7304
rect 2226 7248 2282 7304
rect 1950 6568 2006 6624
rect 1858 6432 1914 6488
rect 2134 6976 2190 7032
rect 2042 6296 2098 6352
rect 2502 7248 2558 7304
rect 2686 7248 2742 7304
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2962 6840 3018 6896
rect 3514 8472 3570 8528
rect 3422 8064 3478 8120
rect 3422 7928 3478 7984
rect 3422 7520 3478 7576
rect 3330 7112 3386 7168
rect 3146 6976 3202 7032
rect 3146 6432 3202 6488
rect 2594 5208 2650 5264
rect 2502 5072 2558 5128
rect 2686 4392 2742 4448
rect 3054 6296 3110 6352
rect 3330 5752 3386 5808
rect 3146 5616 3202 5672
rect 3514 6568 3570 6624
rect 4122 9818 4178 9820
rect 4202 9818 4258 9820
rect 4282 9818 4338 9820
rect 4362 9818 4418 9820
rect 4122 9766 4168 9818
rect 4168 9766 4178 9818
rect 4202 9766 4232 9818
rect 4232 9766 4244 9818
rect 4244 9766 4258 9818
rect 4282 9766 4296 9818
rect 4296 9766 4308 9818
rect 4308 9766 4338 9818
rect 4362 9766 4372 9818
rect 4372 9766 4418 9818
rect 4122 9764 4178 9766
rect 4202 9764 4258 9766
rect 4282 9764 4338 9766
rect 4362 9764 4418 9766
rect 3790 9288 3846 9344
rect 4526 9152 4582 9208
rect 4122 8730 4178 8732
rect 4202 8730 4258 8732
rect 4282 8730 4338 8732
rect 4362 8730 4418 8732
rect 4122 8678 4168 8730
rect 4168 8678 4178 8730
rect 4202 8678 4232 8730
rect 4232 8678 4244 8730
rect 4244 8678 4258 8730
rect 4282 8678 4296 8730
rect 4296 8678 4308 8730
rect 4308 8678 4338 8730
rect 4362 8678 4372 8730
rect 4372 8678 4418 8730
rect 4122 8676 4178 8678
rect 4202 8676 4258 8678
rect 4282 8676 4338 8678
rect 4362 8676 4418 8678
rect 4526 8200 4582 8256
rect 3790 7656 3846 7712
rect 3882 7384 3938 7440
rect 4122 7642 4178 7644
rect 4202 7642 4258 7644
rect 4282 7642 4338 7644
rect 4362 7642 4418 7644
rect 4122 7590 4168 7642
rect 4168 7590 4178 7642
rect 4202 7590 4232 7642
rect 4232 7590 4244 7642
rect 4244 7590 4258 7642
rect 4282 7590 4296 7642
rect 4296 7590 4308 7642
rect 4308 7590 4338 7642
rect 4362 7590 4372 7642
rect 4372 7590 4418 7642
rect 4122 7588 4178 7590
rect 4202 7588 4258 7590
rect 4282 7588 4338 7590
rect 4362 7588 4418 7590
rect 3790 7268 3846 7304
rect 3790 7248 3792 7268
rect 3792 7248 3844 7268
rect 3844 7248 3846 7268
rect 3698 6024 3754 6080
rect 4526 6840 4582 6896
rect 4122 6554 4178 6556
rect 4202 6554 4258 6556
rect 4282 6554 4338 6556
rect 4362 6554 4418 6556
rect 4122 6502 4168 6554
rect 4168 6502 4178 6554
rect 4202 6502 4232 6554
rect 4232 6502 4244 6554
rect 4244 6502 4258 6554
rect 4282 6502 4296 6554
rect 4296 6502 4308 6554
rect 4308 6502 4338 6554
rect 4362 6502 4372 6554
rect 4372 6502 4418 6554
rect 4122 6500 4178 6502
rect 4202 6500 4258 6502
rect 4282 6500 4338 6502
rect 4362 6500 4418 6502
rect 4158 6316 4214 6352
rect 4158 6296 4160 6316
rect 4160 6296 4212 6316
rect 4212 6296 4214 6316
rect 4434 6296 4490 6352
rect 4158 6024 4214 6080
rect 4434 5888 4490 5944
rect 4122 5466 4178 5468
rect 4202 5466 4258 5468
rect 4282 5466 4338 5468
rect 4362 5466 4418 5468
rect 4122 5414 4168 5466
rect 4168 5414 4178 5466
rect 4202 5414 4232 5466
rect 4232 5414 4244 5466
rect 4244 5414 4258 5466
rect 4282 5414 4296 5466
rect 4296 5414 4308 5466
rect 4308 5414 4338 5466
rect 4362 5414 4372 5466
rect 4372 5414 4418 5466
rect 4122 5412 4178 5414
rect 4202 5412 4258 5414
rect 4282 5412 4338 5414
rect 4362 5412 4418 5414
rect 4618 4664 4674 4720
rect 4122 4378 4178 4380
rect 4202 4378 4258 4380
rect 4282 4378 4338 4380
rect 4362 4378 4418 4380
rect 4122 4326 4168 4378
rect 4168 4326 4178 4378
rect 4202 4326 4232 4378
rect 4232 4326 4244 4378
rect 4244 4326 4258 4378
rect 4282 4326 4296 4378
rect 4296 4326 4308 4378
rect 4308 4326 4338 4378
rect 4362 4326 4372 4378
rect 4372 4326 4418 4378
rect 4122 4324 4178 4326
rect 4202 4324 4258 4326
rect 4282 4324 4338 4326
rect 4362 4324 4418 4326
rect 5078 9424 5134 9480
rect 5672 11450 5728 11452
rect 5752 11450 5808 11452
rect 5832 11450 5888 11452
rect 5912 11450 5968 11452
rect 5672 11398 5718 11450
rect 5718 11398 5728 11450
rect 5752 11398 5782 11450
rect 5782 11398 5794 11450
rect 5794 11398 5808 11450
rect 5832 11398 5846 11450
rect 5846 11398 5858 11450
rect 5858 11398 5888 11450
rect 5912 11398 5922 11450
rect 5922 11398 5968 11450
rect 5672 11396 5728 11398
rect 5752 11396 5808 11398
rect 5832 11396 5888 11398
rect 5912 11396 5968 11398
rect 5672 10362 5728 10364
rect 5752 10362 5808 10364
rect 5832 10362 5888 10364
rect 5912 10362 5968 10364
rect 5672 10310 5718 10362
rect 5718 10310 5728 10362
rect 5752 10310 5782 10362
rect 5782 10310 5794 10362
rect 5794 10310 5808 10362
rect 5832 10310 5846 10362
rect 5846 10310 5858 10362
rect 5858 10310 5888 10362
rect 5912 10310 5922 10362
rect 5922 10310 5968 10362
rect 5672 10308 5728 10310
rect 5752 10308 5808 10310
rect 5832 10308 5888 10310
rect 5912 10308 5968 10310
rect 5906 10140 5908 10160
rect 5908 10140 5960 10160
rect 5960 10140 5962 10160
rect 5906 10104 5962 10140
rect 5446 9560 5502 9616
rect 4894 8744 4950 8800
rect 4802 6976 4858 7032
rect 4986 8064 5042 8120
rect 5078 7656 5134 7712
rect 6090 10512 6146 10568
rect 5672 9274 5728 9276
rect 5752 9274 5808 9276
rect 5832 9274 5888 9276
rect 5912 9274 5968 9276
rect 5672 9222 5718 9274
rect 5718 9222 5728 9274
rect 5752 9222 5782 9274
rect 5782 9222 5794 9274
rect 5794 9222 5808 9274
rect 5832 9222 5846 9274
rect 5846 9222 5858 9274
rect 5858 9222 5888 9274
rect 5912 9222 5922 9274
rect 5922 9222 5968 9274
rect 5672 9220 5728 9222
rect 5752 9220 5808 9222
rect 5832 9220 5888 9222
rect 5912 9220 5968 9222
rect 5998 8744 6054 8800
rect 5672 8186 5728 8188
rect 5752 8186 5808 8188
rect 5832 8186 5888 8188
rect 5912 8186 5968 8188
rect 5672 8134 5718 8186
rect 5718 8134 5728 8186
rect 5752 8134 5782 8186
rect 5782 8134 5794 8186
rect 5794 8134 5808 8186
rect 5832 8134 5846 8186
rect 5846 8134 5858 8186
rect 5858 8134 5888 8186
rect 5912 8134 5922 8186
rect 5922 8134 5968 8186
rect 5672 8132 5728 8134
rect 5752 8132 5808 8134
rect 5832 8132 5888 8134
rect 5912 8132 5968 8134
rect 5446 6840 5502 6896
rect 5170 5752 5226 5808
rect 5354 5752 5410 5808
rect 4710 3984 4766 4040
rect 3422 448 3478 504
rect 4122 3290 4178 3292
rect 4202 3290 4258 3292
rect 4282 3290 4338 3292
rect 4362 3290 4418 3292
rect 4122 3238 4168 3290
rect 4168 3238 4178 3290
rect 4202 3238 4232 3290
rect 4232 3238 4244 3290
rect 4244 3238 4258 3290
rect 4282 3238 4296 3290
rect 4296 3238 4308 3290
rect 4308 3238 4338 3290
rect 4362 3238 4372 3290
rect 4372 3238 4418 3290
rect 4122 3236 4178 3238
rect 4202 3236 4258 3238
rect 4282 3236 4338 3238
rect 4362 3236 4418 3238
rect 4122 2202 4178 2204
rect 4202 2202 4258 2204
rect 4282 2202 4338 2204
rect 4362 2202 4418 2204
rect 4122 2150 4168 2202
rect 4168 2150 4178 2202
rect 4202 2150 4232 2202
rect 4232 2150 4244 2202
rect 4244 2150 4258 2202
rect 4282 2150 4296 2202
rect 4296 2150 4308 2202
rect 4308 2150 4338 2202
rect 4362 2150 4372 2202
rect 4372 2150 4418 2202
rect 4122 2148 4178 2150
rect 4202 2148 4258 2150
rect 4282 2148 4338 2150
rect 4362 2148 4418 2150
rect 5672 7098 5728 7100
rect 5752 7098 5808 7100
rect 5832 7098 5888 7100
rect 5912 7098 5968 7100
rect 5672 7046 5718 7098
rect 5718 7046 5728 7098
rect 5752 7046 5782 7098
rect 5782 7046 5794 7098
rect 5794 7046 5808 7098
rect 5832 7046 5846 7098
rect 5846 7046 5858 7098
rect 5858 7046 5888 7098
rect 5912 7046 5922 7098
rect 5922 7046 5968 7098
rect 5672 7044 5728 7046
rect 5752 7044 5808 7046
rect 5832 7044 5888 7046
rect 5912 7044 5968 7046
rect 5672 6010 5728 6012
rect 5752 6010 5808 6012
rect 5832 6010 5888 6012
rect 5912 6010 5968 6012
rect 5672 5958 5718 6010
rect 5718 5958 5728 6010
rect 5752 5958 5782 6010
rect 5782 5958 5794 6010
rect 5794 5958 5808 6010
rect 5832 5958 5846 6010
rect 5846 5958 5858 6010
rect 5858 5958 5888 6010
rect 5912 5958 5922 6010
rect 5922 5958 5968 6010
rect 5672 5956 5728 5958
rect 5752 5956 5808 5958
rect 5832 5956 5888 5958
rect 5912 5956 5968 5958
rect 5906 5752 5962 5808
rect 5722 5652 5724 5672
rect 5724 5652 5776 5672
rect 5776 5652 5778 5672
rect 5722 5616 5778 5652
rect 5672 4922 5728 4924
rect 5752 4922 5808 4924
rect 5832 4922 5888 4924
rect 5912 4922 5968 4924
rect 5672 4870 5718 4922
rect 5718 4870 5728 4922
rect 5752 4870 5782 4922
rect 5782 4870 5794 4922
rect 5794 4870 5808 4922
rect 5832 4870 5846 4922
rect 5846 4870 5858 4922
rect 5858 4870 5888 4922
rect 5912 4870 5922 4922
rect 5922 4870 5968 4922
rect 5672 4868 5728 4870
rect 5752 4868 5808 4870
rect 5832 4868 5888 4870
rect 5912 4868 5968 4870
rect 6274 11328 6330 11384
rect 6366 10104 6422 10160
rect 6550 10784 6606 10840
rect 7746 10920 7802 10976
rect 7222 10906 7278 10908
rect 7302 10906 7358 10908
rect 7382 10906 7438 10908
rect 7462 10906 7518 10908
rect 7222 10854 7268 10906
rect 7268 10854 7278 10906
rect 7302 10854 7332 10906
rect 7332 10854 7344 10906
rect 7344 10854 7358 10906
rect 7382 10854 7396 10906
rect 7396 10854 7408 10906
rect 7408 10854 7438 10906
rect 7462 10854 7472 10906
rect 7472 10854 7518 10906
rect 7222 10852 7278 10854
rect 7302 10852 7358 10854
rect 7382 10852 7438 10854
rect 7462 10852 7518 10854
rect 8772 11450 8828 11452
rect 8852 11450 8908 11452
rect 8932 11450 8988 11452
rect 9012 11450 9068 11452
rect 8772 11398 8818 11450
rect 8818 11398 8828 11450
rect 8852 11398 8882 11450
rect 8882 11398 8894 11450
rect 8894 11398 8908 11450
rect 8932 11398 8946 11450
rect 8946 11398 8958 11450
rect 8958 11398 8988 11450
rect 9012 11398 9022 11450
rect 9022 11398 9068 11450
rect 8772 11396 8828 11398
rect 8852 11396 8908 11398
rect 8932 11396 8988 11398
rect 9012 11396 9068 11398
rect 8390 11328 8446 11384
rect 8574 11192 8630 11248
rect 8206 10648 8262 10704
rect 7222 9818 7278 9820
rect 7302 9818 7358 9820
rect 7382 9818 7438 9820
rect 7462 9818 7518 9820
rect 7222 9766 7268 9818
rect 7268 9766 7278 9818
rect 7302 9766 7332 9818
rect 7332 9766 7344 9818
rect 7344 9766 7358 9818
rect 7382 9766 7396 9818
rect 7396 9766 7408 9818
rect 7408 9766 7438 9818
rect 7462 9766 7472 9818
rect 7472 9766 7518 9818
rect 7222 9764 7278 9766
rect 7302 9764 7358 9766
rect 7382 9764 7438 9766
rect 7462 9764 7518 9766
rect 6458 6296 6514 6352
rect 5672 3834 5728 3836
rect 5752 3834 5808 3836
rect 5832 3834 5888 3836
rect 5912 3834 5968 3836
rect 5672 3782 5718 3834
rect 5718 3782 5728 3834
rect 5752 3782 5782 3834
rect 5782 3782 5794 3834
rect 5794 3782 5808 3834
rect 5832 3782 5846 3834
rect 5846 3782 5858 3834
rect 5858 3782 5888 3834
rect 5912 3782 5922 3834
rect 5922 3782 5968 3834
rect 5672 3780 5728 3782
rect 5752 3780 5808 3782
rect 5832 3780 5888 3782
rect 5912 3780 5968 3782
rect 5630 3460 5686 3496
rect 5630 3440 5632 3460
rect 5632 3440 5684 3460
rect 5684 3440 5686 3460
rect 5672 2746 5728 2748
rect 5752 2746 5808 2748
rect 5832 2746 5888 2748
rect 5912 2746 5968 2748
rect 5672 2694 5718 2746
rect 5718 2694 5728 2746
rect 5752 2694 5782 2746
rect 5782 2694 5794 2746
rect 5794 2694 5808 2746
rect 5832 2694 5846 2746
rect 5846 2694 5858 2746
rect 5858 2694 5888 2746
rect 5912 2694 5922 2746
rect 5922 2694 5968 2746
rect 5672 2692 5728 2694
rect 5752 2692 5808 2694
rect 5832 2692 5888 2694
rect 5912 2692 5968 2694
rect 7562 9016 7618 9072
rect 7222 8730 7278 8732
rect 7302 8730 7358 8732
rect 7382 8730 7438 8732
rect 7462 8730 7518 8732
rect 7222 8678 7268 8730
rect 7268 8678 7278 8730
rect 7302 8678 7332 8730
rect 7332 8678 7344 8730
rect 7344 8678 7358 8730
rect 7382 8678 7396 8730
rect 7396 8678 7408 8730
rect 7408 8678 7438 8730
rect 7462 8678 7472 8730
rect 7472 8678 7518 8730
rect 7222 8676 7278 8678
rect 7302 8676 7358 8678
rect 7382 8676 7438 8678
rect 7462 8676 7518 8678
rect 6918 7656 6974 7712
rect 6642 5752 6698 5808
rect 6274 2932 6276 2952
rect 6276 2932 6328 2952
rect 6328 2932 6330 2952
rect 6274 2896 6330 2932
rect 7222 7642 7278 7644
rect 7302 7642 7358 7644
rect 7382 7642 7438 7644
rect 7462 7642 7518 7644
rect 7222 7590 7268 7642
rect 7268 7590 7278 7642
rect 7302 7590 7332 7642
rect 7332 7590 7344 7642
rect 7344 7590 7358 7642
rect 7382 7590 7396 7642
rect 7396 7590 7408 7642
rect 7408 7590 7438 7642
rect 7462 7590 7472 7642
rect 7472 7590 7518 7642
rect 7222 7588 7278 7590
rect 7302 7588 7358 7590
rect 7382 7588 7438 7590
rect 7462 7588 7518 7590
rect 7222 6554 7278 6556
rect 7302 6554 7358 6556
rect 7382 6554 7438 6556
rect 7462 6554 7518 6556
rect 7222 6502 7268 6554
rect 7268 6502 7278 6554
rect 7302 6502 7332 6554
rect 7332 6502 7344 6554
rect 7344 6502 7358 6554
rect 7382 6502 7396 6554
rect 7396 6502 7408 6554
rect 7408 6502 7438 6554
rect 7462 6502 7472 6554
rect 7472 6502 7518 6554
rect 7222 6500 7278 6502
rect 7302 6500 7358 6502
rect 7382 6500 7438 6502
rect 7462 6500 7518 6502
rect 7010 6196 7012 6216
rect 7012 6196 7064 6216
rect 7064 6196 7066 6216
rect 7010 6160 7066 6196
rect 9402 10784 9458 10840
rect 8482 9560 8538 9616
rect 8482 9424 8538 9480
rect 8022 6740 8024 6760
rect 8024 6740 8076 6760
rect 8076 6740 8078 6760
rect 8022 6704 8078 6740
rect 6918 5616 6974 5672
rect 7222 5466 7278 5468
rect 7302 5466 7358 5468
rect 7382 5466 7438 5468
rect 7462 5466 7518 5468
rect 7222 5414 7268 5466
rect 7268 5414 7278 5466
rect 7302 5414 7332 5466
rect 7332 5414 7344 5466
rect 7344 5414 7358 5466
rect 7382 5414 7396 5466
rect 7396 5414 7408 5466
rect 7408 5414 7438 5466
rect 7462 5414 7472 5466
rect 7472 5414 7518 5466
rect 7222 5412 7278 5414
rect 7302 5412 7358 5414
rect 7382 5412 7438 5414
rect 7462 5412 7518 5414
rect 7222 4378 7278 4380
rect 7302 4378 7358 4380
rect 7382 4378 7438 4380
rect 7462 4378 7518 4380
rect 7222 4326 7268 4378
rect 7268 4326 7278 4378
rect 7302 4326 7332 4378
rect 7332 4326 7344 4378
rect 7344 4326 7358 4378
rect 7382 4326 7396 4378
rect 7396 4326 7408 4378
rect 7408 4326 7438 4378
rect 7462 4326 7472 4378
rect 7472 4326 7518 4378
rect 7222 4324 7278 4326
rect 7302 4324 7358 4326
rect 7382 4324 7438 4326
rect 7462 4324 7518 4326
rect 7222 3290 7278 3292
rect 7302 3290 7358 3292
rect 7382 3290 7438 3292
rect 7462 3290 7518 3292
rect 7222 3238 7268 3290
rect 7268 3238 7278 3290
rect 7302 3238 7332 3290
rect 7332 3238 7344 3290
rect 7344 3238 7358 3290
rect 7382 3238 7396 3290
rect 7396 3238 7408 3290
rect 7408 3238 7438 3290
rect 7462 3238 7472 3290
rect 7472 3238 7518 3290
rect 7222 3236 7278 3238
rect 7302 3236 7358 3238
rect 7382 3236 7438 3238
rect 7462 3236 7518 3238
rect 6826 2896 6882 2952
rect 7930 3576 7986 3632
rect 8574 7792 8630 7848
rect 8772 10362 8828 10364
rect 8852 10362 8908 10364
rect 8932 10362 8988 10364
rect 9012 10362 9068 10364
rect 8772 10310 8818 10362
rect 8818 10310 8828 10362
rect 8852 10310 8882 10362
rect 8882 10310 8894 10362
rect 8894 10310 8908 10362
rect 8932 10310 8946 10362
rect 8946 10310 8958 10362
rect 8958 10310 8988 10362
rect 9012 10310 9022 10362
rect 9022 10310 9068 10362
rect 8772 10308 8828 10310
rect 8852 10308 8908 10310
rect 8932 10308 8988 10310
rect 9012 10308 9068 10310
rect 9402 10376 9458 10432
rect 9218 9988 9274 10024
rect 9218 9968 9220 9988
rect 9220 9968 9272 9988
rect 9272 9968 9274 9988
rect 8772 9274 8828 9276
rect 8852 9274 8908 9276
rect 8932 9274 8988 9276
rect 9012 9274 9068 9276
rect 8772 9222 8818 9274
rect 8818 9222 8828 9274
rect 8852 9222 8882 9274
rect 8882 9222 8894 9274
rect 8894 9222 8908 9274
rect 8932 9222 8946 9274
rect 8946 9222 8958 9274
rect 8958 9222 8988 9274
rect 9012 9222 9022 9274
rect 9022 9222 9068 9274
rect 8772 9220 8828 9222
rect 8852 9220 8908 9222
rect 8932 9220 8988 9222
rect 9012 9220 9068 9222
rect 8772 8186 8828 8188
rect 8852 8186 8908 8188
rect 8932 8186 8988 8188
rect 9012 8186 9068 8188
rect 8772 8134 8818 8186
rect 8818 8134 8828 8186
rect 8852 8134 8882 8186
rect 8882 8134 8894 8186
rect 8894 8134 8908 8186
rect 8932 8134 8946 8186
rect 8946 8134 8958 8186
rect 8958 8134 8988 8186
rect 9012 8134 9022 8186
rect 9022 8134 9068 8186
rect 8772 8132 8828 8134
rect 8852 8132 8908 8134
rect 8932 8132 8988 8134
rect 9012 8132 9068 8134
rect 8758 7828 8760 7848
rect 8760 7828 8812 7848
rect 8812 7828 8814 7848
rect 8758 7792 8814 7828
rect 8772 7098 8828 7100
rect 8852 7098 8908 7100
rect 8932 7098 8988 7100
rect 9012 7098 9068 7100
rect 8772 7046 8818 7098
rect 8818 7046 8828 7098
rect 8852 7046 8882 7098
rect 8882 7046 8894 7098
rect 8894 7046 8908 7098
rect 8932 7046 8946 7098
rect 8946 7046 8958 7098
rect 8958 7046 8988 7098
rect 9012 7046 9022 7098
rect 9022 7046 9068 7098
rect 8772 7044 8828 7046
rect 8852 7044 8908 7046
rect 8932 7044 8988 7046
rect 9012 7044 9068 7046
rect 8772 6010 8828 6012
rect 8852 6010 8908 6012
rect 8932 6010 8988 6012
rect 9012 6010 9068 6012
rect 8772 5958 8818 6010
rect 8818 5958 8828 6010
rect 8852 5958 8882 6010
rect 8882 5958 8894 6010
rect 8894 5958 8908 6010
rect 8932 5958 8946 6010
rect 8946 5958 8958 6010
rect 8958 5958 8988 6010
rect 9012 5958 9022 6010
rect 9022 5958 9068 6010
rect 8772 5956 8828 5958
rect 8852 5956 8908 5958
rect 8932 5956 8988 5958
rect 9012 5956 9068 5958
rect 8206 5072 8262 5128
rect 8206 3576 8262 3632
rect 8298 3440 8354 3496
rect 8574 5072 8630 5128
rect 8772 4922 8828 4924
rect 8852 4922 8908 4924
rect 8932 4922 8988 4924
rect 9012 4922 9068 4924
rect 8772 4870 8818 4922
rect 8818 4870 8828 4922
rect 8852 4870 8882 4922
rect 8882 4870 8894 4922
rect 8894 4870 8908 4922
rect 8932 4870 8946 4922
rect 8946 4870 8958 4922
rect 8958 4870 8988 4922
rect 9012 4870 9022 4922
rect 9022 4870 9068 4922
rect 8772 4868 8828 4870
rect 8852 4868 8908 4870
rect 8932 4868 8988 4870
rect 9012 4868 9068 4870
rect 13266 10376 13322 10432
rect 9770 8200 9826 8256
rect 8772 3834 8828 3836
rect 8852 3834 8908 3836
rect 8932 3834 8988 3836
rect 9012 3834 9068 3836
rect 8772 3782 8818 3834
rect 8818 3782 8828 3834
rect 8852 3782 8882 3834
rect 8882 3782 8894 3834
rect 8894 3782 8908 3834
rect 8932 3782 8946 3834
rect 8946 3782 8958 3834
rect 8958 3782 8988 3834
rect 9012 3782 9022 3834
rect 9022 3782 9068 3834
rect 8772 3780 8828 3782
rect 8852 3780 8908 3782
rect 8932 3780 8988 3782
rect 9012 3780 9068 3782
rect 9586 4528 9642 4584
rect 13450 8064 13506 8120
rect 13450 7964 13452 7984
rect 13452 7964 13504 7984
rect 13504 7964 13506 7984
rect 13450 7928 13506 7964
rect 13358 7656 13414 7712
rect 13450 7384 13506 7440
rect 22098 11192 22154 11248
rect 13818 9288 13874 9344
rect 13726 8880 13782 8936
rect 13726 8492 13782 8528
rect 13726 8472 13728 8492
rect 13728 8472 13780 8492
rect 13780 8472 13782 8492
rect 13818 8372 13820 8392
rect 13820 8372 13872 8392
rect 13872 8372 13874 8392
rect 13818 8336 13874 8372
rect 13634 7248 13690 7304
rect 13818 7132 13874 7168
rect 13818 7112 13820 7132
rect 13820 7112 13872 7132
rect 13872 7112 13874 7132
rect 13542 6976 13598 7032
rect 13542 6568 13598 6624
rect 13726 6296 13782 6352
rect 13818 6024 13874 6080
rect 13634 4936 13690 4992
rect 13450 3712 13506 3768
rect 13266 3304 13322 3360
rect 8772 2746 8828 2748
rect 8852 2746 8908 2748
rect 8932 2746 8988 2748
rect 9012 2746 9068 2748
rect 8772 2694 8818 2746
rect 8818 2694 8828 2746
rect 8852 2694 8882 2746
rect 8882 2694 8894 2746
rect 8894 2694 8908 2746
rect 8932 2694 8946 2746
rect 8946 2694 8958 2746
rect 8958 2694 8988 2746
rect 9012 2694 9022 2746
rect 9022 2694 9068 2746
rect 8772 2692 8828 2694
rect 8852 2692 8908 2694
rect 8932 2692 8988 2694
rect 9012 2692 9068 2694
rect 7222 2202 7278 2204
rect 7302 2202 7358 2204
rect 7382 2202 7438 2204
rect 7462 2202 7518 2204
rect 7222 2150 7268 2202
rect 7268 2150 7278 2202
rect 7302 2150 7332 2202
rect 7332 2150 7344 2202
rect 7344 2150 7358 2202
rect 7382 2150 7396 2202
rect 7396 2150 7408 2202
rect 7408 2150 7438 2202
rect 7462 2150 7472 2202
rect 7472 2150 7518 2202
rect 7222 2148 7278 2150
rect 7302 2148 7358 2150
rect 7382 2148 7438 2150
rect 7462 2148 7518 2150
rect 4710 1400 4766 1456
rect 22190 2760 22246 2816
rect 22282 2352 22338 2408
rect 22466 3032 22522 3088
rect 22742 2080 22798 2136
rect 22374 1672 22430 1728
rect 19798 1128 19854 1184
rect 9310 720 9366 776
rect 3974 176 4030 232
<< metal3 >>
rect 2037 13834 2103 13837
rect 14000 13834 34000 13864
rect 2037 13832 34000 13834
rect 2037 13776 2042 13832
rect 2098 13776 34000 13832
rect 2037 13774 34000 13776
rect 2037 13771 2103 13774
rect 14000 13744 34000 13774
rect 14000 13560 34000 13592
rect 14000 13504 16670 13560
rect 16726 13504 34000 13560
rect 14000 13472 34000 13504
rect 3969 13154 4035 13157
rect 14000 13154 34000 13184
rect 3969 13152 34000 13154
rect 3969 13096 3974 13152
rect 4030 13096 34000 13152
rect 3969 13094 34000 13096
rect 3969 13091 4035 13094
rect 14000 13064 34000 13094
rect 4613 12882 4679 12885
rect 14000 12882 34000 12912
rect 4613 12880 34000 12882
rect 4613 12824 4618 12880
rect 4674 12824 34000 12880
rect 4613 12822 34000 12824
rect 4613 12819 4679 12822
rect 14000 12792 34000 12822
rect 14000 12610 34000 12640
rect 6870 12550 34000 12610
rect 1945 12474 2011 12477
rect 6870 12474 6930 12550
rect 14000 12520 34000 12550
rect 1945 12472 6930 12474
rect 1945 12416 1950 12472
rect 2006 12416 6930 12472
rect 1945 12414 6930 12416
rect 1945 12411 2011 12414
rect 4797 12202 4863 12205
rect 14000 12202 34000 12232
rect 4797 12200 34000 12202
rect 4797 12144 4802 12200
rect 4858 12144 34000 12200
rect 4797 12142 34000 12144
rect 4797 12139 4863 12142
rect 14000 12112 34000 12142
rect 14000 11930 34000 11960
rect 2730 11870 34000 11930
rect 2221 11794 2287 11797
rect 2730 11794 2790 11870
rect 14000 11840 34000 11870
rect 2221 11792 2790 11794
rect 2221 11736 2226 11792
rect 2282 11736 2790 11792
rect 2221 11734 2790 11736
rect 2221 11731 2287 11734
rect 1669 11658 1735 11661
rect 4521 11658 4587 11661
rect 1669 11656 4587 11658
rect 1669 11600 1674 11656
rect 1730 11600 4526 11656
rect 4582 11600 4587 11656
rect 1669 11598 4587 11600
rect 1669 11595 1735 11598
rect 4521 11595 4587 11598
rect 3417 11522 3483 11525
rect 5349 11522 5415 11525
rect 14000 11522 34000 11552
rect 3417 11520 5415 11522
rect 3417 11464 3422 11520
rect 3478 11464 5354 11520
rect 5410 11464 5415 11520
rect 3417 11462 5415 11464
rect 3417 11459 3483 11462
rect 5349 11459 5415 11462
rect 12390 11462 34000 11522
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 5660 11456 5980 11457
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 11391 5980 11392
rect 8760 11456 9080 11457
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 8760 11391 9080 11392
rect 3509 11386 3575 11389
rect 4705 11386 4771 11389
rect 3509 11384 4771 11386
rect 3509 11328 3514 11384
rect 3570 11328 4710 11384
rect 4766 11328 4771 11384
rect 3509 11326 4771 11328
rect 3509 11323 3575 11326
rect 4705 11323 4771 11326
rect 6269 11386 6335 11389
rect 8385 11386 8451 11389
rect 6269 11384 8451 11386
rect 6269 11328 6274 11384
rect 6330 11328 8390 11384
rect 8446 11328 8451 11384
rect 6269 11326 8451 11328
rect 6269 11323 6335 11326
rect 8385 11323 8451 11326
rect 2681 11250 2747 11253
rect 8569 11250 8635 11253
rect 2681 11248 8635 11250
rect 2681 11192 2686 11248
rect 2742 11192 8574 11248
rect 8630 11192 8635 11248
rect 2681 11190 8635 11192
rect 2681 11187 2747 11190
rect 8569 11187 8635 11190
rect 1209 11114 1275 11117
rect 12390 11114 12450 11462
rect 14000 11432 34000 11462
rect 14000 11248 34000 11280
rect 14000 11192 22098 11248
rect 22154 11192 34000 11248
rect 14000 11160 34000 11192
rect 1209 11112 12450 11114
rect 1209 11056 1214 11112
rect 1270 11056 12450 11112
rect 1209 11054 12450 11056
rect 1209 11051 1275 11054
rect 7741 10978 7807 10981
rect 14000 10978 34000 11008
rect 7741 10976 34000 10978
rect 7741 10920 7746 10976
rect 7802 10920 34000 10976
rect 7741 10918 34000 10920
rect 7741 10915 7807 10918
rect 4110 10912 4430 10913
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 10847 4430 10848
rect 7210 10912 7530 10913
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 14000 10888 34000 10918
rect 7210 10847 7530 10848
rect 3049 10842 3115 10845
rect 3417 10842 3483 10845
rect 3049 10840 3483 10842
rect 3049 10784 3054 10840
rect 3110 10784 3422 10840
rect 3478 10784 3483 10840
rect 3049 10782 3483 10784
rect 3049 10779 3115 10782
rect 3417 10779 3483 10782
rect 5073 10842 5139 10845
rect 6545 10842 6611 10845
rect 9397 10842 9463 10845
rect 5073 10840 6611 10842
rect 5073 10784 5078 10840
rect 5134 10784 6550 10840
rect 6606 10784 6611 10840
rect 5073 10782 6611 10784
rect 5073 10779 5139 10782
rect 6545 10779 6611 10782
rect 7606 10840 9463 10842
rect 7606 10784 9402 10840
rect 9458 10784 9463 10840
rect 7606 10782 9463 10784
rect 1393 10706 1459 10709
rect 2773 10706 2839 10709
rect 7606 10706 7666 10782
rect 9397 10779 9463 10782
rect 1393 10704 2839 10706
rect 1393 10648 1398 10704
rect 1454 10648 2778 10704
rect 2834 10648 2839 10704
rect 1393 10646 2839 10648
rect 1393 10643 1459 10646
rect 2773 10643 2839 10646
rect 3006 10646 7666 10706
rect 8201 10706 8267 10709
rect 8201 10704 13186 10706
rect 8201 10648 8206 10704
rect 8262 10648 13186 10704
rect 8201 10646 13186 10648
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 2497 10162 2563 10165
rect 2865 10162 2931 10165
rect 2497 10160 2931 10162
rect 2497 10104 2502 10160
rect 2558 10104 2870 10160
rect 2926 10104 2931 10160
rect 2497 10102 2931 10104
rect 2497 10099 2563 10102
rect 2865 10099 2931 10102
rect 2313 9754 2379 9757
rect 3006 9754 3066 10646
rect 8201 10643 8267 10646
rect 4061 10570 4127 10573
rect 4613 10570 4679 10573
rect 4061 10568 4679 10570
rect 4061 10512 4066 10568
rect 4122 10512 4618 10568
rect 4674 10512 4679 10568
rect 4061 10510 4679 10512
rect 4061 10507 4127 10510
rect 4613 10507 4679 10510
rect 6085 10570 6151 10573
rect 13126 10570 13186 10646
rect 14000 10570 34000 10600
rect 6085 10568 9322 10570
rect 6085 10512 6090 10568
rect 6146 10512 9322 10568
rect 6085 10510 9322 10512
rect 13126 10510 34000 10570
rect 6085 10507 6151 10510
rect 5660 10368 5980 10369
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 10303 5980 10304
rect 8760 10368 9080 10369
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 10303 9080 10304
rect 4153 10298 4219 10301
rect 4797 10298 4863 10301
rect 4153 10296 4863 10298
rect 4153 10240 4158 10296
rect 4214 10240 4802 10296
rect 4858 10240 4863 10296
rect 4153 10238 4863 10240
rect 9262 10298 9322 10510
rect 14000 10480 34000 10510
rect 9397 10434 9463 10437
rect 13261 10434 13327 10437
rect 9397 10432 13327 10434
rect 9397 10376 9402 10432
rect 9458 10376 13266 10432
rect 13322 10376 13327 10432
rect 9397 10374 13327 10376
rect 9397 10371 9463 10374
rect 13261 10371 13327 10374
rect 14000 10298 34000 10328
rect 9262 10238 34000 10298
rect 4153 10235 4219 10238
rect 4797 10235 4863 10238
rect 14000 10208 34000 10238
rect 3969 10162 4035 10165
rect 5901 10162 5967 10165
rect 3969 10160 5967 10162
rect 3969 10104 3974 10160
rect 4030 10104 5906 10160
rect 5962 10104 5967 10160
rect 3969 10102 5967 10104
rect 3969 10099 4035 10102
rect 5901 10099 5967 10102
rect 6361 10162 6427 10165
rect 6361 10160 12450 10162
rect 6361 10104 6366 10160
rect 6422 10104 12450 10160
rect 6361 10102 12450 10104
rect 6361 10099 6427 10102
rect 3233 10026 3299 10029
rect 9213 10026 9279 10029
rect 3233 10024 9279 10026
rect 3233 9968 3238 10024
rect 3294 9968 9218 10024
rect 9274 9968 9279 10024
rect 3233 9966 9279 9968
rect 3233 9963 3299 9966
rect 9213 9963 9279 9966
rect 12390 9890 12450 10102
rect 14000 9890 34000 9920
rect 12390 9830 34000 9890
rect 4110 9824 4430 9825
rect 4110 9760 4118 9824
rect 4182 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4430 9824
rect 4110 9759 4430 9760
rect 7210 9824 7530 9825
rect 7210 9760 7218 9824
rect 7282 9760 7298 9824
rect 7362 9760 7378 9824
rect 7442 9760 7458 9824
rect 7522 9760 7530 9824
rect 14000 9800 34000 9830
rect 7210 9759 7530 9760
rect 2313 9752 3066 9754
rect 2313 9696 2318 9752
rect 2374 9696 3066 9752
rect 2313 9694 3066 9696
rect 2313 9691 2379 9694
rect 2865 9618 2931 9621
rect 5441 9618 5507 9621
rect 2865 9616 5507 9618
rect 2865 9560 2870 9616
rect 2926 9560 5446 9616
rect 5502 9560 5507 9616
rect 2865 9558 5507 9560
rect 2865 9555 2931 9558
rect 5441 9555 5507 9558
rect 8477 9618 8543 9621
rect 14000 9618 34000 9648
rect 8477 9616 34000 9618
rect 8477 9560 8482 9616
rect 8538 9560 34000 9616
rect 8477 9558 34000 9560
rect 8477 9555 8543 9558
rect 14000 9528 34000 9558
rect 2129 9482 2195 9485
rect 5073 9482 5139 9485
rect 8477 9482 8543 9485
rect 2129 9480 5139 9482
rect 2129 9424 2134 9480
rect 2190 9424 5078 9480
rect 5134 9424 5139 9480
rect 2129 9422 5139 9424
rect 2129 9419 2195 9422
rect 5073 9419 5139 9422
rect 5398 9480 8543 9482
rect 5398 9424 8482 9480
rect 8538 9424 8543 9480
rect 5398 9422 8543 9424
rect 3785 9346 3851 9349
rect 5398 9346 5458 9422
rect 8477 9419 8543 9422
rect 3785 9344 5458 9346
rect 3785 9288 3790 9344
rect 3846 9288 5458 9344
rect 3785 9286 5458 9288
rect 13813 9346 13879 9349
rect 14000 9346 34000 9376
rect 13813 9344 34000 9346
rect 13813 9288 13818 9344
rect 13874 9288 34000 9344
rect 13813 9286 34000 9288
rect 3785 9283 3851 9286
rect 13813 9283 13879 9286
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 5660 9280 5980 9281
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 9215 5980 9216
rect 8760 9280 9080 9281
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 14000 9256 34000 9286
rect 8760 9215 9080 9216
rect 3325 9210 3391 9213
rect 4521 9210 4587 9213
rect 3325 9208 4587 9210
rect 3325 9152 3330 9208
rect 3386 9152 4526 9208
rect 4582 9152 4587 9208
rect 3325 9150 4587 9152
rect 3325 9147 3391 9150
rect 4521 9147 4587 9150
rect 7557 9074 7623 9077
rect 2316 9072 7623 9074
rect 2316 9016 7562 9072
rect 7618 9016 7623 9072
rect 2316 9014 7623 9016
rect 2316 8941 2376 9014
rect 7557 9011 7623 9014
rect 2313 8936 2379 8941
rect 2313 8880 2318 8936
rect 2374 8880 2379 8936
rect 2313 8875 2379 8880
rect 2589 8938 2655 8941
rect 13721 8938 13787 8941
rect 14000 8938 34000 8968
rect 2589 8936 12450 8938
rect 2589 8880 2594 8936
rect 2650 8880 12450 8936
rect 2589 8878 12450 8880
rect 2589 8875 2655 8878
rect 4889 8802 4955 8805
rect 5993 8802 6059 8805
rect 4889 8800 6059 8802
rect 4889 8744 4894 8800
rect 4950 8744 5998 8800
rect 6054 8744 6059 8800
rect 4889 8742 6059 8744
rect 4889 8739 4955 8742
rect 5993 8739 6059 8742
rect 4110 8736 4430 8737
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 8671 4430 8672
rect 7210 8736 7530 8737
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 8671 7530 8672
rect 12390 8666 12450 8878
rect 13721 8936 34000 8938
rect 13721 8880 13726 8936
rect 13782 8880 34000 8936
rect 13721 8878 34000 8880
rect 13721 8875 13787 8878
rect 14000 8848 34000 8878
rect 14000 8666 34000 8696
rect 12390 8606 34000 8666
rect 14000 8576 34000 8606
rect 2773 8530 2839 8533
rect 3509 8530 3575 8533
rect 13721 8530 13787 8533
rect 2773 8528 13787 8530
rect 2773 8472 2778 8528
rect 2834 8472 3514 8528
rect 3570 8472 13726 8528
rect 13782 8472 13787 8528
rect 2773 8470 13787 8472
rect 2773 8467 2839 8470
rect 3509 8467 3575 8470
rect 13721 8467 13787 8470
rect 2221 8394 2287 8397
rect 13813 8394 13879 8397
rect 2221 8392 13879 8394
rect 2221 8336 2226 8392
rect 2282 8336 13818 8392
rect 13874 8336 13879 8392
rect 2221 8334 13879 8336
rect 2221 8331 2287 8334
rect 13813 8331 13879 8334
rect 4521 8258 4587 8261
rect 2960 8256 4587 8258
rect 2960 8200 4526 8256
rect 4582 8200 4587 8256
rect 2960 8198 4587 8200
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 2405 7986 2471 7989
rect 2960 7986 3020 8198
rect 4521 8195 4587 8198
rect 9765 8258 9831 8261
rect 14000 8258 34000 8288
rect 9765 8256 34000 8258
rect 9765 8200 9770 8256
rect 9826 8200 34000 8256
rect 9765 8198 34000 8200
rect 9765 8195 9831 8198
rect 5660 8192 5980 8193
rect 5660 8128 5668 8192
rect 5732 8128 5748 8192
rect 5812 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5980 8192
rect 5660 8127 5980 8128
rect 8760 8192 9080 8193
rect 8760 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 9008 8192
rect 9072 8128 9080 8192
rect 14000 8168 34000 8198
rect 8760 8127 9080 8128
rect 3417 8122 3483 8125
rect 4981 8122 5047 8125
rect 3417 8120 5047 8122
rect 3417 8064 3422 8120
rect 3478 8064 4986 8120
rect 5042 8064 5047 8120
rect 3417 8062 5047 8064
rect 3417 8059 3483 8062
rect 4981 8059 5047 8062
rect 13445 8122 13511 8125
rect 13445 8120 13922 8122
rect 13445 8064 13450 8120
rect 13506 8064 13922 8120
rect 13445 8062 13922 8064
rect 13445 8059 13511 8062
rect 2405 7984 3020 7986
rect 2405 7928 2410 7984
rect 2466 7928 3020 7984
rect 2405 7926 3020 7928
rect 3417 7986 3483 7989
rect 13445 7986 13511 7989
rect 3417 7984 13511 7986
rect 3417 7928 3422 7984
rect 3478 7928 13450 7984
rect 13506 7928 13511 7984
rect 3417 7926 13511 7928
rect 13862 7986 13922 8062
rect 14000 7986 34000 8016
rect 13862 7926 34000 7986
rect 2405 7923 2471 7926
rect 3417 7923 3483 7926
rect 13445 7923 13511 7926
rect 14000 7896 34000 7926
rect 1669 7850 1735 7853
rect 8569 7850 8635 7853
rect 8753 7850 8819 7853
rect 1669 7848 8819 7850
rect 1669 7792 1674 7848
rect 1730 7792 8574 7848
rect 8630 7792 8758 7848
rect 8814 7792 8819 7848
rect 1669 7790 8819 7792
rect 1669 7787 1735 7790
rect 8569 7787 8635 7790
rect 8753 7787 8819 7790
rect 1209 7714 1275 7717
rect 3785 7714 3851 7717
rect 1209 7712 3851 7714
rect 1209 7656 1214 7712
rect 1270 7656 3790 7712
rect 3846 7656 3851 7712
rect 1209 7654 3851 7656
rect 1209 7651 1275 7654
rect 3785 7651 3851 7654
rect 5073 7714 5139 7717
rect 6913 7714 6979 7717
rect 5073 7712 6979 7714
rect 5073 7656 5078 7712
rect 5134 7656 6918 7712
rect 6974 7656 6979 7712
rect 5073 7654 6979 7656
rect 5073 7651 5139 7654
rect 6913 7651 6979 7654
rect 13353 7714 13419 7717
rect 14000 7714 34000 7744
rect 13353 7712 34000 7714
rect 13353 7656 13358 7712
rect 13414 7656 34000 7712
rect 13353 7654 34000 7656
rect 13353 7651 13419 7654
rect 4110 7648 4430 7649
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 7583 4430 7584
rect 7210 7648 7530 7649
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 14000 7624 34000 7654
rect 7210 7583 7530 7584
rect 1669 7578 1735 7581
rect 3417 7578 3483 7581
rect 1669 7576 3483 7578
rect 1669 7520 1674 7576
rect 1730 7520 3422 7576
rect 3478 7520 3483 7576
rect 1669 7518 3483 7520
rect 1669 7515 1735 7518
rect 3417 7515 3483 7518
rect 1853 7442 1919 7445
rect 2129 7442 2195 7445
rect 1853 7440 2195 7442
rect 1853 7384 1858 7440
rect 1914 7384 2134 7440
rect 2190 7384 2195 7440
rect 1853 7382 2195 7384
rect 1853 7379 1919 7382
rect 2129 7379 2195 7382
rect 3877 7442 3943 7445
rect 13445 7442 13511 7445
rect 3877 7440 13511 7442
rect 3877 7384 3882 7440
rect 3938 7384 13450 7440
rect 13506 7384 13511 7440
rect 3877 7382 13511 7384
rect 3877 7379 3943 7382
rect 13445 7379 13511 7382
rect 2037 7306 2103 7309
rect 2221 7306 2287 7309
rect 2497 7306 2563 7309
rect 2037 7304 2146 7306
rect 2037 7248 2042 7304
rect 2098 7248 2146 7304
rect 2037 7243 2146 7248
rect 2221 7304 2563 7306
rect 2221 7248 2226 7304
rect 2282 7248 2502 7304
rect 2558 7248 2563 7304
rect 2221 7246 2563 7248
rect 2221 7243 2287 7246
rect 2497 7243 2563 7246
rect 2681 7306 2747 7309
rect 3785 7306 3851 7309
rect 13629 7306 13695 7309
rect 14000 7306 34000 7336
rect 2681 7304 3388 7306
rect 2681 7248 2686 7304
rect 2742 7248 3388 7304
rect 2681 7246 3388 7248
rect 2681 7243 2747 7246
rect 2086 7037 2146 7243
rect 3328 7173 3388 7246
rect 3785 7304 12450 7306
rect 3785 7248 3790 7304
rect 3846 7248 12450 7304
rect 3785 7246 12450 7248
rect 3785 7243 3851 7246
rect 3325 7168 3391 7173
rect 3325 7112 3330 7168
rect 3386 7112 3391 7168
rect 3325 7107 3391 7112
rect 12390 7170 12450 7246
rect 13629 7304 34000 7306
rect 13629 7248 13634 7304
rect 13690 7248 34000 7304
rect 13629 7246 34000 7248
rect 13629 7243 13695 7246
rect 14000 7216 34000 7246
rect 13813 7170 13879 7173
rect 12390 7168 13879 7170
rect 12390 7112 13818 7168
rect 13874 7112 13879 7168
rect 12390 7110 13879 7112
rect 13813 7107 13879 7110
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 5660 7104 5980 7105
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 7039 5980 7040
rect 8760 7104 9080 7105
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 7039 9080 7040
rect 2086 7032 2195 7037
rect 2086 6976 2134 7032
rect 2190 6976 2195 7032
rect 2086 6974 2195 6976
rect 2129 6971 2195 6974
rect 3141 7034 3207 7037
rect 4797 7034 4863 7037
rect 3141 7032 4863 7034
rect 3141 6976 3146 7032
rect 3202 6976 4802 7032
rect 4858 6976 4863 7032
rect 3141 6974 4863 6976
rect 3141 6971 3207 6974
rect 4797 6971 4863 6974
rect 13537 7034 13603 7037
rect 14000 7034 34000 7064
rect 13537 7032 34000 7034
rect 13537 6976 13542 7032
rect 13598 6976 34000 7032
rect 13537 6974 34000 6976
rect 13537 6971 13603 6974
rect 14000 6944 34000 6974
rect 2957 6898 3023 6901
rect 4521 6898 4587 6901
rect 5441 6898 5507 6901
rect 2957 6896 5507 6898
rect 2957 6840 2962 6896
rect 3018 6840 4526 6896
rect 4582 6840 5446 6896
rect 5502 6840 5507 6896
rect 2957 6838 5507 6840
rect 2957 6835 3023 6838
rect 4521 6835 4587 6838
rect 5441 6835 5507 6838
rect 1117 6762 1183 6765
rect 8017 6762 8083 6765
rect 1117 6760 8083 6762
rect 1117 6704 1122 6760
rect 1178 6704 8022 6760
rect 8078 6704 8083 6760
rect 1117 6702 8083 6704
rect 1117 6699 1183 6702
rect 8017 6699 8083 6702
rect 1945 6626 2011 6629
rect 3509 6626 3575 6629
rect 1945 6624 3575 6626
rect 1945 6568 1950 6624
rect 2006 6568 3514 6624
rect 3570 6568 3575 6624
rect 1945 6566 3575 6568
rect 1945 6563 2011 6566
rect 3509 6563 3575 6566
rect 13537 6626 13603 6629
rect 14000 6626 34000 6656
rect 13537 6624 34000 6626
rect 13537 6568 13542 6624
rect 13598 6568 34000 6624
rect 13537 6566 34000 6568
rect 13537 6563 13603 6566
rect 4110 6560 4430 6561
rect 4110 6496 4118 6560
rect 4182 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4430 6560
rect 4110 6495 4430 6496
rect 7210 6560 7530 6561
rect 7210 6496 7218 6560
rect 7282 6496 7298 6560
rect 7362 6496 7378 6560
rect 7442 6496 7458 6560
rect 7522 6496 7530 6560
rect 14000 6536 34000 6566
rect 7210 6495 7530 6496
rect 1853 6490 1919 6493
rect 3141 6490 3207 6493
rect 1853 6488 3207 6490
rect 1853 6432 1858 6488
rect 1914 6432 3146 6488
rect 3202 6432 3207 6488
rect 1853 6430 3207 6432
rect 1853 6427 1919 6430
rect 3141 6427 3207 6430
rect 2037 6354 2103 6357
rect 3049 6354 3115 6357
rect 4153 6354 4219 6357
rect 2037 6352 2790 6354
rect 2037 6296 2042 6352
rect 2098 6296 2790 6352
rect 2037 6294 2790 6296
rect 2037 6291 2103 6294
rect 2730 6218 2790 6294
rect 3049 6352 4219 6354
rect 3049 6296 3054 6352
rect 3110 6296 4158 6352
rect 4214 6296 4219 6352
rect 3049 6294 4219 6296
rect 3049 6291 3115 6294
rect 4153 6291 4219 6294
rect 4429 6354 4495 6357
rect 6453 6354 6519 6357
rect 4429 6352 6519 6354
rect 4429 6296 4434 6352
rect 4490 6296 6458 6352
rect 6514 6296 6519 6352
rect 4429 6294 6519 6296
rect 4429 6291 4495 6294
rect 6453 6291 6519 6294
rect 13721 6354 13787 6357
rect 14000 6354 34000 6384
rect 13721 6352 34000 6354
rect 13721 6296 13726 6352
rect 13782 6296 34000 6352
rect 13721 6294 34000 6296
rect 13721 6291 13787 6294
rect 14000 6264 34000 6294
rect 7005 6218 7071 6221
rect 2730 6216 7071 6218
rect 2730 6160 7010 6216
rect 7066 6160 7071 6216
rect 2730 6158 7071 6160
rect 7005 6155 7071 6158
rect 3693 6082 3759 6085
rect 4153 6082 4219 6085
rect 3693 6080 4219 6082
rect 3693 6024 3698 6080
rect 3754 6024 4158 6080
rect 4214 6024 4219 6080
rect 3693 6022 4219 6024
rect 3693 6019 3759 6022
rect 4153 6019 4219 6022
rect 13813 6082 13879 6085
rect 14000 6082 34000 6112
rect 13813 6080 34000 6082
rect 13813 6024 13818 6080
rect 13874 6024 34000 6080
rect 13813 6022 34000 6024
rect 13813 6019 13879 6022
rect 5660 6016 5980 6017
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 5951 5980 5952
rect 8760 6016 9080 6017
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 14000 5992 34000 6022
rect 8760 5951 9080 5952
rect 1025 5946 1091 5949
rect 4429 5946 4495 5949
rect 1025 5944 4495 5946
rect 1025 5888 1030 5944
rect 1086 5888 4434 5944
rect 4490 5888 4495 5944
rect 1025 5886 4495 5888
rect 1025 5883 1091 5886
rect 4429 5883 4495 5886
rect 3325 5810 3391 5813
rect 5165 5810 5231 5813
rect 5349 5810 5415 5813
rect 3325 5808 5415 5810
rect 3325 5752 3330 5808
rect 3386 5752 5170 5808
rect 5226 5752 5354 5808
rect 5410 5752 5415 5808
rect 3325 5750 5415 5752
rect 3325 5747 3391 5750
rect 5165 5747 5231 5750
rect 5349 5747 5415 5750
rect 5901 5810 5967 5813
rect 6637 5810 6703 5813
rect 5901 5808 6703 5810
rect 5901 5752 5906 5808
rect 5962 5752 6642 5808
rect 6698 5752 6703 5808
rect 5901 5750 6703 5752
rect 5901 5747 5967 5750
rect 6637 5747 6703 5750
rect 3141 5674 3207 5677
rect 5717 5674 5783 5677
rect 3141 5672 5783 5674
rect 3141 5616 3146 5672
rect 3202 5616 5722 5672
rect 5778 5616 5783 5672
rect 3141 5614 5783 5616
rect 3141 5611 3207 5614
rect 5717 5611 5783 5614
rect 6913 5674 6979 5677
rect 14000 5674 34000 5704
rect 6913 5672 34000 5674
rect 6913 5616 6918 5672
rect 6974 5616 34000 5672
rect 6913 5614 34000 5616
rect 6913 5611 6979 5614
rect 14000 5584 34000 5614
rect 4110 5472 4430 5473
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 5407 4430 5408
rect 7210 5472 7530 5473
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 5407 7530 5408
rect 14000 5402 34000 5432
rect 12390 5342 34000 5402
rect 2589 5266 2655 5269
rect 12390 5266 12450 5342
rect 14000 5312 34000 5342
rect 2589 5264 12450 5266
rect 2589 5208 2594 5264
rect 2650 5208 12450 5264
rect 2589 5206 12450 5208
rect 2589 5203 2655 5206
rect 2497 5130 2563 5133
rect 8201 5130 8267 5133
rect 8569 5130 8635 5133
rect 2497 5128 8635 5130
rect 2497 5072 2502 5128
rect 2558 5072 8206 5128
rect 8262 5072 8574 5128
rect 8630 5072 8635 5128
rect 2497 5070 8635 5072
rect 2497 5067 2563 5070
rect 8201 5067 8267 5070
rect 8569 5067 8635 5070
rect 13629 4994 13695 4997
rect 14000 4994 34000 5024
rect 13629 4992 34000 4994
rect 13629 4936 13634 4992
rect 13690 4936 34000 4992
rect 13629 4934 34000 4936
rect 13629 4931 13695 4934
rect 5660 4928 5980 4929
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 4863 5980 4864
rect 8760 4928 9080 4929
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 14000 4904 34000 4934
rect 8760 4863 9080 4864
rect 4613 4722 4679 4725
rect 14000 4722 34000 4752
rect 4613 4720 34000 4722
rect 4613 4664 4618 4720
rect 4674 4664 34000 4720
rect 4613 4662 34000 4664
rect 4613 4659 4679 4662
rect 14000 4632 34000 4662
rect 9581 4586 9647 4589
rect 9581 4584 12450 4586
rect 9581 4528 9586 4584
rect 9642 4528 12450 4584
rect 9581 4526 12450 4528
rect 9581 4523 9647 4526
rect 2681 4450 2747 4453
rect 2484 4448 2747 4450
rect 2484 4392 2686 4448
rect 2742 4392 2747 4448
rect 2484 4390 2747 4392
rect 12390 4450 12450 4526
rect 14000 4450 34000 4480
rect 12390 4390 34000 4450
rect 2681 4387 2747 4390
rect 4110 4384 4430 4385
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 4319 4430 4320
rect 7210 4384 7530 4385
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 14000 4360 34000 4390
rect 7210 4319 7530 4320
rect 4705 4042 4771 4045
rect 14000 4042 34000 4072
rect 4705 4040 34000 4042
rect 4705 3984 4710 4040
rect 4766 3984 34000 4040
rect 4705 3982 34000 3984
rect 4705 3979 4771 3982
rect 14000 3952 34000 3982
rect 5660 3840 5980 3841
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 3775 5980 3776
rect 8760 3840 9080 3841
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 3775 9080 3776
rect 13445 3770 13511 3773
rect 14000 3770 34000 3800
rect 13445 3768 34000 3770
rect 13445 3712 13450 3768
rect 13506 3712 34000 3768
rect 13445 3710 34000 3712
rect 13445 3707 13511 3710
rect 14000 3680 34000 3710
rect 7925 3634 7991 3637
rect 8201 3634 8267 3637
rect 7925 3632 8267 3634
rect 7925 3576 7930 3632
rect 7986 3576 8206 3632
rect 8262 3576 8267 3632
rect 7925 3574 8267 3576
rect 7925 3571 7991 3574
rect 8201 3571 8267 3574
rect 5625 3498 5691 3501
rect 8293 3498 8359 3501
rect 5625 3496 8359 3498
rect 5625 3440 5630 3496
rect 5686 3440 8298 3496
rect 8354 3440 8359 3496
rect 5625 3438 8359 3440
rect 5625 3435 5691 3438
rect 8293 3435 8359 3438
rect 13261 3362 13327 3365
rect 14000 3362 34000 3392
rect 13261 3360 34000 3362
rect 13261 3304 13266 3360
rect 13322 3304 34000 3360
rect 13261 3302 34000 3304
rect 13261 3299 13327 3302
rect 4110 3296 4430 3297
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 3231 4430 3232
rect 7210 3296 7530 3297
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 14000 3272 34000 3302
rect 7210 3231 7530 3232
rect 14000 3088 34000 3120
rect 14000 3032 22466 3088
rect 22522 3032 34000 3088
rect 14000 3000 34000 3032
rect 6269 2954 6335 2957
rect 6821 2954 6887 2957
rect 6269 2952 6887 2954
rect 6269 2896 6274 2952
rect 6330 2896 6826 2952
rect 6882 2896 6887 2952
rect 6269 2894 6887 2896
rect 6269 2891 6335 2894
rect 6821 2891 6887 2894
rect 14000 2816 34000 2848
rect 14000 2760 22190 2816
rect 22246 2760 34000 2816
rect 5660 2752 5980 2753
rect 5660 2688 5668 2752
rect 5732 2688 5748 2752
rect 5812 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5980 2752
rect 5660 2687 5980 2688
rect 8760 2752 9080 2753
rect 8760 2688 8768 2752
rect 8832 2688 8848 2752
rect 8912 2688 8928 2752
rect 8992 2688 9008 2752
rect 9072 2688 9080 2752
rect 14000 2728 34000 2760
rect 8760 2687 9080 2688
rect 14000 2408 34000 2440
rect 14000 2352 22282 2408
rect 22338 2352 34000 2408
rect 14000 2320 34000 2352
rect 4110 2208 4430 2209
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 2143 4430 2144
rect 7210 2208 7530 2209
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 2143 7530 2144
rect 14000 2136 34000 2168
rect 14000 2080 22742 2136
rect 22798 2080 34000 2136
rect 14000 2048 34000 2080
rect 14000 1728 34000 1760
rect 14000 1672 22374 1728
rect 22430 1672 34000 1728
rect 14000 1640 34000 1672
rect 4705 1458 4771 1461
rect 14000 1458 34000 1488
rect 4705 1456 34000 1458
rect 4705 1400 4710 1456
rect 4766 1400 34000 1456
rect 4705 1398 34000 1400
rect 4705 1395 4771 1398
rect 14000 1368 34000 1398
rect 14000 1184 34000 1216
rect 14000 1128 19798 1184
rect 19854 1128 34000 1184
rect 14000 1096 34000 1128
rect 9305 778 9371 781
rect 14000 778 34000 808
rect 9305 776 34000 778
rect 9305 720 9310 776
rect 9366 720 34000 776
rect 9305 718 34000 720
rect 9305 715 9371 718
rect 14000 688 34000 718
rect 3417 506 3483 509
rect 14000 506 34000 536
rect 3417 504 34000 506
rect 3417 448 3422 504
rect 3478 448 34000 504
rect 3417 446 34000 448
rect 3417 443 3483 446
rect 14000 416 34000 446
rect 3969 234 4035 237
rect 14000 234 34000 264
rect 3969 232 34000 234
rect 3969 176 3974 232
rect 4030 176 34000 232
rect 3969 174 34000 176
rect 3969 171 4035 174
rect 14000 144 34000 174
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 5668 11452 5732 11456
rect 5668 11396 5672 11452
rect 5672 11396 5728 11452
rect 5728 11396 5732 11452
rect 5668 11392 5732 11396
rect 5748 11452 5812 11456
rect 5748 11396 5752 11452
rect 5752 11396 5808 11452
rect 5808 11396 5812 11452
rect 5748 11392 5812 11396
rect 5828 11452 5892 11456
rect 5828 11396 5832 11452
rect 5832 11396 5888 11452
rect 5888 11396 5892 11452
rect 5828 11392 5892 11396
rect 5908 11452 5972 11456
rect 5908 11396 5912 11452
rect 5912 11396 5968 11452
rect 5968 11396 5972 11452
rect 5908 11392 5972 11396
rect 8768 11452 8832 11456
rect 8768 11396 8772 11452
rect 8772 11396 8828 11452
rect 8828 11396 8832 11452
rect 8768 11392 8832 11396
rect 8848 11452 8912 11456
rect 8848 11396 8852 11452
rect 8852 11396 8908 11452
rect 8908 11396 8912 11452
rect 8848 11392 8912 11396
rect 8928 11452 8992 11456
rect 8928 11396 8932 11452
rect 8932 11396 8988 11452
rect 8988 11396 8992 11452
rect 8928 11392 8992 11396
rect 9008 11452 9072 11456
rect 9008 11396 9012 11452
rect 9012 11396 9068 11452
rect 9068 11396 9072 11452
rect 9008 11392 9072 11396
rect 4118 10908 4182 10912
rect 4118 10852 4122 10908
rect 4122 10852 4178 10908
rect 4178 10852 4182 10908
rect 4118 10848 4182 10852
rect 4198 10908 4262 10912
rect 4198 10852 4202 10908
rect 4202 10852 4258 10908
rect 4258 10852 4262 10908
rect 4198 10848 4262 10852
rect 4278 10908 4342 10912
rect 4278 10852 4282 10908
rect 4282 10852 4338 10908
rect 4338 10852 4342 10908
rect 4278 10848 4342 10852
rect 4358 10908 4422 10912
rect 4358 10852 4362 10908
rect 4362 10852 4418 10908
rect 4418 10852 4422 10908
rect 4358 10848 4422 10852
rect 7218 10908 7282 10912
rect 7218 10852 7222 10908
rect 7222 10852 7278 10908
rect 7278 10852 7282 10908
rect 7218 10848 7282 10852
rect 7298 10908 7362 10912
rect 7298 10852 7302 10908
rect 7302 10852 7358 10908
rect 7358 10852 7362 10908
rect 7298 10848 7362 10852
rect 7378 10908 7442 10912
rect 7378 10852 7382 10908
rect 7382 10852 7438 10908
rect 7438 10852 7442 10908
rect 7378 10848 7442 10852
rect 7458 10908 7522 10912
rect 7458 10852 7462 10908
rect 7462 10852 7518 10908
rect 7518 10852 7522 10908
rect 7458 10848 7522 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 5668 10364 5732 10368
rect 5668 10308 5672 10364
rect 5672 10308 5728 10364
rect 5728 10308 5732 10364
rect 5668 10304 5732 10308
rect 5748 10364 5812 10368
rect 5748 10308 5752 10364
rect 5752 10308 5808 10364
rect 5808 10308 5812 10364
rect 5748 10304 5812 10308
rect 5828 10364 5892 10368
rect 5828 10308 5832 10364
rect 5832 10308 5888 10364
rect 5888 10308 5892 10364
rect 5828 10304 5892 10308
rect 5908 10364 5972 10368
rect 5908 10308 5912 10364
rect 5912 10308 5968 10364
rect 5968 10308 5972 10364
rect 5908 10304 5972 10308
rect 8768 10364 8832 10368
rect 8768 10308 8772 10364
rect 8772 10308 8828 10364
rect 8828 10308 8832 10364
rect 8768 10304 8832 10308
rect 8848 10364 8912 10368
rect 8848 10308 8852 10364
rect 8852 10308 8908 10364
rect 8908 10308 8912 10364
rect 8848 10304 8912 10308
rect 8928 10364 8992 10368
rect 8928 10308 8932 10364
rect 8932 10308 8988 10364
rect 8988 10308 8992 10364
rect 8928 10304 8992 10308
rect 9008 10364 9072 10368
rect 9008 10308 9012 10364
rect 9012 10308 9068 10364
rect 9068 10308 9072 10364
rect 9008 10304 9072 10308
rect 4118 9820 4182 9824
rect 4118 9764 4122 9820
rect 4122 9764 4178 9820
rect 4178 9764 4182 9820
rect 4118 9760 4182 9764
rect 4198 9820 4262 9824
rect 4198 9764 4202 9820
rect 4202 9764 4258 9820
rect 4258 9764 4262 9820
rect 4198 9760 4262 9764
rect 4278 9820 4342 9824
rect 4278 9764 4282 9820
rect 4282 9764 4338 9820
rect 4338 9764 4342 9820
rect 4278 9760 4342 9764
rect 4358 9820 4422 9824
rect 4358 9764 4362 9820
rect 4362 9764 4418 9820
rect 4418 9764 4422 9820
rect 4358 9760 4422 9764
rect 7218 9820 7282 9824
rect 7218 9764 7222 9820
rect 7222 9764 7278 9820
rect 7278 9764 7282 9820
rect 7218 9760 7282 9764
rect 7298 9820 7362 9824
rect 7298 9764 7302 9820
rect 7302 9764 7358 9820
rect 7358 9764 7362 9820
rect 7298 9760 7362 9764
rect 7378 9820 7442 9824
rect 7378 9764 7382 9820
rect 7382 9764 7438 9820
rect 7438 9764 7442 9820
rect 7378 9760 7442 9764
rect 7458 9820 7522 9824
rect 7458 9764 7462 9820
rect 7462 9764 7518 9820
rect 7518 9764 7522 9820
rect 7458 9760 7522 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 5668 9276 5732 9280
rect 5668 9220 5672 9276
rect 5672 9220 5728 9276
rect 5728 9220 5732 9276
rect 5668 9216 5732 9220
rect 5748 9276 5812 9280
rect 5748 9220 5752 9276
rect 5752 9220 5808 9276
rect 5808 9220 5812 9276
rect 5748 9216 5812 9220
rect 5828 9276 5892 9280
rect 5828 9220 5832 9276
rect 5832 9220 5888 9276
rect 5888 9220 5892 9276
rect 5828 9216 5892 9220
rect 5908 9276 5972 9280
rect 5908 9220 5912 9276
rect 5912 9220 5968 9276
rect 5968 9220 5972 9276
rect 5908 9216 5972 9220
rect 8768 9276 8832 9280
rect 8768 9220 8772 9276
rect 8772 9220 8828 9276
rect 8828 9220 8832 9276
rect 8768 9216 8832 9220
rect 8848 9276 8912 9280
rect 8848 9220 8852 9276
rect 8852 9220 8908 9276
rect 8908 9220 8912 9276
rect 8848 9216 8912 9220
rect 8928 9276 8992 9280
rect 8928 9220 8932 9276
rect 8932 9220 8988 9276
rect 8988 9220 8992 9276
rect 8928 9216 8992 9220
rect 9008 9276 9072 9280
rect 9008 9220 9012 9276
rect 9012 9220 9068 9276
rect 9068 9220 9072 9276
rect 9008 9216 9072 9220
rect 4118 8732 4182 8736
rect 4118 8676 4122 8732
rect 4122 8676 4178 8732
rect 4178 8676 4182 8732
rect 4118 8672 4182 8676
rect 4198 8732 4262 8736
rect 4198 8676 4202 8732
rect 4202 8676 4258 8732
rect 4258 8676 4262 8732
rect 4198 8672 4262 8676
rect 4278 8732 4342 8736
rect 4278 8676 4282 8732
rect 4282 8676 4338 8732
rect 4338 8676 4342 8732
rect 4278 8672 4342 8676
rect 4358 8732 4422 8736
rect 4358 8676 4362 8732
rect 4362 8676 4418 8732
rect 4418 8676 4422 8732
rect 4358 8672 4422 8676
rect 7218 8732 7282 8736
rect 7218 8676 7222 8732
rect 7222 8676 7278 8732
rect 7278 8676 7282 8732
rect 7218 8672 7282 8676
rect 7298 8732 7362 8736
rect 7298 8676 7302 8732
rect 7302 8676 7358 8732
rect 7358 8676 7362 8732
rect 7298 8672 7362 8676
rect 7378 8732 7442 8736
rect 7378 8676 7382 8732
rect 7382 8676 7438 8732
rect 7438 8676 7442 8732
rect 7378 8672 7442 8676
rect 7458 8732 7522 8736
rect 7458 8676 7462 8732
rect 7462 8676 7518 8732
rect 7518 8676 7522 8732
rect 7458 8672 7522 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 5668 8188 5732 8192
rect 5668 8132 5672 8188
rect 5672 8132 5728 8188
rect 5728 8132 5732 8188
rect 5668 8128 5732 8132
rect 5748 8188 5812 8192
rect 5748 8132 5752 8188
rect 5752 8132 5808 8188
rect 5808 8132 5812 8188
rect 5748 8128 5812 8132
rect 5828 8188 5892 8192
rect 5828 8132 5832 8188
rect 5832 8132 5888 8188
rect 5888 8132 5892 8188
rect 5828 8128 5892 8132
rect 5908 8188 5972 8192
rect 5908 8132 5912 8188
rect 5912 8132 5968 8188
rect 5968 8132 5972 8188
rect 5908 8128 5972 8132
rect 8768 8188 8832 8192
rect 8768 8132 8772 8188
rect 8772 8132 8828 8188
rect 8828 8132 8832 8188
rect 8768 8128 8832 8132
rect 8848 8188 8912 8192
rect 8848 8132 8852 8188
rect 8852 8132 8908 8188
rect 8908 8132 8912 8188
rect 8848 8128 8912 8132
rect 8928 8188 8992 8192
rect 8928 8132 8932 8188
rect 8932 8132 8988 8188
rect 8988 8132 8992 8188
rect 8928 8128 8992 8132
rect 9008 8188 9072 8192
rect 9008 8132 9012 8188
rect 9012 8132 9068 8188
rect 9068 8132 9072 8188
rect 9008 8128 9072 8132
rect 4118 7644 4182 7648
rect 4118 7588 4122 7644
rect 4122 7588 4178 7644
rect 4178 7588 4182 7644
rect 4118 7584 4182 7588
rect 4198 7644 4262 7648
rect 4198 7588 4202 7644
rect 4202 7588 4258 7644
rect 4258 7588 4262 7644
rect 4198 7584 4262 7588
rect 4278 7644 4342 7648
rect 4278 7588 4282 7644
rect 4282 7588 4338 7644
rect 4338 7588 4342 7644
rect 4278 7584 4342 7588
rect 4358 7644 4422 7648
rect 4358 7588 4362 7644
rect 4362 7588 4418 7644
rect 4418 7588 4422 7644
rect 4358 7584 4422 7588
rect 7218 7644 7282 7648
rect 7218 7588 7222 7644
rect 7222 7588 7278 7644
rect 7278 7588 7282 7644
rect 7218 7584 7282 7588
rect 7298 7644 7362 7648
rect 7298 7588 7302 7644
rect 7302 7588 7358 7644
rect 7358 7588 7362 7644
rect 7298 7584 7362 7588
rect 7378 7644 7442 7648
rect 7378 7588 7382 7644
rect 7382 7588 7438 7644
rect 7438 7588 7442 7644
rect 7378 7584 7442 7588
rect 7458 7644 7522 7648
rect 7458 7588 7462 7644
rect 7462 7588 7518 7644
rect 7518 7588 7522 7644
rect 7458 7584 7522 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 5668 7100 5732 7104
rect 5668 7044 5672 7100
rect 5672 7044 5728 7100
rect 5728 7044 5732 7100
rect 5668 7040 5732 7044
rect 5748 7100 5812 7104
rect 5748 7044 5752 7100
rect 5752 7044 5808 7100
rect 5808 7044 5812 7100
rect 5748 7040 5812 7044
rect 5828 7100 5892 7104
rect 5828 7044 5832 7100
rect 5832 7044 5888 7100
rect 5888 7044 5892 7100
rect 5828 7040 5892 7044
rect 5908 7100 5972 7104
rect 5908 7044 5912 7100
rect 5912 7044 5968 7100
rect 5968 7044 5972 7100
rect 5908 7040 5972 7044
rect 8768 7100 8832 7104
rect 8768 7044 8772 7100
rect 8772 7044 8828 7100
rect 8828 7044 8832 7100
rect 8768 7040 8832 7044
rect 8848 7100 8912 7104
rect 8848 7044 8852 7100
rect 8852 7044 8908 7100
rect 8908 7044 8912 7100
rect 8848 7040 8912 7044
rect 8928 7100 8992 7104
rect 8928 7044 8932 7100
rect 8932 7044 8988 7100
rect 8988 7044 8992 7100
rect 8928 7040 8992 7044
rect 9008 7100 9072 7104
rect 9008 7044 9012 7100
rect 9012 7044 9068 7100
rect 9068 7044 9072 7100
rect 9008 7040 9072 7044
rect 4118 6556 4182 6560
rect 4118 6500 4122 6556
rect 4122 6500 4178 6556
rect 4178 6500 4182 6556
rect 4118 6496 4182 6500
rect 4198 6556 4262 6560
rect 4198 6500 4202 6556
rect 4202 6500 4258 6556
rect 4258 6500 4262 6556
rect 4198 6496 4262 6500
rect 4278 6556 4342 6560
rect 4278 6500 4282 6556
rect 4282 6500 4338 6556
rect 4338 6500 4342 6556
rect 4278 6496 4342 6500
rect 4358 6556 4422 6560
rect 4358 6500 4362 6556
rect 4362 6500 4418 6556
rect 4418 6500 4422 6556
rect 4358 6496 4422 6500
rect 7218 6556 7282 6560
rect 7218 6500 7222 6556
rect 7222 6500 7278 6556
rect 7278 6500 7282 6556
rect 7218 6496 7282 6500
rect 7298 6556 7362 6560
rect 7298 6500 7302 6556
rect 7302 6500 7358 6556
rect 7358 6500 7362 6556
rect 7298 6496 7362 6500
rect 7378 6556 7442 6560
rect 7378 6500 7382 6556
rect 7382 6500 7438 6556
rect 7438 6500 7442 6556
rect 7378 6496 7442 6500
rect 7458 6556 7522 6560
rect 7458 6500 7462 6556
rect 7462 6500 7518 6556
rect 7518 6500 7522 6556
rect 7458 6496 7522 6500
rect 5668 6012 5732 6016
rect 5668 5956 5672 6012
rect 5672 5956 5728 6012
rect 5728 5956 5732 6012
rect 5668 5952 5732 5956
rect 5748 6012 5812 6016
rect 5748 5956 5752 6012
rect 5752 5956 5808 6012
rect 5808 5956 5812 6012
rect 5748 5952 5812 5956
rect 5828 6012 5892 6016
rect 5828 5956 5832 6012
rect 5832 5956 5888 6012
rect 5888 5956 5892 6012
rect 5828 5952 5892 5956
rect 5908 6012 5972 6016
rect 5908 5956 5912 6012
rect 5912 5956 5968 6012
rect 5968 5956 5972 6012
rect 5908 5952 5972 5956
rect 8768 6012 8832 6016
rect 8768 5956 8772 6012
rect 8772 5956 8828 6012
rect 8828 5956 8832 6012
rect 8768 5952 8832 5956
rect 8848 6012 8912 6016
rect 8848 5956 8852 6012
rect 8852 5956 8908 6012
rect 8908 5956 8912 6012
rect 8848 5952 8912 5956
rect 8928 6012 8992 6016
rect 8928 5956 8932 6012
rect 8932 5956 8988 6012
rect 8988 5956 8992 6012
rect 8928 5952 8992 5956
rect 9008 6012 9072 6016
rect 9008 5956 9012 6012
rect 9012 5956 9068 6012
rect 9068 5956 9072 6012
rect 9008 5952 9072 5956
rect 4118 5468 4182 5472
rect 4118 5412 4122 5468
rect 4122 5412 4178 5468
rect 4178 5412 4182 5468
rect 4118 5408 4182 5412
rect 4198 5468 4262 5472
rect 4198 5412 4202 5468
rect 4202 5412 4258 5468
rect 4258 5412 4262 5468
rect 4198 5408 4262 5412
rect 4278 5468 4342 5472
rect 4278 5412 4282 5468
rect 4282 5412 4338 5468
rect 4338 5412 4342 5468
rect 4278 5408 4342 5412
rect 4358 5468 4422 5472
rect 4358 5412 4362 5468
rect 4362 5412 4418 5468
rect 4418 5412 4422 5468
rect 4358 5408 4422 5412
rect 7218 5468 7282 5472
rect 7218 5412 7222 5468
rect 7222 5412 7278 5468
rect 7278 5412 7282 5468
rect 7218 5408 7282 5412
rect 7298 5468 7362 5472
rect 7298 5412 7302 5468
rect 7302 5412 7358 5468
rect 7358 5412 7362 5468
rect 7298 5408 7362 5412
rect 7378 5468 7442 5472
rect 7378 5412 7382 5468
rect 7382 5412 7438 5468
rect 7438 5412 7442 5468
rect 7378 5408 7442 5412
rect 7458 5468 7522 5472
rect 7458 5412 7462 5468
rect 7462 5412 7518 5468
rect 7518 5412 7522 5468
rect 7458 5408 7522 5412
rect 5668 4924 5732 4928
rect 5668 4868 5672 4924
rect 5672 4868 5728 4924
rect 5728 4868 5732 4924
rect 5668 4864 5732 4868
rect 5748 4924 5812 4928
rect 5748 4868 5752 4924
rect 5752 4868 5808 4924
rect 5808 4868 5812 4924
rect 5748 4864 5812 4868
rect 5828 4924 5892 4928
rect 5828 4868 5832 4924
rect 5832 4868 5888 4924
rect 5888 4868 5892 4924
rect 5828 4864 5892 4868
rect 5908 4924 5972 4928
rect 5908 4868 5912 4924
rect 5912 4868 5968 4924
rect 5968 4868 5972 4924
rect 5908 4864 5972 4868
rect 8768 4924 8832 4928
rect 8768 4868 8772 4924
rect 8772 4868 8828 4924
rect 8828 4868 8832 4924
rect 8768 4864 8832 4868
rect 8848 4924 8912 4928
rect 8848 4868 8852 4924
rect 8852 4868 8908 4924
rect 8908 4868 8912 4924
rect 8848 4864 8912 4868
rect 8928 4924 8992 4928
rect 8928 4868 8932 4924
rect 8932 4868 8988 4924
rect 8988 4868 8992 4924
rect 8928 4864 8992 4868
rect 9008 4924 9072 4928
rect 9008 4868 9012 4924
rect 9012 4868 9068 4924
rect 9068 4868 9072 4924
rect 9008 4864 9072 4868
rect 4118 4380 4182 4384
rect 4118 4324 4122 4380
rect 4122 4324 4178 4380
rect 4178 4324 4182 4380
rect 4118 4320 4182 4324
rect 4198 4380 4262 4384
rect 4198 4324 4202 4380
rect 4202 4324 4258 4380
rect 4258 4324 4262 4380
rect 4198 4320 4262 4324
rect 4278 4380 4342 4384
rect 4278 4324 4282 4380
rect 4282 4324 4338 4380
rect 4338 4324 4342 4380
rect 4278 4320 4342 4324
rect 4358 4380 4422 4384
rect 4358 4324 4362 4380
rect 4362 4324 4418 4380
rect 4418 4324 4422 4380
rect 4358 4320 4422 4324
rect 7218 4380 7282 4384
rect 7218 4324 7222 4380
rect 7222 4324 7278 4380
rect 7278 4324 7282 4380
rect 7218 4320 7282 4324
rect 7298 4380 7362 4384
rect 7298 4324 7302 4380
rect 7302 4324 7358 4380
rect 7358 4324 7362 4380
rect 7298 4320 7362 4324
rect 7378 4380 7442 4384
rect 7378 4324 7382 4380
rect 7382 4324 7438 4380
rect 7438 4324 7442 4380
rect 7378 4320 7442 4324
rect 7458 4380 7522 4384
rect 7458 4324 7462 4380
rect 7462 4324 7518 4380
rect 7518 4324 7522 4380
rect 7458 4320 7522 4324
rect 5668 3836 5732 3840
rect 5668 3780 5672 3836
rect 5672 3780 5728 3836
rect 5728 3780 5732 3836
rect 5668 3776 5732 3780
rect 5748 3836 5812 3840
rect 5748 3780 5752 3836
rect 5752 3780 5808 3836
rect 5808 3780 5812 3836
rect 5748 3776 5812 3780
rect 5828 3836 5892 3840
rect 5828 3780 5832 3836
rect 5832 3780 5888 3836
rect 5888 3780 5892 3836
rect 5828 3776 5892 3780
rect 5908 3836 5972 3840
rect 5908 3780 5912 3836
rect 5912 3780 5968 3836
rect 5968 3780 5972 3836
rect 5908 3776 5972 3780
rect 8768 3836 8832 3840
rect 8768 3780 8772 3836
rect 8772 3780 8828 3836
rect 8828 3780 8832 3836
rect 8768 3776 8832 3780
rect 8848 3836 8912 3840
rect 8848 3780 8852 3836
rect 8852 3780 8908 3836
rect 8908 3780 8912 3836
rect 8848 3776 8912 3780
rect 8928 3836 8992 3840
rect 8928 3780 8932 3836
rect 8932 3780 8988 3836
rect 8988 3780 8992 3836
rect 8928 3776 8992 3780
rect 9008 3836 9072 3840
rect 9008 3780 9012 3836
rect 9012 3780 9068 3836
rect 9068 3780 9072 3836
rect 9008 3776 9072 3780
rect 4118 3292 4182 3296
rect 4118 3236 4122 3292
rect 4122 3236 4178 3292
rect 4178 3236 4182 3292
rect 4118 3232 4182 3236
rect 4198 3292 4262 3296
rect 4198 3236 4202 3292
rect 4202 3236 4258 3292
rect 4258 3236 4262 3292
rect 4198 3232 4262 3236
rect 4278 3292 4342 3296
rect 4278 3236 4282 3292
rect 4282 3236 4338 3292
rect 4338 3236 4342 3292
rect 4278 3232 4342 3236
rect 4358 3292 4422 3296
rect 4358 3236 4362 3292
rect 4362 3236 4418 3292
rect 4418 3236 4422 3292
rect 4358 3232 4422 3236
rect 7218 3292 7282 3296
rect 7218 3236 7222 3292
rect 7222 3236 7278 3292
rect 7278 3236 7282 3292
rect 7218 3232 7282 3236
rect 7298 3292 7362 3296
rect 7298 3236 7302 3292
rect 7302 3236 7358 3292
rect 7358 3236 7362 3292
rect 7298 3232 7362 3236
rect 7378 3292 7442 3296
rect 7378 3236 7382 3292
rect 7382 3236 7438 3292
rect 7438 3236 7442 3292
rect 7378 3232 7442 3236
rect 7458 3292 7522 3296
rect 7458 3236 7462 3292
rect 7462 3236 7518 3292
rect 7518 3236 7522 3292
rect 7458 3232 7522 3236
rect 5668 2748 5732 2752
rect 5668 2692 5672 2748
rect 5672 2692 5728 2748
rect 5728 2692 5732 2748
rect 5668 2688 5732 2692
rect 5748 2748 5812 2752
rect 5748 2692 5752 2748
rect 5752 2692 5808 2748
rect 5808 2692 5812 2748
rect 5748 2688 5812 2692
rect 5828 2748 5892 2752
rect 5828 2692 5832 2748
rect 5832 2692 5888 2748
rect 5888 2692 5892 2748
rect 5828 2688 5892 2692
rect 5908 2748 5972 2752
rect 5908 2692 5912 2748
rect 5912 2692 5968 2748
rect 5968 2692 5972 2748
rect 5908 2688 5972 2692
rect 8768 2748 8832 2752
rect 8768 2692 8772 2748
rect 8772 2692 8828 2748
rect 8828 2692 8832 2748
rect 8768 2688 8832 2692
rect 8848 2748 8912 2752
rect 8848 2692 8852 2748
rect 8852 2692 8908 2748
rect 8908 2692 8912 2748
rect 8848 2688 8912 2692
rect 8928 2748 8992 2752
rect 8928 2692 8932 2748
rect 8932 2692 8988 2748
rect 8988 2692 8992 2748
rect 8928 2688 8992 2692
rect 9008 2748 9072 2752
rect 9008 2692 9012 2748
rect 9012 2692 9068 2748
rect 9068 2692 9072 2748
rect 9008 2688 9072 2692
rect 4118 2204 4182 2208
rect 4118 2148 4122 2204
rect 4122 2148 4178 2204
rect 4178 2148 4182 2204
rect 4118 2144 4182 2148
rect 4198 2204 4262 2208
rect 4198 2148 4202 2204
rect 4202 2148 4258 2204
rect 4258 2148 4262 2204
rect 4198 2144 4262 2148
rect 4278 2204 4342 2208
rect 4278 2148 4282 2204
rect 4282 2148 4338 2204
rect 4338 2148 4342 2204
rect 4278 2144 4342 2148
rect 4358 2204 4422 2208
rect 4358 2148 4362 2204
rect 4362 2148 4418 2204
rect 4418 2148 4422 2204
rect 4358 2144 4422 2148
rect 7218 2204 7282 2208
rect 7218 2148 7222 2204
rect 7222 2148 7278 2204
rect 7278 2148 7282 2204
rect 7218 2144 7282 2148
rect 7298 2204 7362 2208
rect 7298 2148 7302 2204
rect 7302 2148 7358 2204
rect 7358 2148 7362 2204
rect 7298 2144 7362 2148
rect 7378 2204 7442 2208
rect 7378 2148 7382 2204
rect 7382 2148 7438 2204
rect 7438 2148 7442 2204
rect 7378 2144 7442 2148
rect 7458 2204 7522 2208
rect 7458 2148 7462 2204
rect 7462 2148 7518 2204
rect 7518 2148 7522 2204
rect 7458 2144 7522 2148
<< metal4 >>
rect -1620 13922 -1300 13964
rect -1620 13686 -1578 13922
rect -1342 13686 -1300 13922
rect -1620 8244 -1300 13686
rect 12064 13922 12384 13964
rect 12064 13686 12106 13922
rect 12342 13686 12384 13922
rect -1620 8008 -1578 8244
rect -1342 8008 -1300 8244
rect -1620 5144 -1300 8008
rect -1620 4908 -1578 5144
rect -1342 4908 -1300 5144
rect -1620 -86 -1300 4908
rect -960 13262 -640 13304
rect -960 13026 -918 13262
rect -682 13026 -640 13262
rect -960 9794 -640 13026
rect 11404 13262 11724 13304
rect 11404 13026 11446 13262
rect 11682 13026 11724 13262
rect -960 9558 -918 9794
rect -682 9558 -640 9794
rect -960 6694 -640 9558
rect -960 6458 -918 6694
rect -682 6458 -640 6694
rect -960 3594 -640 6458
rect -960 3358 -918 3594
rect -682 3358 -640 3594
rect -960 574 -640 3358
rect -300 12602 20 12644
rect -300 12366 -258 12602
rect -22 12366 20 12602
rect -300 10444 20 12366
rect -300 10208 -258 10444
rect -22 10208 20 10444
rect -300 7344 20 10208
rect -300 7108 -258 7344
rect -22 7108 20 7344
rect -300 4244 20 7108
rect -300 4008 -258 4244
rect -22 4008 20 4244
rect -300 1234 20 4008
rect 360 11942 680 11984
rect 360 11706 402 11942
rect 638 11706 680 11942
rect 360 8894 680 11706
rect 360 8658 402 8894
rect 638 8658 680 8894
rect 360 5794 680 8658
rect 360 5558 402 5794
rect 638 5558 680 5794
rect 360 2694 680 5558
rect 2560 11942 2880 12644
rect 2560 11706 2602 11942
rect 2838 11706 2880 11942
rect 2560 11456 2880 11706
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8894 2880 9216
rect 2560 8658 2602 8894
rect 2838 8658 2880 8894
rect 2560 8192 2880 8658
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 7104 2880 8128
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 5794 2880 7040
rect 2560 5558 2602 5794
rect 2838 5558 2880 5794
rect 1996 5144 2276 5186
rect 1996 4908 2018 5144
rect 2254 4908 2276 5144
rect 1996 4866 2276 4908
rect 1256 3594 1536 3636
rect 1256 3358 1278 3594
rect 1514 3358 1536 3594
rect 1256 3316 1536 3358
rect 360 2458 402 2694
rect 638 2458 680 2694
rect 360 1894 680 2458
rect 360 1658 402 1894
rect 638 1658 680 1894
rect 360 1616 680 1658
rect 2560 2694 2880 5558
rect 2560 2458 2602 2694
rect 2838 2458 2880 2694
rect 2560 1894 2880 2458
rect 2560 1658 2602 1894
rect 2838 1658 2880 1894
rect -300 998 -258 1234
rect -22 998 20 1234
rect -300 956 20 998
rect 2560 956 2880 1658
rect 4110 12602 4430 12644
rect 4110 12366 4152 12602
rect 4388 12366 4430 12602
rect 4110 10912 4430 12366
rect 4110 10848 4118 10912
rect 4182 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4430 10912
rect 4110 10444 4430 10848
rect 4110 10208 4152 10444
rect 4388 10208 4430 10444
rect 4110 9824 4430 10208
rect 4110 9760 4118 9824
rect 4182 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4430 9824
rect 4110 8736 4430 9760
rect 4110 8672 4118 8736
rect 4182 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4430 8736
rect 4110 7648 4430 8672
rect 4110 7584 4118 7648
rect 4182 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4430 7648
rect 4110 7344 4430 7584
rect 4110 7108 4152 7344
rect 4388 7108 4430 7344
rect 4110 6560 4430 7108
rect 4110 6496 4118 6560
rect 4182 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4430 6560
rect 4110 5472 4430 6496
rect 4110 5408 4118 5472
rect 4182 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4430 5472
rect 4110 4384 4430 5408
rect 4110 4320 4118 4384
rect 4182 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4430 4384
rect 4110 4244 4430 4320
rect 4110 4008 4152 4244
rect 4388 4008 4430 4244
rect 4110 3296 4430 4008
rect 4110 3232 4118 3296
rect 4182 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4430 3296
rect 4110 2208 4430 3232
rect 4110 2144 4118 2208
rect 4182 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4430 2208
rect 4110 1234 4430 2144
rect 4110 998 4152 1234
rect 4388 998 4430 1234
rect 4110 956 4430 998
rect 5660 11942 5980 12644
rect 5660 11706 5702 11942
rect 5938 11706 5980 11942
rect 5660 11456 5980 11706
rect 5660 11392 5668 11456
rect 5732 11392 5748 11456
rect 5812 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5980 11456
rect 5660 10368 5980 11392
rect 5660 10304 5668 10368
rect 5732 10304 5748 10368
rect 5812 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5980 10368
rect 5660 9280 5980 10304
rect 5660 9216 5668 9280
rect 5732 9216 5748 9280
rect 5812 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5980 9280
rect 5660 8894 5980 9216
rect 5660 8658 5702 8894
rect 5938 8658 5980 8894
rect 5660 8192 5980 8658
rect 5660 8128 5668 8192
rect 5732 8128 5748 8192
rect 5812 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5980 8192
rect 5660 7104 5980 8128
rect 5660 7040 5668 7104
rect 5732 7040 5748 7104
rect 5812 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5980 7104
rect 5660 6016 5980 7040
rect 5660 5952 5668 6016
rect 5732 5952 5748 6016
rect 5812 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5980 6016
rect 5660 5794 5980 5952
rect 5660 5558 5702 5794
rect 5938 5558 5980 5794
rect 5660 4928 5980 5558
rect 5660 4864 5668 4928
rect 5732 4864 5748 4928
rect 5812 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5980 4928
rect 5660 3840 5980 4864
rect 5660 3776 5668 3840
rect 5732 3776 5748 3840
rect 5812 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5980 3840
rect 5660 2752 5980 3776
rect 5660 2688 5668 2752
rect 5732 2694 5748 2752
rect 5812 2694 5828 2752
rect 5892 2694 5908 2752
rect 5972 2688 5980 2752
rect 5660 2458 5702 2688
rect 5938 2458 5980 2688
rect 5660 1894 5980 2458
rect 5660 1658 5702 1894
rect 5938 1658 5980 1894
rect 5660 956 5980 1658
rect 7210 12602 7530 12644
rect 7210 12366 7252 12602
rect 7488 12366 7530 12602
rect 7210 10912 7530 12366
rect 7210 10848 7218 10912
rect 7282 10848 7298 10912
rect 7362 10848 7378 10912
rect 7442 10848 7458 10912
rect 7522 10848 7530 10912
rect 7210 10444 7530 10848
rect 7210 10208 7252 10444
rect 7488 10208 7530 10444
rect 7210 9824 7530 10208
rect 7210 9760 7218 9824
rect 7282 9760 7298 9824
rect 7362 9760 7378 9824
rect 7442 9760 7458 9824
rect 7522 9760 7530 9824
rect 7210 8736 7530 9760
rect 7210 8672 7218 8736
rect 7282 8672 7298 8736
rect 7362 8672 7378 8736
rect 7442 8672 7458 8736
rect 7522 8672 7530 8736
rect 7210 7648 7530 8672
rect 7210 7584 7218 7648
rect 7282 7584 7298 7648
rect 7362 7584 7378 7648
rect 7442 7584 7458 7648
rect 7522 7584 7530 7648
rect 7210 7344 7530 7584
rect 7210 7108 7252 7344
rect 7488 7108 7530 7344
rect 7210 6560 7530 7108
rect 7210 6496 7218 6560
rect 7282 6496 7298 6560
rect 7362 6496 7378 6560
rect 7442 6496 7458 6560
rect 7522 6496 7530 6560
rect 7210 5472 7530 6496
rect 7210 5408 7218 5472
rect 7282 5408 7298 5472
rect 7362 5408 7378 5472
rect 7442 5408 7458 5472
rect 7522 5408 7530 5472
rect 7210 4384 7530 5408
rect 7210 4320 7218 4384
rect 7282 4320 7298 4384
rect 7362 4320 7378 4384
rect 7442 4320 7458 4384
rect 7522 4320 7530 4384
rect 7210 4244 7530 4320
rect 7210 4008 7252 4244
rect 7488 4008 7530 4244
rect 7210 3296 7530 4008
rect 7210 3232 7218 3296
rect 7282 3232 7298 3296
rect 7362 3232 7378 3296
rect 7442 3232 7458 3296
rect 7522 3232 7530 3296
rect 7210 2208 7530 3232
rect 7210 2144 7218 2208
rect 7282 2144 7298 2208
rect 7362 2144 7378 2208
rect 7442 2144 7458 2208
rect 7522 2144 7530 2208
rect 7210 1234 7530 2144
rect 7210 998 7252 1234
rect 7488 998 7530 1234
rect 7210 956 7530 998
rect 8760 11942 9080 12644
rect 10744 12602 11064 12644
rect 10744 12366 10786 12602
rect 11022 12366 11064 12602
rect 8760 11706 8802 11942
rect 9038 11706 9080 11942
rect 8760 11456 9080 11706
rect 8760 11392 8768 11456
rect 8832 11392 8848 11456
rect 8912 11392 8928 11456
rect 8992 11392 9008 11456
rect 9072 11392 9080 11456
rect 8760 10368 9080 11392
rect 8760 10304 8768 10368
rect 8832 10304 8848 10368
rect 8912 10304 8928 10368
rect 8992 10304 9008 10368
rect 9072 10304 9080 10368
rect 8760 9280 9080 10304
rect 8760 9216 8768 9280
rect 8832 9216 8848 9280
rect 8912 9216 8928 9280
rect 8992 9216 9008 9280
rect 9072 9216 9080 9280
rect 8760 8894 9080 9216
rect 8760 8658 8802 8894
rect 9038 8658 9080 8894
rect 8760 8192 9080 8658
rect 8760 8128 8768 8192
rect 8832 8128 8848 8192
rect 8912 8128 8928 8192
rect 8992 8128 9008 8192
rect 9072 8128 9080 8192
rect 8760 7104 9080 8128
rect 8760 7040 8768 7104
rect 8832 7040 8848 7104
rect 8912 7040 8928 7104
rect 8992 7040 9008 7104
rect 9072 7040 9080 7104
rect 8760 6016 9080 7040
rect 8760 5952 8768 6016
rect 8832 5952 8848 6016
rect 8912 5952 8928 6016
rect 8992 5952 9008 6016
rect 9072 5952 9080 6016
rect 8760 5794 9080 5952
rect 8760 5558 8802 5794
rect 9038 5558 9080 5794
rect 8760 4928 9080 5558
rect 8760 4864 8768 4928
rect 8832 4864 8848 4928
rect 8912 4864 8928 4928
rect 8992 4864 9008 4928
rect 9072 4864 9080 4928
rect 8760 3840 9080 4864
rect 8760 3776 8768 3840
rect 8832 3776 8848 3840
rect 8912 3776 8928 3840
rect 8992 3776 9008 3840
rect 9072 3776 9080 3840
rect 8760 2752 9080 3776
rect 8760 2688 8768 2752
rect 8832 2694 8848 2752
rect 8912 2694 8928 2752
rect 8992 2694 9008 2752
rect 9072 2688 9080 2752
rect 8760 2458 8802 2688
rect 9038 2458 9080 2688
rect 8760 1894 9080 2458
rect 8760 1658 8802 1894
rect 9038 1658 9080 1894
rect 8760 956 9080 1658
rect 10084 11942 10404 11984
rect 10084 11706 10126 11942
rect 10362 11706 10404 11942
rect 10084 8894 10404 11706
rect 10084 8658 10126 8894
rect 10362 8658 10404 8894
rect 10084 5794 10404 8658
rect 10084 5558 10126 5794
rect 10362 5558 10404 5794
rect 10084 2694 10404 5558
rect 10084 2458 10126 2694
rect 10362 2458 10404 2694
rect 10084 1894 10404 2458
rect 10084 1658 10126 1894
rect 10362 1658 10404 1894
rect 10084 1616 10404 1658
rect 10744 10444 11064 12366
rect 10744 10208 10786 10444
rect 11022 10208 11064 10444
rect 10744 7344 11064 10208
rect 10744 7108 10786 7344
rect 11022 7108 11064 7344
rect 10744 4244 11064 7108
rect 10744 4008 10786 4244
rect 11022 4008 11064 4244
rect 10744 1234 11064 4008
rect 10744 998 10786 1234
rect 11022 998 11064 1234
rect 10744 956 11064 998
rect 11404 9794 11724 13026
rect 11404 9558 11446 9794
rect 11682 9558 11724 9794
rect 11404 6694 11724 9558
rect 11404 6458 11446 6694
rect 11682 6458 11724 6694
rect 11404 3594 11724 6458
rect 11404 3358 11446 3594
rect 11682 3358 11724 3594
rect -960 338 -918 574
rect -682 338 -640 574
rect -960 296 -640 338
rect 11404 574 11724 3358
rect 11404 338 11446 574
rect 11682 338 11724 574
rect 11404 296 11724 338
rect 12064 8244 12384 13686
rect 12064 8008 12106 8244
rect 12342 8008 12384 8244
rect 12064 5144 12384 8008
rect 12064 4908 12106 5144
rect 12342 4908 12384 5144
rect -1620 -322 -1578 -86
rect -1342 -322 -1300 -86
rect -1620 -364 -1300 -322
rect 12064 -86 12384 4908
rect 12064 -322 12106 -86
rect 12342 -322 12384 -86
rect 12064 -364 12384 -322
<< via4 >>
rect -1578 13686 -1342 13922
rect 12106 13686 12342 13922
rect -1578 8008 -1342 8244
rect -1578 4908 -1342 5144
rect -918 13026 -682 13262
rect 11446 13026 11682 13262
rect -918 9558 -682 9794
rect -918 6458 -682 6694
rect -918 3358 -682 3594
rect -258 12366 -22 12602
rect -258 10208 -22 10444
rect -258 7108 -22 7344
rect -258 4008 -22 4244
rect 402 11706 638 11942
rect 402 8658 638 8894
rect 402 5558 638 5794
rect 2602 11706 2838 11942
rect 2602 8658 2838 8894
rect 2602 5558 2838 5794
rect 2018 4908 2254 5144
rect 1278 3358 1514 3594
rect 402 2458 638 2694
rect 402 1658 638 1894
rect 2602 2458 2838 2694
rect 2602 1658 2838 1894
rect -258 998 -22 1234
rect 4152 12366 4388 12602
rect 4152 10208 4388 10444
rect 4152 7108 4388 7344
rect 4152 4008 4388 4244
rect 4152 998 4388 1234
rect 5702 11706 5938 11942
rect 5702 8658 5938 8894
rect 5702 5558 5938 5794
rect 5702 2688 5732 2694
rect 5732 2688 5748 2694
rect 5748 2688 5812 2694
rect 5812 2688 5828 2694
rect 5828 2688 5892 2694
rect 5892 2688 5908 2694
rect 5908 2688 5938 2694
rect 5702 2458 5938 2688
rect 5702 1658 5938 1894
rect 7252 12366 7488 12602
rect 7252 10208 7488 10444
rect 7252 7108 7488 7344
rect 7252 4008 7488 4244
rect 7252 998 7488 1234
rect 10786 12366 11022 12602
rect 8802 11706 9038 11942
rect 8802 8658 9038 8894
rect 8802 5558 9038 5794
rect 8802 2688 8832 2694
rect 8832 2688 8848 2694
rect 8848 2688 8912 2694
rect 8912 2688 8928 2694
rect 8928 2688 8992 2694
rect 8992 2688 9008 2694
rect 9008 2688 9038 2694
rect 8802 2458 9038 2688
rect 8802 1658 9038 1894
rect 10126 11706 10362 11942
rect 10126 8658 10362 8894
rect 10126 5558 10362 5794
rect 10126 2458 10362 2694
rect 10126 1658 10362 1894
rect 10786 10208 11022 10444
rect 10786 7108 11022 7344
rect 10786 4008 11022 4244
rect 10786 998 11022 1234
rect 11446 9558 11682 9794
rect 11446 6458 11682 6694
rect 11446 3358 11682 3594
rect -918 338 -682 574
rect 11446 338 11682 574
rect 12106 8008 12342 8244
rect 12106 4908 12342 5144
rect -1578 -322 -1342 -86
rect 12106 -322 12342 -86
<< metal5 >>
rect -1620 13922 12384 13964
rect -1620 13686 -1578 13922
rect -1342 13686 12106 13922
rect 12342 13686 12384 13922
rect -1620 13644 12384 13686
rect -960 13262 11724 13304
rect -960 13026 -918 13262
rect -682 13026 11446 13262
rect 11682 13026 11724 13262
rect -960 12984 11724 13026
rect -300 12602 11064 12644
rect -300 12366 -258 12602
rect -22 12366 4152 12602
rect 4388 12366 7252 12602
rect 7488 12366 10786 12602
rect 11022 12366 11064 12602
rect -300 12324 11064 12366
rect 360 11942 10404 11984
rect 360 11706 402 11942
rect 638 11706 2602 11942
rect 2838 11706 5702 11942
rect 5938 11706 8802 11942
rect 9038 11706 10126 11942
rect 10362 11706 10404 11942
rect 360 11664 10404 11706
rect -300 10444 11064 10486
rect -300 10208 -258 10444
rect -22 10208 4152 10444
rect 4388 10208 7252 10444
rect 7488 10208 10786 10444
rect 11022 10208 11064 10444
rect -300 10166 11064 10208
rect -1620 9794 12384 9836
rect -1620 9558 -918 9794
rect -682 9558 11446 9794
rect 11682 9558 12384 9794
rect -1620 9516 12384 9558
rect -300 8894 11064 8936
rect -300 8658 402 8894
rect 638 8658 2602 8894
rect 2838 8658 5702 8894
rect 5938 8658 8802 8894
rect 9038 8658 10126 8894
rect 10362 8658 11064 8894
rect -300 8616 11064 8658
rect -1620 8244 12384 8286
rect -1620 8008 -1578 8244
rect -1342 8008 12106 8244
rect 12342 8008 12384 8244
rect -1620 7966 12384 8008
rect -300 7344 11064 7386
rect -300 7108 -258 7344
rect -22 7108 4152 7344
rect 4388 7108 7252 7344
rect 7488 7108 10786 7344
rect 11022 7108 11064 7344
rect -300 7066 11064 7108
rect -1620 6694 12384 6736
rect -1620 6458 -918 6694
rect -682 6458 11446 6694
rect 11682 6458 12384 6694
rect -1620 6416 12384 6458
rect -300 5794 11064 5836
rect -300 5558 402 5794
rect 638 5558 2602 5794
rect 2838 5558 5702 5794
rect 5938 5558 8802 5794
rect 9038 5558 10126 5794
rect 10362 5558 11064 5794
rect -300 5516 11064 5558
rect -1620 5144 12384 5186
rect -1620 4908 -1578 5144
rect -1342 4908 2018 5144
rect 2254 4908 12106 5144
rect 12342 4908 12384 5144
rect -1620 4866 12384 4908
rect -300 4244 11064 4286
rect -300 4008 -258 4244
rect -22 4008 4152 4244
rect 4388 4008 7252 4244
rect 7488 4008 10786 4244
rect 11022 4008 11064 4244
rect -300 3966 11064 4008
rect -1620 3594 12384 3636
rect -1620 3358 -918 3594
rect -682 3358 1278 3594
rect 1514 3358 11446 3594
rect 11682 3358 12384 3594
rect -1620 3316 12384 3358
rect -300 2694 11064 2736
rect -300 2458 402 2694
rect 638 2458 2602 2694
rect 2838 2458 5702 2694
rect 5938 2458 8802 2694
rect 9038 2458 10126 2694
rect 10362 2458 11064 2694
rect -300 2416 11064 2458
rect 360 1894 10404 1936
rect 360 1658 402 1894
rect 638 1658 2602 1894
rect 2838 1658 5702 1894
rect 5938 1658 8802 1894
rect 9038 1658 10126 1894
rect 10362 1658 10404 1894
rect 360 1616 10404 1658
rect -300 1234 11064 1276
rect -300 998 -258 1234
rect -22 998 4152 1234
rect 4388 998 7252 1234
rect 7488 998 10786 1234
rect 11022 998 11064 1234
rect -300 956 11064 998
rect -960 574 11724 616
rect -960 338 -918 574
rect -682 338 11446 574
rect 11682 338 11724 574
rect -960 296 11724 338
rect -1620 -86 12384 -44
rect -1620 -322 -1578 -86
rect -1342 -322 12106 -86
rect 12342 -322 12384 -86
rect -1620 -364 12384 -322
use sky130_fd_sc_hd__clkbuf_1  _150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635271187
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635271187
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1635271187
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635271187
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635271187
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635271187
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1635271187
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform -1 0 3496 0 1 4352
box -38 -48 222 592
use gpio_logic_high  gpio_logic_high
timestamp 1636035201
transform 1 0 1196 0 1 2680
box -38 -48 1418 2768
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1635271187
transform 1 0 3864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1635271187
transform 1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46
timestamp 1635271187
transform 1 0 5152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50
timestamp 1635271187
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52
timestamp 1635271187
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1635271187
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 4692 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__dfbbn_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3496 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__dfrtp_1  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3404 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfbbn_1  _203_
timestamp 1635271187
transform 1 0 5704 0 1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1635271187
transform 1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1635271187
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1635271187
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _204_
timestamp 1635271187
transform 1 0 4416 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1635271187
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1635271187
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1635271187
transform 1 0 3772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_34
timestamp 1635271187
transform 1 0 4048 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3496 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 1635271187
transform 1 0 3772 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _102_
timestamp 1635271187
transform 1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1635271187
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _217_
timestamp 1635271187
transform 1 0 3956 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfbbn_1  _209_
timestamp 1635271187
transform 1 0 5796 0 -1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1635271187
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_32
timestamp 1635271187
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59
timestamp 1635271187
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1635271187
transform 1 0 6440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1635271187
transform 1 0 6440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _139_
timestamp 1635271187
transform 1 0 5888 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 1635271187
transform 1 0 5888 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1635271187
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1635271187
transform 1 0 6716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _145_
timestamp 1635271187
transform 1 0 6808 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _147_
timestamp 1635271187
transform 1 0 6992 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1635271187
transform 1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1635271187
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1635271187
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _179_
timestamp 1635271187
transform 1 0 7636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1635271187
transform 1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1635271187
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1635271187
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1635271187
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1635271187
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1635271187
transform 1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1635271187
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1635271187
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1635271187
transform 1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _108_
timestamp 1635271187
transform 1 0 8280 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1635271187
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_64
timestamp 1635271187
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfbbn_1  _208_
timestamp 1635271187
transform 1 0 7176 0 1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1635271187
transform 1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1635271187
transform 1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1635271187
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1635271187
transform 1 0 6532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1635271187
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1635271187
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8648 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1635271187
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1635271187
transform 1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1635271187
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_83
timestamp 1635271187
transform 1 0 8556 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635271187
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635271187
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1635271187
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92
timestamp 1635271187
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _116_
timestamp 1635271187
transform 1 0 8924 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _114_
timestamp 1635271187
transform 1 0 8372 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635271187
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_92
timestamp 1635271187
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__and2_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8832 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1635271187
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635271187
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635271187
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 1635271187
transform 1 0 9108 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _110_
timestamp 1635271187
transform 1 0 8648 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635271187
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _214_
timestamp 1635271187
transform 1 0 3312 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635271187
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635271187
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635271187
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _213_
timestamp 1635271187
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635271187
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1635271187
transform -1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1635271187
transform 1 0 1196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635271187
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635271187
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635271187
transform 1 0 1288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635271187
transform 1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635271187
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_16
timestamp 1635271187
transform 1 0 2392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635271187
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1635271187
transform -1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_20
timestamp 1635271187
transform 1 0 2760 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1635271187
transform -1 0 3312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1635271187
transform -1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1635271187
transform 1 0 1196 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635271187
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635271187
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635271187
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635271187
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635271187
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1635271187
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1635271187
transform 1 0 3036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635271187
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1635271187
transform -1 0 3404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1635271187
transform 1 0 5704 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp 1635271187
transform 1 0 5152 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1635271187
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _210_
timestamp 1635271187
transform 1 0 4140 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__or2_1  _171_
timestamp 1635271187
transform 1 0 3680 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__dfbbn_1  _199_
timestamp 1635271187
transform 1 0 3588 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1635271187
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _218_
timestamp 1635271187
transform 1 0 4048 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1635271187
transform -1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1635271187
transform -1 0 3864 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1635271187
transform -1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _222_
timestamp 1635271187
transform 1 0 4692 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1635271187
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_39
timestamp 1635271187
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1635271187
transform 1 0 3404 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1635271187
transform -1 0 4140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1635271187
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1635271187
transform -1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1635271187
transform -1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1635271187
transform -1 0 4324 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfbbn_1  _205_
timestamp 1635271187
transform 1 0 6624 0 1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1635271187
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_61
timestamp 1635271187
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1635271187
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _126_
timestamp 1635271187
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6532 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1635271187
transform 1 0 8188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_77
timestamp 1635271187
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6164 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _132_
timestamp 1635271187
transform 1 0 8004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1635271187
transform 1 0 6072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1635271187
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _206_
timestamp 1635271187
transform 1 0 6164 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1635271187
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1635271187
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1635271187
transform 1 0 6532 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__or2_1  _128_
timestamp 1635271187
transform 1 0 9016 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635271187
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1635271187
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8648 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635271187
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp 1635271187
transform 1 0 9476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1635271187
transform 1 0 8740 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1635271187
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1635271187
transform 1 0 8556 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635271187
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _183_
timestamp 1635271187
transform 1 0 8740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1635271187
transform 1 0 8556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1635271187
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635271187
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _120_
timestamp 1635271187
transform 1 0 8740 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1635271187
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1635271187
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1635271187
transform 1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635271187
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635271187
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _219_
timestamp 1635271187
transform 1 0 2576 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1635271187
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1635271187
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635271187
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1635271187
transform 1 0 1196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1635271187
transform 1 0 1932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1635271187
transform -1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635271187
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1635271187
transform 1 0 1196 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635271187
transform 1 0 1472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1635271187
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1635271187
transform -1 0 2392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_12
timestamp 1635271187
transform 1 0 2024 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1635271187
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635271187
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1635271187
transform 1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1635271187
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1635271187
transform 1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1635271187
transform 1 0 3128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635271187
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1196 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_22
timestamp 1635271187
transform 1 0 2944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_11
timestamp 1635271187
transform 1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1635271187
transform 1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1635271187
transform 1 0 1196 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635271187
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635271187
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 1196 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1635271187
transform 1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1635271187
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1635271187
transform 1 0 1564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1635271187
transform 1 0 1656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635271187
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635271187
transform 1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1635271187
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1635271187
transform -1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1635271187
transform 1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1635271187
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1635271187
transform 1 0 2944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1635271187
transform 1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _212_
timestamp 1635271187
transform 1 0 2392 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__or2b_1  _163_
timestamp 1635271187
transform 1 0 5336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_
timestamp 1635271187
transform 1 0 4416 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1635271187
transform 1 0 5428 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1635271187
transform 1 0 3588 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1635271187
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _200_
timestamp 1635271187
transform 1 0 3680 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1635271187
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _211_
timestamp 1635271187
transform 1 0 4232 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfbbn_1  _201_
timestamp 1635271187
transform 1 0 4600 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1635271187
transform 1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1635271187
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1635271187
transform 1 0 4232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1635271187
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_39
timestamp 1635271187
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1635271187
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 6440 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dfbbn_1  _207_
timestamp 1635271187
transform 1 0 7176 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1635271187
transform 1 0 6164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1635271187
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1635271187
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1635271187
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _186_
timestamp 1635271187
transform 1 0 8188 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_12_75
timestamp 1635271187
transform 1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_69
timestamp 1635271187
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1635271187
transform -1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_12  input17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 8096 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__einvp_2  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635271187
transform 1 0 7452 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1635271187
transform 1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _165_
timestamp 1635271187
transform 1 0 6716 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _157_
timestamp 1635271187
transform 1 0 6164 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1635271187
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfbbn_1  _198_
timestamp 1635271187
transform 1 0 6256 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__or2_1  _177_
timestamp 1635271187
transform 1 0 8004 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _175_
timestamp 1635271187
transform 1 0 7452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _159_
timestamp 1635271187
transform 1 0 6992 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1635271187
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1635271187
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635271187
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1635271187
transform 1 0 9200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1635271187
transform 1 0 8740 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1635271187
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635271187
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp 1635271187
transform 1 0 8740 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1635271187
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1635271187
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635271187
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635271187
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp 1635271187
transform 1 0 8648 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635271187
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_93
timestamp 1635271187
transform 1 0 9476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635271187
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635271187
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1635271187
transform 1 0 1564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1635271187
transform 1 0 1196 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1635271187
transform -1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1635271187
transform 1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_15
timestamp 1635271187
transform 1 0 2300 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1635271187
transform 1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1635271187
transform -1 0 2300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp 1635271187
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1635271187
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1635271187
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1635271187
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1635271187
transform 1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1635271187
transform 1 0 5336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1635271187
transform 1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1635271187
transform 1 0 4968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1635271187
transform 1 0 4600 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1635271187
transform 1 0 4232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1635271187
transform 1 0 3864 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_77
timestamp 1635271187
transform 1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1635271187
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1635271187
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1635271187
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1635271187
transform 1 0 6900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1635271187
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1635271187
transform 1 0 8280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1635271187
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1635271187
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635271187
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1635271187
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _191_
timestamp 1635271187
transform 1 0 8832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1635271187
transform 1 0 9200 0 1 10880
box -38 -48 406 592
<< labels >>
rlabel metal3 s 14000 1640 34000 1760 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal3 s 14000 4904 34000 5024 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal3 s 14000 5312 34000 5432 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal3 s 14000 5584 34000 5704 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal3 s 14000 2320 34000 2440 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal3 s 14000 2728 34000 2848 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal3 s 14000 3000 34000 3120 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal3 s 14000 3272 34000 3392 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal3 s 14000 3680 34000 3800 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal3 s 14000 3952 34000 4072 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal3 s 14000 4360 34000 4480 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal3 s 14000 4632 34000 4752 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 688 34000 808 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1096 34000 1216 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 1368 34000 1488 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 416 34000 536 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 5992 34000 6112 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 6264 34000 6384 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 7216 34000 7336 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 7896 34000 8016 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 8576 34000 8696 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 8848 34000 8968 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 9256 34000 9376 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 9528 34000 9648 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 10208 34000 10328 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 10480 34000 10600 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 10888 34000 11008 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 11160 34000 11280 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 11432 34000 11552 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 12112 34000 12232 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 12520 34000 12640 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 12792 34000 12912 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 13472 34000 13592 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 13744 34000 13864 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 360 1616 10404 1936 6 vccd
port 42 nsew power input
rlabel metal5 s -300 2416 11064 2736 6 vccd
port 42 nsew power input
rlabel metal5 s -300 5516 11064 5836 6 vccd
port 42 nsew power input
rlabel metal5 s -300 8616 11064 8936 6 vccd
port 42 nsew power input
rlabel metal5 s 360 11664 10404 11984 6 vccd
port 42 nsew power input
rlabel metal4 s 360 1616 680 11984 6 vccd
port 42 nsew power input
rlabel metal4 s 10084 1616 10404 11984 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 956 2880 12644 6 vccd
port 42 nsew power input
rlabel metal4 s 5660 956 5980 12644 6 vccd
port 42 nsew power input
rlabel metal4 s 8760 956 9080 12644 6 vccd
port 42 nsew power input
rlabel metal5 s -960 296 11724 616 6 vccd1
port 43 nsew power input
rlabel metal5 s -1620 3316 12384 3636 6 vccd1
port 43 nsew power input
rlabel metal5 s -1620 6416 12384 6736 6 vccd1
port 43 nsew power input
rlabel metal5 s -1620 9516 12384 9836 6 vccd1
port 43 nsew power input
rlabel metal5 s -960 12984 11724 13304 6 vccd1
port 43 nsew power input
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 43 nsew power input
rlabel metal4 s 11404 296 11724 13304 6 vccd1
port 43 nsew power input
rlabel metal5 s -300 956 11064 1276 6 vssd
port 44 nsew ground input
rlabel metal5 s -300 3966 11064 4286 6 vssd
port 44 nsew ground input
rlabel metal5 s -300 7066 11064 7386 6 vssd
port 44 nsew ground input
rlabel metal5 s -300 10166 11064 10486 6 vssd
port 44 nsew ground input
rlabel metal5 s -300 12324 11064 12644 6 vssd
port 44 nsew ground input
rlabel metal4 s -300 956 20 12644 4 vssd
port 44 nsew ground input
rlabel metal4 s 4110 956 4430 12644 6 vssd
port 44 nsew ground input
rlabel metal4 s 7210 956 7530 12644 6 vssd
port 44 nsew ground input
rlabel metal4 s 10744 956 11064 12644 6 vssd
port 44 nsew ground input
rlabel metal5 s -1620 -364 12384 -44 8 vssd1
port 45 nsew ground input
rlabel metal5 s -1620 4866 12384 5186 6 vssd1
port 45 nsew ground input
rlabel metal5 s -1620 7966 12384 8286 6 vssd1
port 45 nsew ground input
rlabel metal5 s -1620 13644 12384 13964 6 vssd1
port 45 nsew ground input
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 45 nsew ground input
rlabel metal4 s 12064 -364 12384 13964 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 144 34000 264 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 14000
<< end >>
