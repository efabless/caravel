module caravan_signal_routing();
endmodule