VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan_core
  CLASS BLOCK ;
  FOREIGN caravan_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END caravan_core
END LIBRARY

