* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv vccd vssd vdda1 vssa1 vdda2 vssa2 mprj2_vdd_logic1 mprj_vdd_logic1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufbuf_8 abstract view
.subckt sky130_fd_sc_hd__bufbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1_uq1 vccd2_uq0 vdda1_uq0 vdda2_uq0 vssd vssd2_uq0
+ vssa1_uq0 vssa2_uq0 vssd1_uq1
XANTENNA_wire1828_A wire1828/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_4541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1902 wire1902/A vssd vssd vccd vccd wire1902/X sky130_fd_sc_hd__buf_6
XFILLER_41_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1913 wire1913/A vssd vssd vccd vccd _257_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1924 wire1924/A vssd vssd vccd vccd _335_/A sky130_fd_sc_hd__buf_6
Xwire1935 wire1935/A vssd vssd vccd vccd _332_/A sky130_fd_sc_hd__buf_6
Xwire1946 wire1947/X vssd vssd vccd vccd _191_/A sky130_fd_sc_hd__buf_6
XTAP_3202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1957 wire1957/A vssd vssd vccd vccd wire1957/X sky130_fd_sc_hd__buf_6
XTAP_3213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1968 wire1969/X vssd vssd vccd vccd _176_/A sky130_fd_sc_hd__buf_6
XFILLER_41_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1979 wire1979/A vssd vssd vccd vccd _169_/A sky130_fd_sc_hd__buf_6
XTAP_3235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input127_A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2044_A wire2044/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_501_ _501_/A _501_/B vssd vssd vccd vccd _501_/X sky130_fd_sc_hd__and2_4
XTAP_2512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 wire1985/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_224 _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_432_ _560_/A _432_/B _432_/C vssd vssd vccd vccd _432_/X sky130_fd_sc_hd__and3b_4
XANTENNA_257 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_363_ _363_/A _363_/B vssd vssd vccd vccd _363_/X sky130_fd_sc_hd__and2_2
XTAP_1888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input92_A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_294_ _294_/A _294_/B vssd vssd vccd vccd _294_/X sky130_fd_sc_hd__and2_2
XFILLER_48_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] max_cap1456/X vssd vssd vccd vccd _122_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output513_A wire1292/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1311_A wire1312/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output882_A wire1066/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1409_A _319_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] _188_/X vssd vssd vccd vccd _008_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1778_A wire1779/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__304__A _304_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1945_A wire1945/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput467 wire1212/X vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__buf_8
Xoutput478 _482_/X vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__buf_8
XFILLER_42_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput489 wire1205/X vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__buf_8
XFILLER_47_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1209 _475_/X vssd vssd vccd vccd wire1209/X sky130_fd_sc_hd__buf_6
XFILLER_25_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__490__A_N _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4242 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__214__A _214_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2161_A wire2162/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input244_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2259_A wire2260/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1710 wire1710/A vssd vssd vccd vccd _559_/A sky130_fd_sc_hd__buf_6
XFILLER_25_2980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1721 wire1721/A vssd vssd vccd vccd _527_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1732 wire1732/A vssd vssd vccd vccd _612_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1743 wire1743/A vssd vssd vccd vccd _191_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1754 wire1754/A vssd vssd vccd vccd _440_/C sky130_fd_sc_hd__buf_6
XFILLER_19_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input411_A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1765 wire1765/A vssd vssd vccd vccd wire1765/X sky130_fd_sc_hd__buf_6
XTAP_3021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1776 wire1777/X vssd vssd vccd vccd _383_/B sky130_fd_sc_hd__buf_6
XFILLER_20_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1787 wire1787/A vssd vssd vccd vccd wire1787/X sky130_fd_sc_hd__buf_6
XTAP_3043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1798 wire1799/X vssd vssd vccd vccd _374_/B sky130_fd_sc_hd__buf_6
XTAP_3054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ _543_/A _415_/B _415_/C vssd vssd vccd vccd _415_/X sky130_fd_sc_hd__and3b_4
XTAP_2397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_346_ _346_/A _346_/B vssd vssd vccd vccd _346_/X sky130_fd_sc_hd__and2_4
XFILLER_30_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_277_ _277_/A _277_/B vssd vssd vccd vccd _277_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output463_A wire1294/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1094_A wire1095/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output728_A _605_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1359_A wire1360/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1526_A wire1527/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1895_A wire1896/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire979_A wire980/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__034__A _034_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1006 wire1007/X vssd vssd vccd vccd wire1006/X sky130_fd_sc_hd__buf_6
XFILLER_25_2276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1017 wire1018/X vssd vssd vccd vccd wire1017/X sky130_fd_sc_hd__buf_6
Xwire1028 wire1029/X vssd vssd vccd vccd wire1028/X sky130_fd_sc_hd__buf_6
XFILLER_38_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1039 wire1040/X vssd vssd vccd vccd wire1039/X sky130_fd_sc_hd__buf_6
XFILLER_28_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__209__A _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_200_ _200_/A _200_/B vssd vssd vccd vccd _200_/X sky130_fd_sc_hd__and2_2
XFILLER_23_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2007_A wire2008/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_131_ _131_/A vssd vssd vccd vccd _131_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input194_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_062_ _062_/A vssd vssd vccd vccd _062_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__386__A_N _514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input361_A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input459_A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input55_A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__598__B _598_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2230 wire2231/X vssd vssd vccd vccd _473_/B sky130_fd_sc_hd__buf_6
Xwire2241 wire2241/A vssd vssd vccd vccd wire2241/X sky130_fd_sc_hd__buf_6
XFILLER_38_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2252 wire2253/X vssd vssd vccd vccd _457_/B sky130_fd_sc_hd__buf_6
Xwire2263 wire2264/X vssd vssd vccd vccd wire2263/X sky130_fd_sc_hd__buf_6
XFILLER_21_4098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2274 wire2274/A vssd vssd vccd vccd wire2274/X sky130_fd_sc_hd__buf_6
XFILLER_47_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1540 wire1541/X vssd vssd vccd vccd _349_/B sky130_fd_sc_hd__buf_6
Xwire2285 wire2285/A vssd vssd vccd vccd _441_/B sky130_fd_sc_hd__buf_6
Xwire1551 wire1552/X vssd vssd vccd vccd wire1551/X sky130_fd_sc_hd__buf_6
XFILLER_21_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2296 wire2296/A vssd vssd vccd vccd _432_/B sky130_fd_sc_hd__buf_6
Xwire1562 wire1563/X vssd vssd vccd vccd wire1562/X sky130_fd_sc_hd__buf_6
Xwire1573 wire1574/X vssd vssd vccd vccd wire1573/X sky130_fd_sc_hd__buf_6
XFILLER_19_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1584 wire1585/X vssd vssd vccd vccd wire1584/X sky130_fd_sc_hd__buf_6
Xwire1595 wire1596/X vssd vssd vccd vccd wire1595/X sky130_fd_sc_hd__buf_6
XFILLER_1_2768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__119__A _119_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output580_A wire1223/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1107_A wire1108/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_329_ _329_/A _329_/B vssd vssd vccd vccd _329_/X sky130_fd_sc_hd__and2_4
XFILLER_30_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output845_A _596_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1476_A _246_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] wire1467/X vssd vssd vccd vccd wire1125/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_45_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1643_A wire1644/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__301__B _301_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1810_A wire1811/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__029__A _029_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__211__B _211_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2124_A wire2125/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input207_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_114_ _114_/A vssd vssd vccd vccd _114_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_045_ _045_/A vssd vssd vccd vccd _045_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2060 wire2061/X vssd vssd vccd vccd _599_/B sky130_fd_sc_hd__buf_6
Xwire2071 wire2072/X vssd vssd vccd vccd wire2071/X sky130_fd_sc_hd__buf_6
XFILLER_21_3172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2082 wire2082/A vssd vssd vccd vccd _590_/B sky130_fd_sc_hd__buf_6
XFILLER_38_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1057_A wire1058/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2093 wire2094/X vssd vssd vccd vccd wire2093/X sky130_fd_sc_hd__buf_6
XFILLER_1_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__401__A_N _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1370 wire1371/X vssd vssd vccd vccd wire1370/X sky130_fd_sc_hd__buf_6
XFILLER_19_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1381 _343_/X vssd vssd vccd vccd wire1381/X sky130_fd_sc_hd__buf_6
XFILLER_53_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1392 _339_/X vssd vssd vccd vccd wire1392/X sky130_fd_sc_hd__buf_6
XFILLER_1_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1224_A _458_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output795_A wire1156/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3820 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] load_slew1458/X vssd vssd vccd vccd _134_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_15_2264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1593_A wire1594/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1760_A wire1760/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__312__A _312_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1338 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__206__B _206_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2074_A wire2075/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input157_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput301 la_oenb_mprj[21] vssd vssd vccd vccd _518_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__424__A_N _552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput312 la_oenb_mprj[31] vssd vssd vccd vccd _400_/A_N sky130_fd_sc_hd__buf_6
XFILLER_7_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput323 la_oenb_mprj[41] vssd vssd vccd vccd _538_/A sky130_fd_sc_hd__buf_4
XFILLER_44_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput334 la_oenb_mprj[51] vssd vssd vccd vccd wire1712/A sky130_fd_sc_hd__buf_6
XFILLER_2_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput345 la_oenb_mprj[61] vssd vssd vccd vccd _558_/A sky130_fd_sc_hd__clkbuf_4
Xinput356 la_oenb_mprj[71] vssd vssd vccd vccd wire1701/A sky130_fd_sc_hd__buf_6
Xinput367 la_oenb_mprj[81] vssd vssd vccd vccd wire1691/A sky130_fd_sc_hd__buf_6
XANTENNA_input324_A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput378 la_oenb_mprj[91] vssd vssd vccd vccd _588_/A sky130_fd_sc_hd__buf_4
XFILLER_40_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput389 mprj_adr_o_core[10] vssd vssd vccd vccd wire1674/A sky130_fd_sc_hd__buf_6
XFILLER_2_3597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input18_A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_594_ _594_/A _594_/B vssd vssd vccd vccd _594_/X sky130_fd_sc_hd__and2_4
XFILLER_21_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1774 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_5 _554_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput808 _562_/X vssd vssd vccd vccd la_oenb_core[65] sky130_fd_sc_hd__buf_8
Xoutput819 _572_/X vssd vssd vccd vccd la_oenb_core[75] sky130_fd_sc_hd__buf_8
X_028_ _028_/A vssd vssd vccd vccd _028_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output543_A wire1231/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__132__A _132_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1174_A _523_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output710_A _075_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1341_A wire1342/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1439_A _302_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] _218_/X vssd vssd vccd vccd _038_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1606_A wire1606/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3926 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__307__A _307_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1975_A wire1975/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire961_A wire962/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__447__A_N _447_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__217__A _217_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input274_A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2191_A wire2192/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2289_A wire2290/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input441_A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput120 la_data_out_mprj[8] vssd vssd vccd vccd _377_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput131 la_data_out_mprj[9] vssd vssd vccd vccd _378_/C sky130_fd_sc_hd__clkbuf_4
Xinput142 la_iena_mprj[109] vssd vssd vccd vccd _272_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput153 la_iena_mprj[119] vssd vssd vccd vccd _282_/B sky130_fd_sc_hd__buf_4
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput164 la_iena_mprj[13] vssd vssd vccd vccd _176_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 la_iena_mprj[23] vssd vssd vccd vccd _186_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 la_iena_mprj[33] vssd vssd vccd vccd _196_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput197 la_iena_mprj[43] vssd vssd vccd vccd _206_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_577_ _577_/A _577_/B vssd vssd vccd vccd _577_/X sky130_fd_sc_hd__and2_4
XFILLER_32_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output493_A wire1201/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output660_A _030_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output758_A wire1199/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1291_A _372_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1389_A wire1390/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput605 _095_/Y vssd vssd vccd vccd la_data_in_mprj[112] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[43\]_B _206_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput616 _105_/Y vssd vssd vccd vccd la_data_in_mprj[122] sky130_fd_sc_hd__buf_8
XFILLER_29_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput627 _000_/Y vssd vssd vccd vccd la_data_in_mprj[17] sky130_fd_sc_hd__buf_8
XFILLER_29_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput638 _010_/Y vssd vssd vccd vccd la_data_in_mprj[27] sky130_fd_sc_hd__buf_8
XANTENNA_output925_A wire1337/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput649 _020_/Y vssd vssd vccd vccd la_data_in_mprj[37] sky130_fd_sc_hd__buf_8
XFILLER_29_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1556_A wire1557/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1723_A wire1724/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__037__A _037_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[34\]_B _197_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1903 wire1904/X vssd vssd vccd vccd _263_/A sky130_fd_sc_hd__buf_6
XANTENNA__500__A _500_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1914 wire1914/A vssd vssd vccd vccd _256_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1925 wire1925/A vssd vssd vccd vccd _242_/A sky130_fd_sc_hd__buf_4
XFILLER_41_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1936 wire1936/A vssd vssd vccd vccd _209_/A sky130_fd_sc_hd__buf_4
Xwire1947 wire1947/A vssd vssd vccd vccd wire1947/X sky130_fd_sc_hd__buf_6
XTAP_3203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1958 wire1958/A vssd vssd vccd vccd _329_/A sky130_fd_sc_hd__buf_6
XFILLER_19_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1969 wire1969/A vssd vssd vccd vccd wire1969/X sky130_fd_sc_hd__buf_6
XTAP_3225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_500_ _500_/A _500_/B vssd vssd vccd vccd _500_/X sky130_fd_sc_hd__and2_4
XFILLER_22_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_225 _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_431_ _559_/A _431_/B _431_/C vssd vssd vccd vccd _431_/X sky130_fd_sc_hd__and3b_2
XTAP_2557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ _362_/A _362_/B vssd vssd vccd vccd _362_/X sky130_fd_sc_hd__and2_2
XANTENNA_wire2204_A wire2205/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_293_ _293_/A _293_/B vssd vssd vccd vccd _293_/X sky130_fd_sc_hd__and2_1
XANTENNA_input391_A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input85_A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4102 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output506_A wire1271/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1137_A wire1137/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_2421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1304_A wire1305/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output875_A _310_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] _181_/X vssd vssd vccd vccd _001_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1673_A wire1674/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[100\]_B _263_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__304__B _304_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1840_A wire1840/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput468 wire1211/X vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__buf_8
XFILLER_9_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput479 _483_/X vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__buf_8
XFILLER_42_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__320__A _320_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4254 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__214__B _214_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__230__A _230_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1700 wire1700/A vssd vssd vccd vccd _569_/A sky130_fd_sc_hd__buf_8
Xwire1711 wire1711/A vssd vssd vccd vccd _555_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1722 wire1722/A vssd vssd vccd vccd _526_/A sky130_fd_sc_hd__buf_6
XANTENNA_input237_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1733 wire1733/A vssd vssd vccd vccd _611_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1744 input18/X vssd vssd vccd vccd _481_/C sky130_fd_sc_hd__buf_4
XFILLER_46_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1755 wire1755/A vssd vssd vccd vccd _304_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1766 wire1767/X vssd vssd vccd vccd _387_/B sky130_fd_sc_hd__buf_6
XTAP_3011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1777 wire1777/A vssd vssd vccd vccd wire1777/X sky130_fd_sc_hd__buf_6
XTAP_3033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1788 wire1789/X vssd vssd vccd vccd _377_/B sky130_fd_sc_hd__buf_6
XFILLER_41_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1799 wire1799/A vssd vssd vccd vccd wire1799/X sky130_fd_sc_hd__buf_6
XTAP_3055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input404_A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _542_/A _414_/B _414_/C vssd vssd vccd vccd _414_/X sky130_fd_sc_hd__and3b_4
XFILLER_19_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _345_/A _345_/B vssd vssd vccd vccd _345_/X sky130_fd_sc_hd__and2_4
XFILLER_50_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_276_ _276_/A _276_/B vssd vssd vccd vccd _276_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1087_A wire1088/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1254_A _408_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_2355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1421_A _314_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1519_A wire1519/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1790_A wire1791/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1888_A wire1888/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__315__A _315_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__050__A _050_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1007 wire1008/X vssd vssd vccd vccd wire1007/X sky130_fd_sc_hd__buf_6
Xwire1018 wire1019/X vssd vssd vccd vccd wire1018/X sky130_fd_sc_hd__buf_6
XFILLER_0_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1029 wire1030/X vssd vssd vccd vccd wire1029/X sky130_fd_sc_hd__buf_6
XFILLER_38_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__209__B _209_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_582 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_130_ _130_/A vssd vssd vccd vccd _130_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_7_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1082 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__225__A _225_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_061_ _061_/A vssd vssd vccd vccd _061_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input187_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input354_A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2271_A wire2272/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input48_A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2220 wire2221/X vssd vssd vccd vccd _478_/B sky130_fd_sc_hd__buf_6
Xwire2231 wire2231/A vssd vssd vccd vccd wire2231/X sky130_fd_sc_hd__buf_6
XFILLER_43_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2242 wire2243/X vssd vssd vccd vccd _466_/B sky130_fd_sc_hd__buf_6
XFILLER_21_4088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2253 wire2254/X vssd vssd vccd vccd wire2253/X sky130_fd_sc_hd__buf_6
XFILLER_21_3354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2264 wire2264/A vssd vssd vccd vccd wire2264/X sky130_fd_sc_hd__buf_6
XFILLER_5_2861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1530 wire1531/X vssd vssd vccd vccd _354_/B sky130_fd_sc_hd__buf_6
Xwire2275 wire2276/X vssd vssd vccd vccd _449_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1541 wire1541/A vssd vssd vccd vccd wire1541/X sky130_fd_sc_hd__buf_6
Xwire2286 wire2286/A vssd vssd vccd vccd _440_/B sky130_fd_sc_hd__buf_6
XFILLER_47_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1552 wire1552/A vssd vssd vccd vccd wire1552/X sky130_fd_sc_hd__buf_6
Xwire2297 wire2297/A vssd vssd vccd vccd _307_/A sky130_fd_sc_hd__buf_6
XFILLER_46_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1563 wire1563/A vssd vssd vccd vccd wire1563/X sky130_fd_sc_hd__buf_6
XFILLER_4_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1574 wire1575/X vssd vssd vccd vccd wire1574/X sky130_fd_sc_hd__buf_6
XFILLER_38_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1585 wire1586/X vssd vssd vccd vccd wire1585/X sky130_fd_sc_hd__buf_6
XFILLER_19_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1596 wire1596/A vssd vssd vccd vccd wire1596/X sky130_fd_sc_hd__buf_6
XFILLER_46_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1002_A wire1003/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_328_ _328_/A _328_/B vssd vssd vccd vccd _328_/X sky130_fd_sc_hd__and2_4
XANTENNA_output573_A _453_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_259_ _259_/A _259_/B vssd vssd vccd vccd _259_/X sky130_fd_sc_hd__and2_2
XFILLER_7_940 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output740_A _616_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output838_A _589_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1371_A wire1372/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1469_A _253_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__480__A_N _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] wire1474/X vssd vssd vccd vccd wire1130/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1636_A wire1636/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1803_A wire1803/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3902 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__045__A _045_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3018 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1723 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input102_A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2117_A wire2117/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_113_ _113_/A vssd vssd vccd vccd _113_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_044_ _044_/A vssd vssd vccd vccd _044_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2050 wire2051/X vssd vssd vccd vccd _604_/B sky130_fd_sc_hd__buf_6
XFILLER_43_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2061 wire2061/A vssd vssd vccd vccd wire2061/X sky130_fd_sc_hd__buf_6
Xwire2072 wire2073/X vssd vssd vccd vccd wire2072/X sky130_fd_sc_hd__buf_6
Xwire2083 wire2083/A vssd vssd vccd vccd _589_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2094 wire2094/A vssd vssd vccd vccd wire2094/X sky130_fd_sc_hd__buf_6
XFILLER_47_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1360 _350_/X vssd vssd vccd vccd wire1360/X sky130_fd_sc_hd__buf_6
Xwire1371 wire1372/X vssd vssd vccd vccd wire1371/X sky130_fd_sc_hd__buf_6
Xwire1382 wire1383/X vssd vssd vccd vccd wire1382/X sky130_fd_sc_hd__buf_6
Xwire1393 wire1394/X vssd vssd vccd vccd wire1393/X sky130_fd_sc_hd__buf_6
XFILLER_19_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output690_A _057_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output788_A _544_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output955_A wire1453/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] split4/A vssd vssd vccd vccd _127_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_28_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__312__B _312_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[1\]_A mprj_dat_i_user[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] _274_/X vssd vssd vccd vccd _094_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_1_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__376__A_N _504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__503__A _503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput302 la_oenb_mprj[22] vssd vssd vccd vccd _519_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput313 la_oenb_mprj[32] vssd vssd vccd vccd wire1719/A sky130_fd_sc_hd__buf_6
XFILLER_2_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput324 la_oenb_mprj[42] vssd vssd vccd vccd _539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput335 la_oenb_mprj[52] vssd vssd vccd vccd _549_/A sky130_fd_sc_hd__buf_4
XANTENNA_wire2067_A wire2067/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput346 la_oenb_mprj[62] vssd vssd vccd vccd wire1710/A sky130_fd_sc_hd__buf_6
XFILLER_22_3471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput357 la_oenb_mprj[72] vssd vssd vccd vccd wire1700/A sky130_fd_sc_hd__buf_6
Xinput368 la_oenb_mprj[82] vssd vssd vccd vccd wire1690/A sky130_fd_sc_hd__buf_6
XFILLER_5_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput379 la_oenb_mprj[92] vssd vssd vccd vccd _589_/A sky130_fd_sc_hd__buf_6
XFILLER_25_1170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input317_A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2234_A wire2235/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_593_ _593_/A _593_/B vssd vssd vccd vccd _593_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_6 _554_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput809 _563_/X vssd vssd vccd vccd la_oenb_core[66] sky130_fd_sc_hd__buf_8
X_027_ _027_/A vssd vssd vccd vccd _027_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_46_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output536_A wire1243/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1167_A wire1168/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__399__A_N _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1334_A wire1335/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1190 _507_/X vssd vssd vccd vccd wire1190/X sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] _211_/X vssd vssd vccd vccd _031_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_34_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3943 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1501_A wire1502/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__307__B _307_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1870_A wire1871/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1968_A wire1969/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__323__A _323_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_850 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1147 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__233__A _233_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2184_A wire2184/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input267_A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2832 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input434_A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput110 la_data_out_mprj[80] vssd vssd vccd vccd wire1753/A sky130_fd_sc_hd__buf_6
XFILLER_4_2926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput121 la_data_out_mprj[90] vssd vssd vccd vccd _459_/C sky130_fd_sc_hd__clkbuf_4
Xinput132 la_iena_mprj[0] vssd vssd vccd vccd _625_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input30_A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput143 la_iena_mprj[10] vssd vssd vccd vccd _173_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput154 la_iena_mprj[11] vssd vssd vccd vccd _174_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput165 la_iena_mprj[14] vssd vssd vccd vccd _177_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput176 la_iena_mprj[24] vssd vssd vccd vccd _187_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput187 la_iena_mprj[34] vssd vssd vccd vccd _197_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput198 la_iena_mprj[44] vssd vssd vccd vccd _207_/B sky130_fd_sc_hd__buf_4
XTAP_4675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_576_ _576_/A _576_/B vssd vssd vccd vccd _576_/X sky130_fd_sc_hd__and2_4
XFILLER_16_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output486_A _489_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output653_A _023_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput606 _096_/Y vssd vssd vccd vccd la_data_in_mprj[113] sky130_fd_sc_hd__buf_8
XANTENNA__143__A _143_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2710 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput617 _106_/Y vssd vssd vccd vccd la_data_in_mprj[123] sky130_fd_sc_hd__buf_8
XANTENNA_wire1284_A _379_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput628 _001_/Y vssd vssd vccd vccd la_data_in_mprj[18] sky130_fd_sc_hd__buf_8
Xoutput639 _011_/Y vssd vssd vccd vccd la_data_in_mprj[28] sky130_fd_sc_hd__buf_8
XFILLER_29_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output820_A _573_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output918_A wire1355/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1451_A _299_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1549_A wire1550/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1716_A _406_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_964 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__318__A _318_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__414__A_N _542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__053__A _053_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1904 wire1904/A vssd vssd vccd vccd wire1904/X sky130_fd_sc_hd__buf_6
XANTENNA__500__B _500_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1915 wire1915/A vssd vssd vccd vccd _255_/A sky130_fd_sc_hd__buf_6
Xwire1926 wire1926/A vssd vssd vccd vccd _238_/A sky130_fd_sc_hd__buf_6
XTAP_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1937 wire1937/A vssd vssd vccd vccd _208_/A sky130_fd_sc_hd__buf_6
Xwire1948 wire1948/A vssd vssd vccd vccd _190_/A sky130_fd_sc_hd__buf_6
XTAP_3204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1959 wire1960/X vssd vssd vccd vccd _182_/A sky130_fd_sc_hd__buf_6
XTAP_3215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 wire2022/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_226 _559_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ _558_/A _430_/B _430_/C vssd vssd vccd vccd _430_/X sky130_fd_sc_hd__and3b_4
XFILLER_19_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_248 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_614 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4071 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_259 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__228__A _228_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_361_ _361_/A _361_/B vssd vssd vccd vccd _361_/X sky130_fd_sc_hd__and2_1
XTAP_1868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_292_ _292_/A _292_/B vssd vssd vccd vccd _292_/X sky130_fd_sc_hd__and2_1
XFILLER_35_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input384_A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input78_A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__B _410_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1032_A wire1033/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__437__A_N _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__138__A _138_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_559_ _559_/A _559_/B vssd vssd vccd vccd _559_/X sky130_fd_sc_hd__and2_4
XFILLER_31_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output868_A _333_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1499_A wire1500/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1666_A wire1667/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput469 wire1210/X vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__buf_8
XFILLER_47_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__601__A _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1833_A wire1833/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__320__B _320_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__048__A _048_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1139 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__511__A _511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__230__B _230_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1701 wire1701/A vssd vssd vccd vccd _568_/A sky130_fd_sc_hd__buf_6
XFILLER_43_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1712 wire1712/A vssd vssd vccd vccd _548_/A sky130_fd_sc_hd__buf_6
Xwire1723 wire1724/X vssd vssd vccd vccd _295_/A_N sky130_fd_sc_hd__buf_6
Xwire1734 wire1734/A vssd vssd vccd vccd _610_/A sky130_fd_sc_hd__buf_6
Xwire1745 wire1745/A vssd vssd vccd vccd _457_/C sky130_fd_sc_hd__buf_6
XFILLER_19_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input132_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1756 wire1757/X vssd vssd vccd vccd _394_/B sky130_fd_sc_hd__buf_6
XFILLER_46_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2147_A wire2148/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4122 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1767 wire1767/A vssd vssd vccd vccd wire1767/X sky130_fd_sc_hd__buf_6
XTAP_3012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1778 wire1779/X vssd vssd vccd vccd _382_/B sky130_fd_sc_hd__buf_6
XTAP_3034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1789 wire1789/A vssd vssd vccd vccd wire1789/X sky130_fd_sc_hd__buf_6
XTAP_3045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1075 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_413_ _541_/A _413_/B _413_/C vssd vssd vccd vccd _413_/X sky130_fd_sc_hd__and3b_4
XTAP_2377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _344_/A _344_/B vssd vssd vccd vccd _344_/X sky130_fd_sc_hd__and2_2
XFILLER_53_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_275_ _275_/A _275_/B vssd vssd vccd vccd _275_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output616_A _105_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1247_A _415_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1414_A wire1415/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] _193_/X vssd vssd vccd vccd _013_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_33_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_904 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1783_A wire1783/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__315__B _315_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1950_A wire1950/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__331__A _331_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1008 wire1009/X vssd vssd vccd vccd wire1008/X sky130_fd_sc_hd__buf_6
XFILLER_5_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1019 wire1020/X vssd vssd vccd vccd wire1019/X sky130_fd_sc_hd__buf_6
XFILLER_9_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_A mprj_ack_i_user vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__506__A _506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__225__B _225_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_060_ _060_/A vssd vssd vccd vccd _060_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2097_A wire2098/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__241__A _241_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2264_A wire2264/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input347_A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2210 wire2211/X vssd vssd vccd vccd wire2210/X sky130_fd_sc_hd__buf_6
XFILLER_21_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2221 wire2221/A vssd vssd vccd vccd wire2221/X sky130_fd_sc_hd__buf_6
XFILLER_25_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2232 wire2233/X vssd vssd vccd vccd _472_/B sky130_fd_sc_hd__buf_6
XFILLER_48_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2243 wire2243/A vssd vssd vccd vccd wire2243/X sky130_fd_sc_hd__buf_6
XFILLER_5_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2254 wire2254/A vssd vssd vccd vccd wire2254/X sky130_fd_sc_hd__buf_6
XFILLER_43_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1520 wire1520/A vssd vssd vccd vccd _361_/B sky130_fd_sc_hd__buf_6
Xwire2265 wire2266/X vssd vssd vccd vccd _453_/B sky130_fd_sc_hd__buf_6
Xwire1531 wire1531/A vssd vssd vccd vccd wire1531/X sky130_fd_sc_hd__buf_6
Xwire2276 wire2276/A vssd vssd vccd vccd wire2276/X sky130_fd_sc_hd__buf_6
XFILLER_48_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1542 wire1543/X vssd vssd vccd vccd _348_/B sky130_fd_sc_hd__buf_6
Xwire2287 wire2287/A vssd vssd vccd vccd _439_/B sky130_fd_sc_hd__buf_6
Xwire1553 wire1554/X vssd vssd vccd vccd _314_/B sky130_fd_sc_hd__buf_6
Xwire2298 wire2298/A vssd vssd vccd vccd _306_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1564 wire1565/X vssd vssd vccd vccd _311_/B sky130_fd_sc_hd__buf_6
XFILLER_0_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1575 wire1576/X vssd vssd vccd vccd wire1575/X sky130_fd_sc_hd__buf_6
Xwire1586 wire1586/A vssd vssd vccd vccd wire1586/X sky130_fd_sc_hd__buf_6
XFILLER_21_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1597 wire1598/X vssd vssd vccd vccd _334_/B sky130_fd_sc_hd__buf_8
XFILLER_47_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2594 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_327_ _327_/A _327_/B vssd vssd vccd vccd _327_/X sky130_fd_sc_hd__and2_4
XFILLER_15_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_258_ _258_/A _258_/B vssd vssd vccd vccd _258_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3760 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output566_A _447_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_189_ _189_/A _189_/B vssd vssd vccd vccd _189_/X sky130_fd_sc_hd__and2_1
XFILLER_6_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1197_A _500_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output733_A _609_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1364_A wire1365/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output900_A wire982/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] wire1481/X vssd vssd vccd vccd wire1137/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_22_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1629_A wire1629/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1998_A wire1999/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire984_A wire985/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__A _326_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__061__A _061_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1735 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2012_A wire2012/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__236__A _236_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input297_A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_112_ _112_/A vssd vssd vccd vccd _112_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_043_ _043_/A vssd vssd vccd vccd _043_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_4243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input60_A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__402__C _402_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2040 wire2041/X vssd vssd vccd vccd _608_/B sky130_fd_sc_hd__buf_6
Xwire2051 wire2051/A vssd vssd vccd vccd wire2051/X sky130_fd_sc_hd__buf_6
XFILLER_43_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2062 wire2063/X vssd vssd vccd vccd _598_/B sky130_fd_sc_hd__buf_6
Xwire2073 wire2073/A vssd vssd vccd vccd wire2073/X sky130_fd_sc_hd__buf_6
XFILLER_5_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2084 wire2085/X vssd vssd vccd vccd _588_/B sky130_fd_sc_hd__buf_6
Xwire1350 wire1351/X vssd vssd vccd vccd wire1350/X sky130_fd_sc_hd__buf_6
XFILLER_21_3196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2095 wire2096/X vssd vssd vccd vccd _582_/B sky130_fd_sc_hd__buf_6
Xwire1361 wire1362/X vssd vssd vccd vccd wire1361/X sky130_fd_sc_hd__buf_6
XFILLER_1_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1372 _346_/X vssd vssd vccd vccd wire1372/X sky130_fd_sc_hd__buf_6
Xwire1383 wire1384/X vssd vssd vccd vccd wire1383/X sky130_fd_sc_hd__buf_6
XFILLER_1_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1394 _338_/X vssd vssd vccd vccd wire1394/X sky130_fd_sc_hd__buf_6
XFILLER_47_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1112_A wire1113/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output683_A _051_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output850_A wire1414/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output948_A wire1426/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1481_A _241_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1579_A wire1580/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1746_A wire1746/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[1\]_B max_cap1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1913_A wire1913/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] _267_/X vssd vssd vccd vccd _087_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__056__A _056_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1610 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__503__B _503_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput303 la_oenb_mprj[23] vssd vssd vccd vccd _520_/A sky130_fd_sc_hd__buf_4
XFILLER_44_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput314 la_oenb_mprj[33] vssd vssd vccd vccd _530_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput325 la_oenb_mprj[43] vssd vssd vccd vccd _540_/A sky130_fd_sc_hd__buf_6
Xinput336 la_oenb_mprj[53] vssd vssd vccd vccd _550_/A sky130_fd_sc_hd__buf_4
XFILLER_40_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput347 la_oenb_mprj[63] vssd vssd vccd vccd wire1709/A sky130_fd_sc_hd__buf_6
Xinput358 la_oenb_mprj[73] vssd vssd vccd vccd wire1699/A sky130_fd_sc_hd__buf_6
XFILLER_22_3483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput369 la_oenb_mprj[83] vssd vssd vccd vccd wire1689/A sky130_fd_sc_hd__buf_6
XFILLER_2_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xload_slew1457 load_slew1458/X vssd vssd vccd vccd split4/A sky130_fd_sc_hd__buf_8
XFILLER_1_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input212_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_592_ _592_/A _592_/B vssd vssd vccd vccd _592_/X sky130_fd_sc_hd__and2_4
XFILLER_43_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2227_A wire2227/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__A_N _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_7 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_026_ _026_/A vssd vssd vccd vccd _026_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__413__B _413_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2502 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output529_A wire1249/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1062_A wire1063/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1180 _517_/X vssd vssd vccd vccd wire1180/X sky130_fd_sc_hd__buf_6
XFILLER_1_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1191 _506_/X vssd vssd vccd vccd wire1191/X sky130_fd_sc_hd__buf_6
XFILLER_1_2364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1327_A wire1328/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output898_A wire992/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__604__A _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__323__B _323_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__493__A_N _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1830 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__514__A _514_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__233__B _233_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input162_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2177_A wire2178/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput100 la_data_out_mprj[71] vssd vssd vccd vccd wire1754/A sky130_fd_sc_hd__buf_6
XFILLER_2_4042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput111 la_data_out_mprj[81] vssd vssd vccd vccd wire1752/A sky130_fd_sc_hd__buf_6
XFILLER_44_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput122 la_data_out_mprj[91] vssd vssd vccd vccd _460_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput133 la_iena_mprj[100] vssd vssd vccd vccd _263_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput144 la_iena_mprj[110] vssd vssd vccd vccd _273_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input427_A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 la_iena_mprj[120] vssd vssd vccd vccd _283_/B sky130_fd_sc_hd__buf_4
XFILLER_24_2888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 la_iena_mprj[15] vssd vssd vccd vccd _178_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input23_A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput177 la_iena_mprj[25] vssd vssd vccd vccd _188_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput188 la_iena_mprj[35] vssd vssd vccd vccd _198_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput199 la_iena_mprj[45] vssd vssd vccd vccd _208_/B sky130_fd_sc_hd__buf_4
XFILLER_17_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_575_ _575_/A _575_/B vssd vssd vccd vccd _575_/X sky130_fd_sc_hd__and2_4
XFILLER_44_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__408__B _408_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output479_A _483_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_29_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput607 _097_/Y vssd vssd vccd vccd la_data_in_mprj[114] sky130_fd_sc_hd__buf_8
XFILLER_9_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput618 _107_/Y vssd vssd vccd vccd la_data_in_mprj[124] sky130_fd_sc_hd__buf_8
Xoutput629 _002_/Y vssd vssd vccd vccd la_data_in_mprj[19] sky130_fd_sc_hd__buf_8
XFILLER_25_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output646_A _017_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_009_ _009_/A vssd vssd vccd vccd _009_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1277_A _386_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output813_A wire1194/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1444_A _301_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] _223_/X vssd vssd vccd vccd _043_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1611_A wire1611/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__318__B _318_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1980_A wire1981/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__334__A _334_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1905 wire1906/X vssd vssd vccd vccd _262_/A sky130_fd_sc_hd__buf_6
XTAP_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1916 wire1916/A vssd vssd vccd vccd _254_/A sky130_fd_sc_hd__buf_6
XFILLER_3_4395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1927 wire1927/A vssd vssd vccd vccd _234_/A sky130_fd_sc_hd__buf_4
XFILLER_41_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1938 wire1938/A vssd vssd vccd vccd _207_/A sky130_fd_sc_hd__buf_6
XTAP_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1949 wire1949/A vssd vssd vccd vccd _189_/A sky130_fd_sc_hd__buf_6
XTAP_3205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_216 wire2063/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_227 wire2164/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__509__A _509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__228__B _228_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_360_ _360_/A _360_/B vssd vssd vccd vccd _360_/X sky130_fd_sc_hd__and2_1
XTAP_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_291_ _291_/A _291_/B vssd vssd vccd vccd _291_/X sky130_fd_sc_hd__and2_1
XFILLER_52_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__A _244_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__389__A_N _517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2294_A wire2294/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input377_A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_751 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_558_ _558_/A _558_/B vssd vssd vccd vccd _558_/X sky130_fd_sc_hd__and2_2
XANTENNA_wire1025_A _133_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output596_A _087_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_489_ _617_/A _489_/B _489_/C vssd vssd vccd vccd _489_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output763_A wire1176/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1394_A _338_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output930_A wire1319/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1561_A wire1562/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1659_A wire1660/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__601__B _601_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1826_A wire1826/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__329__A _329_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__064__A _064_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput960 _295_/X vssd vssd vccd vccd user_reset sky130_fd_sc_hd__buf_8
XANTENNA__511__B _511_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1702 wire1702/A vssd vssd vccd vccd _567_/A sky130_fd_sc_hd__buf_6
Xwire1713 wire1713/A vssd vssd vccd vccd _544_/A sky130_fd_sc_hd__buf_6
XFILLER_25_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1724 wire1725/X vssd vssd vccd vccd wire1724/X sky130_fd_sc_hd__buf_6
Xwire1735 wire1735/A vssd vssd vccd vccd _609_/A sky130_fd_sc_hd__buf_6
XFILLER_19_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1746 wire1746/A vssd vssd vccd vccd _456_/C sky130_fd_sc_hd__buf_6
XTAP_3002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1757 wire1757/A vssd vssd vccd vccd wire1757/X sky130_fd_sc_hd__buf_6
Xwire1768 wire1769/X vssd vssd vccd vccd _386_/B sky130_fd_sc_hd__buf_6
XTAP_3013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1779 wire1779/A vssd vssd vccd vccd wire1779/X sky130_fd_sc_hd__buf_6
XTAP_3035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2042_A wire2043/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__239__A _239_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ _540_/A _412_/B _412_/C vssd vssd vccd vccd _412_/X sky130_fd_sc_hd__and3b_4
XTAP_2367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_343_ _343_/A _343_/B vssd vssd vccd vccd _343_/X sky130_fd_sc_hd__and2_2
XTAP_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input90_A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_274_ _274_/A _274_/B vssd vssd vccd vccd _274_/X sky130_fd_sc_hd__and2_4
XFILLER_52_2391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__405__C _405_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] split4/X vssd vssd vccd vccd _120_/A sky130_fd_sc_hd__nand2_4
XFILLER_48_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4092 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__421__B _421_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__404__A_N _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output511_A wire1265/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output609_A _099_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1407_A _320_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output880_A wire1452/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] _186_/X vssd vssd vccd vccd _006_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3728 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1776_A wire1777/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__612__A _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1943_A wire1943/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__331__B _331_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1009 wire1010/X vssd vssd vccd vccd wire1009/X sky130_fd_sc_hd__buf_6
XFILLER_5_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__059__A _059_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_B max_cap1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__506__B _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__522__A _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__427__A_N _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2200 wire2201/X vssd vssd vccd vccd _485_/B sky130_fd_sc_hd__buf_6
Xoutput790 wire1162/X vssd vssd vccd vccd la_oenb_core[49] sky130_fd_sc_hd__buf_8
XFILLER_5_3542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2211 wire2211/A vssd vssd vccd vccd wire2211/X sky130_fd_sc_hd__buf_6
Xwire2222 wire2223/X vssd vssd vccd vccd _477_/B sky130_fd_sc_hd__buf_6
XANTENNA_input242_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2233 wire2233/A vssd vssd vccd vccd wire2233/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2257_A wire2257/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2244 wire2244/A vssd vssd vccd vccd _465_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1510 wire1510/A vssd vssd vccd vccd wire1510/X sky130_fd_sc_hd__buf_6
Xwire2255 wire2256/X vssd vssd vccd vccd _456_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1521 wire1521/A vssd vssd vccd vccd _360_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2266 wire2267/X vssd vssd vccd vccd wire2266/X sky130_fd_sc_hd__buf_6
XFILLER_4_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1532 wire1533/X vssd vssd vccd vccd _353_/B sky130_fd_sc_hd__buf_6
Xwire2277 wire2277/A vssd vssd vccd vccd _448_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1543 wire1543/A vssd vssd vccd vccd wire1543/X sky130_fd_sc_hd__buf_6
Xwire2288 wire2288/A vssd vssd vccd vccd _438_/B sky130_fd_sc_hd__buf_6
XFILLER_48_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1554 wire1555/X vssd vssd vccd vccd wire1554/X sky130_fd_sc_hd__buf_6
Xwire2299 wire2299/A vssd vssd vccd vccd _305_/A sky130_fd_sc_hd__buf_6
Xwire1565 wire1566/X vssd vssd vccd vccd wire1565/X sky130_fd_sc_hd__buf_6
XFILLER_4_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1576 wire1576/A vssd vssd vccd vccd wire1576/X sky130_fd_sc_hd__buf_6
XFILLER_38_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1587 wire1588/X vssd vssd vccd vccd _335_/B sky130_fd_sc_hd__buf_8
XFILLER_46_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1598 wire1599/X vssd vssd vccd vccd wire1598/X sky130_fd_sc_hd__buf_6
XFILLER_21_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_326_ _326_/A _326_/B vssd vssd vccd vccd _326_/X sky130_fd_sc_hd__and2_4
XFILLER_9_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__416__B _416_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_257_ _257_/A _257_/B vssd vssd vccd vccd _257_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_188_ _188_/A _188_/B vssd vssd vccd vccd _188_/X sky130_fd_sc_hd__and2_1
XFILLER_26_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output559_A _440_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1092_A wire1093/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output726_A _603_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1357_A _351_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1524_A wire1524/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__A _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1893_A wire1894/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__B _326_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire977_A _143_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[91\]_B wire1468/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__342__A _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__517__A _517_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__236__B _236_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2005_A wire2006/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_111_ _111_/A vssd vssd vccd vccd _111_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_input192_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[82\]_B wire1477/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_042_ _042_/A vssd vssd vccd vccd _042_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__252__A _252_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input457_A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input53_A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2030 wire2031/X vssd vssd vccd vccd wire2030/X sky130_fd_sc_hd__buf_6
Xwire2041 wire2041/A vssd vssd vccd vccd wire2041/X sky130_fd_sc_hd__buf_6
Xwire2052 wire2053/X vssd vssd vccd vccd _603_/B sky130_fd_sc_hd__buf_6
XFILLER_38_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2063 wire2063/A vssd vssd vccd vccd wire2063/X sky130_fd_sc_hd__buf_6
Xwire2074 wire2075/X vssd vssd vccd vccd _594_/B sky130_fd_sc_hd__buf_6
Xwire1340 wire1341/X vssd vssd vccd vccd wire1340/X sky130_fd_sc_hd__buf_6
XFILLER_1_2502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2085 wire2085/A vssd vssd vccd vccd wire2085/X sky130_fd_sc_hd__buf_6
Xwire2096 wire2096/A vssd vssd vccd vccd wire2096/X sky130_fd_sc_hd__buf_6
Xwire1351 _353_/X vssd vssd vccd vccd wire1351/X sky130_fd_sc_hd__buf_6
Xwire1362 wire1363/X vssd vssd vccd vccd wire1362/X sky130_fd_sc_hd__buf_6
XFILLER_19_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1373 wire1374/X vssd vssd vccd vccd wire1373/X sky130_fd_sc_hd__buf_6
XFILLER_47_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1384 _342_/X vssd vssd vccd vccd wire1384/X sky130_fd_sc_hd__buf_6
Xwire1395 wire1396/X vssd vssd vccd vccd wire1395/X sky130_fd_sc_hd__buf_6
XFILLER_46_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_309_ _309_/A _309_/B vssd vssd vccd vccd _309_/X sky130_fd_sc_hd__and2_4
XFILLER_12_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[73\]_B _236_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output843_A _594_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__162__A _162_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1474_A _248_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] wire1469/X vssd vssd vccd vccd _073_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_28_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1641_A wire1642/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1739_A input22/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__337__A _337_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2610 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__072__A _072_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput304 la_oenb_mprj[24] vssd vssd vccd vccd _521_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_2081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput315 la_oenb_mprj[34] vssd vssd vccd vccd _531_/A sky130_fd_sc_hd__buf_4
XFILLER_22_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput326 la_oenb_mprj[44] vssd vssd vccd vccd _541_/A sky130_fd_sc_hd__buf_4
XFILLER_6_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput337 la_oenb_mprj[54] vssd vssd vccd vccd _551_/A sky130_fd_sc_hd__buf_8
XFILLER_29_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput348 la_oenb_mprj[64] vssd vssd vccd vccd wire1708/A sky130_fd_sc_hd__buf_6
XFILLER_40_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput359 la_oenb_mprj[74] vssd vssd vccd vccd wire1698/A sky130_fd_sc_hd__buf_6
XFILLER_5_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xload_slew1458 split5/A vssd vssd vccd vccd load_slew1458/X sky130_fd_sc_hd__buf_8
X_591_ _591_/A _591_/B vssd vssd vccd vccd _591_/X sky130_fd_sc_hd__and2_4
XFILLER_35_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2122_A wire2122/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input205_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__247__A _247_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[55\]_B _218_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_025_ _025_/A vssd vssd vccd vccd _025_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_8 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__413__C _413_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3226 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2514 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1055_A _127_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1170 _535_/X vssd vssd vccd vccd wire1170/X sky130_fd_sc_hd__buf_6
Xwire1181 _516_/X vssd vssd vccd vccd wire1181/X sky130_fd_sc_hd__buf_6
XFILLER_47_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1192 _505_/X vssd vssd vccd vccd wire1192/X sky130_fd_sc_hd__buf_6
XFILLER_1_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__295__A_N _295_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1222_A _460_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output793_A _548_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_370 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1591_A wire1591/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1689_A wire1689/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__604__B _604_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1856_A wire1857/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__620__A _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__067__A _067_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__514__B _514_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_B _284_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__A _530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input155_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2072_A wire2073/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput101 la_data_out_mprj[72] vssd vssd vccd vccd _441_/C sky130_fd_sc_hd__buf_4
XFILLER_7_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput112 la_data_out_mprj[82] vssd vssd vccd vccd wire1751/A sky130_fd_sc_hd__buf_6
XFILLER_7_1328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput123 la_data_out_mprj[92] vssd vssd vccd vccd _461_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput134 la_iena_mprj[101] vssd vssd vccd vccd _264_/B sky130_fd_sc_hd__buf_4
XTAP_4611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 la_iena_mprj[111] vssd vssd vccd vccd _274_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput156 la_iena_mprj[121] vssd vssd vccd vccd _284_/B sky130_fd_sc_hd__buf_4
XTAP_4633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input322_A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput167 la_iena_mprj[16] vssd vssd vccd vccd _179_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput178 la_iena_mprj[26] vssd vssd vccd vccd _189_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 la_iena_mprj[36] vssd vssd vccd vccd _199_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_574_ _574_/A _574_/B vssd vssd vccd vccd _574_/X sky130_fd_sc_hd__and2_4
XANTENNA_user_wb_dat_gates\[30\]_A mprj_dat_i_user[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2930 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[112\]_B _275_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__424__B _424_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput608 _098_/Y vssd vssd vccd vccd la_data_in_mprj[115] sky130_fd_sc_hd__buf_8
Xoutput619 _108_/Y vssd vssd vccd vccd la_data_in_mprj[125] sky130_fd_sc_hd__buf_8
X_008_ _008_/A vssd vssd vccd vccd _008_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output541_A wire1234/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output639_A _011_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1172_A _530_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output806_A _560_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1437_A wire1438/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] _216_/X vssd vssd vccd vccd _036_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1604_A wire1605/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[21\]_A mprj_dat_i_user[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3027 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__615__A _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[103\]_B _266_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__334__B _334_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__350__A _350_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__460__A_N _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input8_A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1906 wire1906/A vssd vssd vccd vccd wire1906/X sky130_fd_sc_hd__buf_6
XTAP_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1917 wire1917/A vssd vssd vccd vccd _253_/A sky130_fd_sc_hd__buf_4
XFILLER_6_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1928 wire1928/A vssd vssd vccd vccd _233_/A sky130_fd_sc_hd__buf_6
XTAP_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1939 wire1939/A vssd vssd vccd vccd _331_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 wire2073/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__509__B _509_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_239 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_A mprj_dat_i_user[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_290_ _290_/A _290_/B vssd vssd vccd vccd _290_/X sky130_fd_sc_hd__and2_2
XFILLER_22_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__525__A _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input272_A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2287_A wire2287/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__260__A _260_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2758 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__419__B _419_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_763 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_557_ _557_/A _557_/B vssd vssd vccd vccd _557_/X sky130_fd_sc_hd__and2_4
XFILLER_31_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1018_A wire1019/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_488_ _616_/A _488_/B _488_/C vssd vssd vccd vccd _488_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output491_A wire1203/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output589_A wire1216/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output756_A wire1182/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1387_A _341_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__483__A_N _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output923_A wire1340/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__170__A _170_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1554_A wire1555/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__329__B _329_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__345__A _345_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__080__A _080_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput950 wire1445/X vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__buf_8
XFILLER_25_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1703 wire1703/A vssd vssd vccd vccd _566_/A sky130_fd_sc_hd__buf_6
XFILLER_43_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1725 input3/X vssd vssd vccd vccd wire1725/X sky130_fd_sc_hd__buf_6
Xwire1736 wire1736/A vssd vssd vccd vccd _597_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1747 wire1747/A vssd vssd vccd vccd _455_/C sky130_fd_sc_hd__buf_6
XFILLER_24_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1758 wire1758/A vssd vssd vccd vccd _393_/B sky130_fd_sc_hd__buf_6
XFILLER_41_1551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1769 wire1769/A vssd vssd vccd vccd wire1769/X sky130_fd_sc_hd__buf_6
XTAP_3014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__239__B _239_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2035_A wire2036/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ _539_/A _411_/B _411_/C vssd vssd vccd vccd _411_/X sky130_fd_sc_hd__and3b_4
XTAP_2368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_342_ _342_/A _342_/B vssd vssd vccd vccd _342_/X sky130_fd_sc_hd__and2_2
XANTENNA_wire2202_A wire2202/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__255__A _255_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_273_ _273_/A _273_/B vssd vssd vccd vccd _273_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input83_A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__421__C _421_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output504_A wire1273/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1135_A wire1135/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_609_ _609_/A _609_/B vssd vssd vccd vccd _609_/X sky130_fd_sc_hd__and2_4
XFILLER_53_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1302_A _367_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output873_A _308_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__165__A _165_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] _179_/X vssd vssd vccd vccd _163_/A
+ sky130_fd_sc_hd__nand2_4
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] split5/X vssd vssd vccd vccd _143_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_31_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1671_A wire1672/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1769_A wire1769/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__612__B _612_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] _290_/X vssd vssd vccd vccd _110_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_2021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__379__A_N _507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__075__A _075_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_rebuffer6_A wire1460/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__522__B _522_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput780 wire1197/X vssd vssd vccd vccd la_oenb_core[3] sky130_fd_sc_hd__buf_8
Xwire2201 wire2202/X vssd vssd vccd vccd wire2201/X sky130_fd_sc_hd__buf_6
Xoutput791 wire1196/X vssd vssd vccd vccd la_oenb_core[4] sky130_fd_sc_hd__buf_8
Xwire2212 wire2213/X vssd vssd vccd vccd _481_/B sky130_fd_sc_hd__buf_6
XFILLER_40_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2223 wire2223/A vssd vssd vccd vccd wire2223/X sky130_fd_sc_hd__buf_6
XFILLER_47_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2234 wire2235/X vssd vssd vccd vccd _471_/B sky130_fd_sc_hd__buf_6
Xwire1500 wire1500/A vssd vssd vccd vccd wire1500/X sky130_fd_sc_hd__buf_6
Xwire2245 wire2245/A vssd vssd vccd vccd _464_/B sky130_fd_sc_hd__buf_6
Xwire1511 wire1511/A vssd vssd vccd vccd _368_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2256 wire2257/X vssd vssd vccd vccd wire2256/X sky130_fd_sc_hd__buf_6
XFILLER_48_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input235_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2152_A wire2152/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1522 wire1522/A vssd vssd vccd vccd _359_/B sky130_fd_sc_hd__buf_6
Xwire2267 wire2267/A vssd vssd vccd vccd wire2267/X sky130_fd_sc_hd__buf_6
XFILLER_4_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1533 wire1533/A vssd vssd vccd vccd wire1533/X sky130_fd_sc_hd__buf_6
XFILLER_19_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2278 wire2278/A vssd vssd vccd vccd _447_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1544 wire1545/X vssd vssd vccd vccd _347_/B sky130_fd_sc_hd__buf_6
Xwire2289 wire2290/X vssd vssd vccd vccd _437_/B sky130_fd_sc_hd__buf_6
XFILLER_38_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1555 wire1555/A vssd vssd vccd vccd wire1555/X sky130_fd_sc_hd__buf_6
XFILLER_21_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1566 wire1566/A vssd vssd vccd vccd wire1566/X sky130_fd_sc_hd__buf_6
XFILLER_21_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1577 wire1578/X vssd vssd vccd vccd _308_/B sky130_fd_sc_hd__buf_6
Xwire1588 wire1589/X vssd vssd vccd vccd wire1588/X sky130_fd_sc_hd__buf_6
XFILLER_46_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1599 wire1600/X vssd vssd vccd vccd wire1599/X sky130_fd_sc_hd__buf_6
XTAP_2110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input402_A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _325_/A _325_/B vssd vssd vccd vccd _325_/X sky130_fd_sc_hd__and2_1
XANTENNA__416__C _416_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_256_ _256_/A _256_/B vssd vssd vccd vccd _256_/X sky130_fd_sc_hd__and2_2
XFILLER_10_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_187_ _187_/A _187_/B vssd vssd vccd vccd _187_/X sky130_fd_sc_hd__and2_2
XFILLER_48_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__432__B _432_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1085_A _121_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output621_A _110_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output719_A wire1200/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3042 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1252_A _410_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1517_A wire1517/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__B _607_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1886_A wire1886/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__623__A _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__342__B _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[4\]_A mprj_dat_i_user[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__517__B _517_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_110_ _110_/A vssd vssd vccd vccd _110_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_36_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__533__A _533_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_041_ _041_/A vssd vssd vccd vccd _041_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input352_A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input46_A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2020 wire2021/X vssd vssd vccd vccd _615_/B sky130_fd_sc_hd__buf_6
Xwire2031 wire2031/A vssd vssd vccd vccd wire2031/X sky130_fd_sc_hd__buf_6
XFILLER_43_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2042 wire2043/X vssd vssd vccd vccd _607_/B sky130_fd_sc_hd__buf_6
Xwire2053 wire2053/A vssd vssd vccd vccd wire2053/X sky130_fd_sc_hd__buf_6
Xwire2064 wire2065/X vssd vssd vccd vccd _597_/B sky130_fd_sc_hd__buf_6
Xwire1330 _360_/X vssd vssd vccd vccd wire1330/X sky130_fd_sc_hd__buf_6
Xwire2075 wire2075/A vssd vssd vccd vccd wire2075/X sky130_fd_sc_hd__buf_6
Xwire1341 wire1342/X vssd vssd vccd vccd wire1341/X sky130_fd_sc_hd__buf_6
Xwire2086 wire2086/A vssd vssd vccd vccd _587_/B sky130_fd_sc_hd__buf_6
Xwire1352 wire1353/X vssd vssd vccd vccd wire1352/X sky130_fd_sc_hd__buf_6
Xwire2097 wire2098/X vssd vssd vccd vccd _581_/B sky130_fd_sc_hd__buf_6
XFILLER_46_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1363 _349_/X vssd vssd vccd vccd wire1363/X sky130_fd_sc_hd__buf_6
Xwire1374 wire1375/X vssd vssd vccd vccd wire1374/X sky130_fd_sc_hd__buf_6
Xwire1385 wire1386/X vssd vssd vccd vccd wire1385/X sky130_fd_sc_hd__buf_6
XFILLER_1_2558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1396 _337_/X vssd vssd vccd vccd wire1396/X sky130_fd_sc_hd__buf_6
XFILLER_46_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__427__B _427_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_308_ _308_/A _308_/B vssd vssd vccd vccd _308_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1000_A wire1001/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output571_A _451_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_239_ _239_/A _239_/B vssd vssd vccd vccd _239_/X sky130_fd_sc_hd__and2_4
XFILLER_45_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output836_A wire1146/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1467_A _255_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] wire1476/X vssd vssd vccd vccd wire1132/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1634_A wire1635/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1801_A wire1801/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__618__A _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__337__B _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__417__A_N _545_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__353__A _353_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput305 la_oenb_mprj[25] vssd vssd vccd vccd _522_/A sky130_fd_sc_hd__buf_4
Xinput316 la_oenb_mprj[35] vssd vssd vccd vccd wire1718/A sky130_fd_sc_hd__buf_6
XFILLER_22_4186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput327 la_oenb_mprj[45] vssd vssd vccd vccd _542_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput338 la_oenb_mprj[55] vssd vssd vccd vccd _552_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput349 la_oenb_mprj[65] vssd vssd vccd vccd wire1707/A sky130_fd_sc_hd__buf_6
XFILLER_2_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_590_ _590_/A _590_/B vssd vssd vccd vccd _590_/X sky130_fd_sc_hd__and2_4
XFILLER_2_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xload_slew1459 wire1460/X vssd vssd vccd vccd split5/A sky130_fd_sc_hd__buf_8
XFILLER_44_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__528__A _528_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input100_A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2115_A wire2116/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__263__A _263_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_024_ _024_/A vssd vssd vccd vccd _024_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_9 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1160 wire1161/X vssd vssd vccd vccd wire1160/X sky130_fd_sc_hd__buf_6
Xwire1171 _531_/X vssd vssd vccd vccd wire1171/X sky130_fd_sc_hd__buf_6
Xwire1182 _515_/X vssd vssd vccd vccd wire1182/X sky130_fd_sc_hd__buf_6
XFILLER_1_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1193 _504_/X vssd vssd vccd vccd wire1193/X sky130_fd_sc_hd__buf_6
XFILLER_35_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1048_A wire1049/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output786_A wire1164/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output953_A wire2302/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__173__A _173_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] rebuffer2/X vssd vssd vccd vccd _125_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_51_2991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1584_A wire1585/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1751_A wire1751/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1849_A wire1849/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__620__B _620_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_964 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__348__A _348_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__083__A _083_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__530__B _530_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput102 la_data_out_mprj[73] vssd vssd vccd vccd _442_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput113 la_data_out_mprj[83] vssd vssd vccd vccd wire1750/A sky130_fd_sc_hd__buf_6
XFILLER_24_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput124 la_data_out_mprj[93] vssd vssd vccd vccd _462_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2065_A wire2065/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input148_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput135 la_iena_mprj[102] vssd vssd vccd vccd _265_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput146 la_iena_mprj[112] vssd vssd vccd vccd _275_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 la_iena_mprj[122] vssd vssd vccd vccd _285_/B sky130_fd_sc_hd__buf_4
XTAP_4634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 la_iena_mprj[17] vssd vssd vccd vccd _180_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 la_iena_mprj[27] vssd vssd vccd vccd _190_/B sky130_fd_sc_hd__buf_4
XFILLER_29_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2232_A wire2233/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input315_A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__258__A _258_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_573_ _573_/A _573_/B vssd vssd vccd vccd _573_/X sky130_fd_sc_hd__and2_4
XTAP_3988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_B split5/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2942 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__424__C _424_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput609 _099_/Y vssd vssd vccd vccd la_data_in_mprj[116] sky130_fd_sc_hd__buf_8
XFILLER_29_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_007_ _007_/A vssd vssd vccd vccd _007_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_46_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__440__B _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output534_A wire1244/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1332_A wire1333/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__168__A _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] _209_/X vssd vssd vccd vccd _029_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_36_967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_B load_slew1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1799_A wire1799/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__615__B _615_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] _171_/X vssd vssd vccd vccd _155_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_28_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__350__B _350_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1907 wire1908/X vssd vssd vccd vccd _261_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1918 wire1918/A vssd vssd vccd vccd _252_/A sky130_fd_sc_hd__buf_6
XFILLER_3_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1929 wire1929/A vssd vssd vccd vccd _298_/A sky130_fd_sc_hd__buf_6
XTAP_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_207 _337_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__078__A _078_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 wire2077/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 wire2193/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[12\]_B split4/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__525__B _525_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_672 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__541__A _541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2182_A wire2183/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input265_A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__260__B _260_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input432_A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_625_ _625_/A _625_/B vssd vssd vccd vccd _625_/X sky130_fd_sc_hd__and2_1
XTAP_3763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_556_ _556_/A _556_/B vssd vssd vccd vccd _556_/X sky130_fd_sc_hd__and2_4
XFILLER_45_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_487_ _615_/A _487_/B _487_/C vssd vssd vccd vccd _487_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__435__B _435_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output484_A _488_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3782 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2658 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output651_A _022_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output749_A wire1143/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1282_A _381_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output916_A wire1361/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1547_A wire1548/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__345__B _345_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__361__A _361_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput940 wire1382/X vssd vssd vccd vccd mprj_dat_o_user[5] sky130_fd_sc_hd__buf_8
XFILLER_5_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput951 wire1838/X vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_25_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1704 wire1704/A vssd vssd vccd vccd _565_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1715 _409_/A_N vssd vssd vccd vccd _537_/A sky130_fd_sc_hd__buf_4
XFILLER_41_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1726 wire1726/A vssd vssd vccd vccd _618_/A sky130_fd_sc_hd__buf_6
XTAP_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1737 input24/X vssd vssd vccd vccd _487_/C sky130_fd_sc_hd__buf_6
XTAP_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1748 wire1748/A vssd vssd vccd vccd _454_/C sky130_fd_sc_hd__buf_6
XFILLER_3_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1759 wire1759/A vssd vssd vccd vccd _392_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _538_/A _410_/B _410_/C vssd vssd vccd vccd _410_/X sky130_fd_sc_hd__and3b_4
XTAP_2347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2028_A wire2028/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_341_ _341_/A _341_/B vssd vssd vccd vccd _341_/X sky130_fd_sc_hd__and2_2
XFILLER_36_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_272_ _272_/A _272_/B vssd vssd vccd vccd _272_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3922 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input382_A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input76_A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__271__A _271_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_608_ _608_/A _608_/B vssd vssd vccd vccd _608_/X sky130_fd_sc_hd__and2_4
XTAP_3593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1030_A _132_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1128_A wire1128/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_539_ _539_/A _539_/B vssd vssd vccd vccd _539_/X sky130_fd_sc_hd__and2_4
XTAP_2892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__450__A_N _578_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output866_A _331_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1497_A wire1498/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__181__A _181_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1664_A wire1665/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1831_A wire1831/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1929_A wire1929/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__356__A _356_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4438 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__091__A _091_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput770 _527_/X vssd vssd vccd vccd la_oenb_core[30] sky130_fd_sc_hd__buf_8
Xoutput781 _537_/X vssd vssd vccd vccd la_oenb_core[40] sky130_fd_sc_hd__buf_8
XFILLER_47_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2202 wire2202/A vssd vssd vccd vccd wire2202/X sky130_fd_sc_hd__buf_6
Xoutput792 wire1160/X vssd vssd vccd vccd la_oenb_core[50] sky130_fd_sc_hd__buf_8
Xwire2213 wire2214/X vssd vssd vccd vccd wire2213/X sky130_fd_sc_hd__buf_6
Xwire2224 wire2225/X vssd vssd vccd vccd _476_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2235 wire2235/A vssd vssd vccd vccd wire2235/X sky130_fd_sc_hd__buf_6
XFILLER_25_2760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1501 wire1502/X vssd vssd vccd vccd _344_/B sky130_fd_sc_hd__buf_6
Xwire2246 wire2246/A vssd vssd vccd vccd _463_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1512 wire1512/A vssd vssd vccd vccd _367_/B sky130_fd_sc_hd__buf_6
Xwire2257 wire2257/A vssd vssd vccd vccd wire2257/X sky130_fd_sc_hd__buf_6
XFILLER_38_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1523 wire1523/A vssd vssd vccd vccd _358_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2268 wire2269/X vssd vssd vccd vccd _452_/B sky130_fd_sc_hd__buf_6
XFILLER_48_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1534 wire1535/X vssd vssd vccd vccd _352_/B sky130_fd_sc_hd__buf_6
Xwire2279 wire2279/A vssd vssd vccd vccd _446_/B sky130_fd_sc_hd__buf_6
XFILLER_4_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1545 wire1545/A vssd vssd vccd vccd wire1545/X sky130_fd_sc_hd__buf_6
XFILLER_19_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input130_A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1556 wire1557/X vssd vssd vccd vccd _313_/B sky130_fd_sc_hd__buf_6
XFILLER_38_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2145_A wire2145/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1567 wire1568/X vssd vssd vccd vccd _310_/B sky130_fd_sc_hd__buf_6
XANTENNA_input228_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1578 wire1579/X vssd vssd vccd vccd wire1578/X sky130_fd_sc_hd__buf_6
XFILLER_0_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1589 wire1590/X vssd vssd vccd vccd wire1589/X sky130_fd_sc_hd__buf_6
XTAP_2100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__473__A_N _601_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__266__A _266_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ _324_/A _324_/B vssd vssd vccd vccd _324_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_255_ _255_/A _255_/B vssd vssd vccd vccd _255_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_186_ _186_/A _186_/B vssd vssd vccd vccd _186_/X sky130_fd_sc_hd__and2_1
XFILLER_45_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__432__C _432_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1078_A wire1079/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1245_A _417_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1412_A wire1413/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__176__A _176_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1781_A wire1781/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1879_A wire1880/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__623__B _623_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[4\]_B split4/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__496__A_N _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__086__A _086_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_040_ _040_/A vssd vssd vccd vccd _040_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__533__B _533_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2095_A wire2096/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input178_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input345_A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2262_A wire2263/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2010 wire2011/X vssd vssd vccd vccd _618_/B sky130_fd_sc_hd__buf_6
Xwire2021 wire2022/X vssd vssd vccd vccd wire2021/X sky130_fd_sc_hd__buf_6
Xwire2032 wire2033/X vssd vssd vccd vccd _611_/B sky130_fd_sc_hd__buf_6
XFILLER_25_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input39_A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2043 wire2044/X vssd vssd vccd vccd wire2043/X sky130_fd_sc_hd__buf_6
Xwire2054 wire2055/X vssd vssd vccd vccd _602_/B sky130_fd_sc_hd__buf_6
XFILLER_5_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1320 wire1321/X vssd vssd vccd vccd wire1320/X sky130_fd_sc_hd__buf_6
Xwire2065 wire2065/A vssd vssd vccd vccd wire2065/X sky130_fd_sc_hd__buf_6
Xwire1331 wire1332/X vssd vssd vccd vccd wire1331/X sky130_fd_sc_hd__buf_8
Xwire2076 wire2077/X vssd vssd vccd vccd _593_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2087 wire2087/A vssd vssd vccd vccd _586_/B sky130_fd_sc_hd__buf_6
Xwire1342 _356_/X vssd vssd vccd vccd wire1342/X sky130_fd_sc_hd__buf_6
XFILLER_1_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1353 wire1354/X vssd vssd vccd vccd wire1353/X sky130_fd_sc_hd__buf_6
Xwire2098 wire2098/A vssd vssd vccd vccd wire2098/X sky130_fd_sc_hd__buf_6
Xwire1364 wire1365/X vssd vssd vccd vccd wire1364/X sky130_fd_sc_hd__buf_6
XFILLER_5_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1375 _345_/X vssd vssd vccd vccd wire1375/X sky130_fd_sc_hd__buf_6
Xwire1386 wire1387/X vssd vssd vccd vccd wire1386/X sky130_fd_sc_hd__buf_6
XFILLER_19_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1397 _328_/X vssd vssd vccd vccd wire1397/X sky130_fd_sc_hd__buf_6
XFILLER_1_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__427__C _427_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_307_ _307_/A _307_/B vssd vssd vccd vccd _307_/X sky130_fd_sc_hd__and2_4
XFILLER_50_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_238_ _238_/A _238_/B vssd vssd vccd vccd _238_/X sky130_fd_sc_hd__and2_4
XANTENNA__443__B _443_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output564_A _445_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__369__A_N _497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_169_ _169_/A _169_/B vssd vssd vccd vccd _169_/X sky130_fd_sc_hd__and2_2
XFILLER_32_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1195_A _502_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output731_A _607_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output829_A _581_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1362_A wire1363/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] _239_/X vssd vssd vccd vccd _059_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1627_A wire1628/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__618__B _618_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1996_A wire1997/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire982_A wire983/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__353__B _353_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput306 la_oenb_mprj[26] vssd vssd vccd vccd _523_/A sky130_fd_sc_hd__buf_4
XFILLER_22_4176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput317 la_oenb_mprj[36] vssd vssd vccd vccd _405_/A_N sky130_fd_sc_hd__buf_6
Xinput328 la_oenb_mprj[46] vssd vssd vccd vccd _543_/A sky130_fd_sc_hd__buf_8
XFILLER_22_4198 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput339 la_oenb_mprj[56] vssd vssd vccd vccd _553_/A sky130_fd_sc_hd__buf_4
XFILLER_29_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_884 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2010_A wire2011/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__544__A _544_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_16_2589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input295_A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__263__B _263_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_023_ _023_/A vssd vssd vccd vccd _023_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input462_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1150 wire1151/X vssd vssd vccd vccd wire1150/X sky130_fd_sc_hd__buf_6
XFILLER_1_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1161 _547_/X vssd vssd vccd vccd wire1161/X sky130_fd_sc_hd__buf_6
XFILLER_40_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1172 _530_/X vssd vssd vccd vccd wire1172/X sky130_fd_sc_hd__buf_6
XFILLER_21_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1183 _514_/X vssd vssd vccd vccd wire1183/X sky130_fd_sc_hd__buf_6
XFILLER_34_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1194 _503_/X vssd vssd vccd vccd wire1194/X sky130_fd_sc_hd__buf_6
XFILLER_5_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__438__B _438_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1110_A _116_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output681_A _049_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output779_A wire1169/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4080 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output946_A wire1435/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1577_A wire1578/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1911_A wire1911/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] _265_/X vssd vssd vccd vccd _085_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__348__B _348_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__364__A _364_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_2767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput103 la_data_out_mprj[74] vssd vssd vccd vccd _443_/C sky130_fd_sc_hd__buf_4
Xinput114 la_data_out_mprj[84] vssd vssd vccd vccd wire1749/A sky130_fd_sc_hd__buf_6
XFILLER_49_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput125 la_data_out_mprj[94] vssd vssd vccd vccd _463_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 la_iena_mprj[103] vssd vssd vccd vccd _266_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput147 la_iena_mprj[113] vssd vssd vccd vccd _276_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput158 la_iena_mprj[123] vssd vssd vccd vccd _286_/B sky130_fd_sc_hd__buf_4
XFILLER_5_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2058_A wire2059/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput169 la_iena_mprj[18] vssd vssd vccd vccd _181_/B sky130_fd_sc_hd__buf_4
XTAP_4646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__539__A _539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input210_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_572_ _572_/A _572_/B vssd vssd vccd vccd _572_/X sky130_fd_sc_hd__and2_4
XTAP_3978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2225_A wire2225/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input308_A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2954 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3931 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__274__A _274_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_006_ _006_/A vssd vssd vccd vccd _006_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_2725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__440__C _440_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__407__A_N _535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output527_A wire1251/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1060_A _126_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1158_A wire1159/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1325_A wire1326/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output896_A wire1002/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] _202_/X vssd vssd vccd vccd _022_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_14_3728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__184__A _184_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1694_A _447_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1861_A wire1862/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1959_A wire1960/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1908 wire1908/A vssd vssd vccd vccd wire1908/X sky130_fd_sc_hd__buf_6
XTAP_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1919 wire1919/A vssd vssd vccd vccd _251_/A sky130_fd_sc_hd__buf_6
XFILLER_41_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__359__A _359_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _314_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 wire2079/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__094__A _094_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_150 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_684 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__541__B _541_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input160_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input258_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2175_A wire2175/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input425_A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__269__A _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_624_ _624_/A _624_/B vssd vssd vccd vccd _624_/X sky130_fd_sc_hd__and2_2
XTAP_4498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_555_ _555_/A _555_/B vssd vssd vccd vccd _555_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_938 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_486_ _614_/A _486_/B _486_/C vssd vssd vccd vccd _486_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__435__C _435_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3794 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output477_A _481_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__451__B _451_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output644_A _015_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1275_A _388_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output811_A _565_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output909_A wire1086/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1442_A wire1443/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3754 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__179__A _179_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1707_A wire1707/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_702 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__361__B _361_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput930 wire1319/X vssd vssd vccd vccd mprj_dat_o_user[25] sky130_fd_sc_hd__buf_8
XFILLER_25_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput941 wire1379/X vssd vssd vccd vccd mprj_dat_o_user[6] sky130_fd_sc_hd__buf_8
XFILLER_8_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput952 output952/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_5_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1705 wire1705/A vssd vssd vccd vccd _564_/A sky130_fd_sc_hd__buf_6
XFILLER_3_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1716 _406_/A_N vssd vssd vccd vccd _534_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1727 wire1727/A vssd vssd vccd vccd _617_/A sky130_fd_sc_hd__buf_6
XTAP_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1738 input23/X vssd vssd vccd vccd _486_/C sky130_fd_sc_hd__buf_6
XTAP_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__089__A _089_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1749 wire1749/A vssd vssd vccd vccd _453_/C sky130_fd_sc_hd__buf_6
XTAP_3005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _340_/A _340_/B vssd vssd vccd vccd _340_/X sky130_fd_sc_hd__and2_2
XFILLER_41_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__536__B _536_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_271_ _271_/A _271_/B vssd vssd vccd vccd _271_/X sky130_fd_sc_hd__and2_4
XFILLER_23_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3934 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__552__A _552_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2292_A wire2292/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input375_A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input69_A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_607_ _607_/A _607_/B vssd vssd vccd vccd _607_/X sky130_fd_sc_hd__and2_4
XFILLER_45_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__446__B _446_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1023_A wire1024/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_538_ _538_/A _538_/B vssd vssd vccd vccd _538_/X sky130_fd_sc_hd__and2_2
XTAP_2893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output594_A _085_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_469_ _597_/A _469_/B _469_/C vssd vssd vccd vccd _469_/X sky130_fd_sc_hd__and3b_2
XFILLER_32_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output761_A wire1178/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output859_A _306_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1392_A _339_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__181__B _181_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1657_A wire1658/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1824_A wire1824/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4083 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__356__B _356_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_B _257_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput760 wire1179/X vssd vssd vccd vccd la_oenb_core[21] sky130_fd_sc_hd__buf_8
XFILLER_5_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput771 _528_/X vssd vssd vccd vccd la_oenb_core[31] sky130_fd_sc_hd__buf_8
XFILLER_40_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput782 wire1167/X vssd vssd vccd vccd la_oenb_core[41] sky130_fd_sc_hd__buf_8
XFILLER_8_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2203 wire2204/X vssd vssd vccd vccd _484_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput793 _548_/X vssd vssd vccd vccd la_oenb_core[51] sky130_fd_sc_hd__buf_8
XFILLER_47_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2214 wire2214/A vssd vssd vccd vccd wire2214/X sky130_fd_sc_hd__buf_6
XFILLER_21_3315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2225 wire2225/A vssd vssd vccd vccd wire2225/X sky130_fd_sc_hd__buf_6
XFILLER_28_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2236 wire2236/A vssd vssd vccd vccd _470_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1502 wire1502/A vssd vssd vccd vccd wire1502/X sky130_fd_sc_hd__buf_6
Xwire2247 wire2247/A vssd vssd vccd vccd _462_/B sky130_fd_sc_hd__buf_4
XFILLER_25_2772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1513 wire1514/X vssd vssd vccd vccd _339_/B sky130_fd_sc_hd__buf_6
Xwire2258 wire2259/X vssd vssd vccd vccd _455_/B sky130_fd_sc_hd__buf_6
Xwire1524 wire1524/A vssd vssd vccd vccd _357_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2269 wire2270/X vssd vssd vccd vccd wire2269/X sky130_fd_sc_hd__buf_6
Xwire1535 wire1535/A vssd vssd vccd vccd wire1535/X sky130_fd_sc_hd__buf_6
Xwire1546 wire1547/X vssd vssd vccd vccd _337_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1557 wire1558/X vssd vssd vccd vccd wire1557/X sky130_fd_sc_hd__buf_6
XFILLER_24_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1568 wire1569/X vssd vssd vccd vccd wire1568/X sky130_fd_sc_hd__buf_6
XFILLER_38_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1579 wire1580/X vssd vssd vccd vccd wire1579/X sky130_fd_sc_hd__buf_6
XANTENNA_input123_A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2040_A wire2041/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2138_A wire2138/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__547__A _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__266__B _266_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2305_A wire2306/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_323_ _323_/A _323_/B vssd vssd vccd vccd _323_/X sky130_fd_sc_hd__and2_2
XFILLER_42_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[85\]_B wire1474/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_254_ _254_/A _254_/B vssd vssd vccd vccd _254_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__282__A _282_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_185_ _185_/A _185_/B vssd vssd vccd vccd _185_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2798 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] split4/X vssd vssd vccd vccd _118_/A sky130_fd_sc_hd__nand2_4
XFILLER_7_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1238_A wire1239/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1405_A _322_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] _184_/X vssd vssd vccd vccd _004_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_20_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[76\]_B _239_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__192__A _192_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1774_A wire1775/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1941_A wire1941/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__367__A _367_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2088_A wire2089/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2000 wire2000/A vssd vssd vccd vccd wire2000/X sky130_fd_sc_hd__buf_6
XFILLER_27_2867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput590 wire1285/X vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__buf_8
XFILLER_44_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2011 wire2012/X vssd vssd vccd vccd wire2011/X sky130_fd_sc_hd__buf_6
XFILLER_47_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2022 wire2022/A vssd vssd vccd vccd wire2022/X sky130_fd_sc_hd__buf_6
XANTENNA_input240_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2033 wire2034/X vssd vssd vccd vccd wire2033/X sky130_fd_sc_hd__buf_6
XFILLER_21_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input338_A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2044 wire2044/A vssd vssd vccd vccd wire2044/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2255_A wire2256/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2055 wire2055/A vssd vssd vccd vccd wire2055/X sky130_fd_sc_hd__buf_6
Xwire1310 _365_/X vssd vssd vccd vccd wire1310/X sky130_fd_sc_hd__buf_6
XFILLER_40_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__440__A_N _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1321 wire1322/X vssd vssd vccd vccd wire1321/X sky130_fd_sc_hd__buf_6
Xwire2066 wire2067/X vssd vssd vccd vccd _596_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2422 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1332 wire1333/X vssd vssd vccd vccd wire1332/X sky130_fd_sc_hd__buf_6
XFILLER_8_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2077 wire2077/A vssd vssd vccd vccd wire2077/X sky130_fd_sc_hd__buf_6
Xwire1343 wire1344/X vssd vssd vccd vccd wire1343/X sky130_fd_sc_hd__buf_6
XFILLER_38_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2088 wire2089/X vssd vssd vccd vccd _585_/B sky130_fd_sc_hd__buf_6
Xwire2099 wire2100/X vssd vssd vccd vccd _580_/B sky130_fd_sc_hd__buf_6
Xwire1354 _352_/X vssd vssd vccd vccd wire1354/X sky130_fd_sc_hd__buf_6
Xwire1365 wire1366/X vssd vssd vccd vccd wire1365/X sky130_fd_sc_hd__buf_6
XFILLER_19_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1376 wire1377/X vssd vssd vccd vccd wire1376/X sky130_fd_sc_hd__buf_6
XFILLER_38_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1387 _341_/X vssd vssd vccd vccd wire1387/X sky130_fd_sc_hd__buf_6
Xwire1398 wire1399/X vssd vssd vccd vccd wire1398/X sky130_fd_sc_hd__buf_6
XANTENNA__277__A _277_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3853 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_306_ _306_/A _306_/B vssd vssd vccd vccd _306_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_237_ _237_/A _237_/B vssd vssd vccd vccd _237_/X sky130_fd_sc_hd__and2_4
XANTENNA__443__C _443_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_168_ _168_/A _168_/B vssd vssd vccd vccd _168_/X sky130_fd_sc_hd__and2_1
XANTENNA_output557_A wire1288/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_099_ _099_/A vssd vssd vccd vccd _099_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_3900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output724_A _601_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1355_A wire1356/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] _232_/X vssd vssd vccd vccd _052_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1522_A wire1522/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__187__A _187_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4015 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1891_A wire1892/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1989_A wire1989/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire975_A wire976/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__463__A_N _591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput307 la_oenb_mprj[27] vssd vssd vccd vccd _524_/A sky130_fd_sc_hd__clkbuf_8
Xinput318 la_oenb_mprj[37] vssd vssd vccd vccd _406_/A_N sky130_fd_sc_hd__buf_6
XFILLER_9_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput329 la_oenb_mprj[47] vssd vssd vccd vccd _416_/A_N sky130_fd_sc_hd__buf_6
XFILLER_44_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__097__A _097_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__544__B _544_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_B _287_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input190_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input288_A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_022_ _022_/A vssd vssd vccd vccd _022_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__A _560_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input455_A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input51_A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1140 wire1140/A vssd vssd vccd vccd _105_/A sky130_fd_sc_hd__buf_6
Xwire1151 _555_/X vssd vssd vccd vccd wire1151/X sky130_fd_sc_hd__buf_6
Xwire1162 wire1163/X vssd vssd vccd vccd wire1162/X sky130_fd_sc_hd__buf_6
XFILLER_5_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1173 _525_/X vssd vssd vccd vccd wire1173/X sky130_fd_sc_hd__buf_6
Xwire1184 _513_/X vssd vssd vccd vccd wire1184/X sky130_fd_sc_hd__buf_6
XFILLER_38_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1195 _502_/X vssd vssd vccd vccd wire1195/X sky130_fd_sc_hd__buf_6
XANTENNA__438__C _438_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_638 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3915 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__454__B _454_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[115\]_B _278_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1103_A wire1104/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4092 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__486__A_N _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output841_A _592_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output939_A wire1385/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1472_A _250_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[24\]_A mprj_dat_i_user[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__364__B _364_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_B wire1462/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1731 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput104 la_data_out_mprj[75] vssd vssd vccd vccd _444_/C sky130_fd_sc_hd__buf_4
XFILLER_4_2909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput115 la_data_out_mprj[85] vssd vssd vccd vccd wire1748/A sky130_fd_sc_hd__buf_6
Xinput126 la_data_out_mprj[95] vssd vssd vccd vccd _464_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 la_iena_mprj[104] vssd vssd vccd vccd _267_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 la_iena_mprj[114] vssd vssd vccd vccd _277_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput159 la_iena_mprj[124] vssd vssd vccd vccd _287_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__539__B _539_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[15\]_A mprj_dat_i_user[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_571_ _571_/A _571_/B vssd vssd vccd vccd _571_/X sky130_fd_sc_hd__and2_4
XTAP_3968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input203_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2218_A wire2219/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__555__A _555_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3943 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input99_A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__A _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_005_ _005_/A vssd vssd vccd vccd _005_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__449__B _449_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1053_A wire1054/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1220_A _462_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output791_A wire1196/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output889_A wire1031/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__184__B _184_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_4198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1687_A wire1687/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1854_A wire1855/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1909 wire1910/X vssd vssd vccd vccd _260_/A sky130_fd_sc_hd__buf_6
XTAP_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__359__B _359_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 wire1649/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2070_A wire2071/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input153_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2168_A wire2168/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__269__B _269_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input320_A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input418_A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_623_ _623_/A _623_/B vssd vssd vccd vccd _623_/X sky130_fd_sc_hd__and2_2
XFILLER_22_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_554_ _554_/A _554_/B vssd vssd vccd vccd _554_/X sky130_fd_sc_hd__and2_2
XTAP_3798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__285__A _285_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_485_ _613_/A _485_/B _485_/C vssd vssd vccd vccd _485_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2086 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__451__C _451_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1170_A _535_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output804_A wire1148/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__179__B _179_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3766 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1435_A wire1436/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] _214_/X vssd vssd vccd vccd _034_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_40_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1602_A wire1603/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_714 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__195__A _195_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput920 wire1349/X vssd vssd vccd vccd mprj_dat_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_2_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput931 wire1315/X vssd vssd vccd vccd mprj_dat_o_user[26] sky130_fd_sc_hd__buf_8
XFILLER_9_3852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput942 wire1376/X vssd vssd vccd vccd mprj_dat_o_user[7] sky130_fd_sc_hd__buf_8
XFILLER_25_4367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput953 wire2302/X vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_45_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input6_A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1706 wire1706/A vssd vssd vccd vccd _563_/A sky130_fd_sc_hd__buf_6
XTAP_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1717 _405_/A_N vssd vssd vccd vccd _533_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1728 wire1728/A vssd vssd vccd vccd _616_/A sky130_fd_sc_hd__buf_6
XTAP_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1739 input22/X vssd vssd vccd vccd _485_/C sky130_fd_sc_hd__buf_6
XFILLER_3_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_270_ _270_/A _270_/B vssd vssd vccd vccd _270_/X sky130_fd_sc_hd__and2_4
XFILLER_41_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_460 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__552__B _552_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input270_A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2092 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2285_A wire2285/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input368_A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_606_ _606_/A _606_/B vssd vssd vccd vccd _606_/X sky130_fd_sc_hd__and2_4
XTAP_3573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3960 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_537_ _537_/A _537_/B vssd vssd vccd vccd _537_/X sky130_fd_sc_hd__and2_4
XTAP_2872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__446__C _446_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_468_ _596_/A _468_/B _468_/C vssd vssd vccd vccd _468_/X sky130_fd_sc_hd__and3b_1
XANTENNA_wire1016_A wire1017/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output587_A _466_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_399_ _527_/A _399_/B _399_/C vssd vssd vccd vccd _399_/X sky130_fd_sc_hd__and3b_2
XFILLER_31_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__462__B _462_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output754_A wire1184/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1385_A wire1386/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output921_A wire1346/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] _262_/X vssd vssd vccd vccd wire1121/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_29_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1552_A wire1552/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1817_A wire1817/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2070 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__372__B _372_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[7\]_A mprj_dat_i_user[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_4175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput750 wire1188/X vssd vssd vccd vccd la_oenb_core[12] sky130_fd_sc_hd__buf_8
Xoutput761 wire1178/X vssd vssd vccd vccd la_oenb_core[22] sky130_fd_sc_hd__buf_8
Xoutput772 _529_/X vssd vssd vccd vccd la_oenb_core[32] sky130_fd_sc_hd__buf_8
XFILLER_5_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput783 wire1166/X vssd vssd vccd vccd la_oenb_core[42] sky130_fd_sc_hd__buf_8
XFILLER_40_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2204 wire2205/X vssd vssd vccd vccd wire2204/X sky130_fd_sc_hd__buf_6
Xoutput794 wire1158/X vssd vssd vccd vccd la_oenb_core[52] sky130_fd_sc_hd__buf_8
XFILLER_5_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2215 wire2216/X vssd vssd vccd vccd _480_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2226 wire2227/X vssd vssd vccd vccd _475_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2237 wire2238/X vssd vssd vccd vccd _469_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1503 wire1504/X vssd vssd vccd vccd _343_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2248 wire2248/A vssd vssd vccd vccd _461_/B sky130_fd_sc_hd__buf_6
Xwire1514 wire1514/A vssd vssd vccd vccd wire1514/X sky130_fd_sc_hd__buf_6
XFILLER_43_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2259 wire2260/X vssd vssd vccd vccd wire2259/X sky130_fd_sc_hd__buf_6
XFILLER_24_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1525 wire1526/X vssd vssd vccd vccd _338_/B sky130_fd_sc_hd__buf_6
XTAP_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1536 wire1537/X vssd vssd vccd vccd _351_/B sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1547 wire1548/X vssd vssd vccd vccd wire1547/X sky130_fd_sc_hd__buf_6
XFILLER_41_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1558 wire1559/X vssd vssd vccd vccd wire1558/X sky130_fd_sc_hd__buf_6
Xwire1569 wire1570/X vssd vssd vccd vccd wire1569/X sky130_fd_sc_hd__buf_6
XFILLER_38_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__547__B _547_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2033_A wire2034/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _322_/A _322_/B vssd vssd vccd vccd _322_/X sky130_fd_sc_hd__and2_2
XTAP_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2200_A wire2201/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__563__A _563_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_253_ _253_/A _253_/B vssd vssd vccd vccd _253_/X sky130_fd_sc_hd__and2_2
XFILLER_10_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__282__B _282_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input81_A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_184_ _184_/A _184_/B vssd vssd vccd vccd _184_/X sky130_fd_sc_hd__and2_2
XFILLER_10_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output502_A wire1293/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__457__B _457_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1133_A wire1133/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1300_A wire1301/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output871_A _335_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] split5/X vssd vssd vccd vccd _141_/A
+ sky130_fd_sc_hd__nand2_4
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] _177_/X vssd vssd vccd vccd _161_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_33_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__192__B _192_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1767_A wire1767/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1934_A wire1934/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] _288_/X vssd vssd vccd vccd _108_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_20_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__367__B _367_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3418 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__A_N _520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2608 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_4309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput580 wire1223/X vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__buf_8
XFILLER_40_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2001 wire2002/X vssd vssd vccd vccd _621_/B sky130_fd_sc_hd__buf_6
Xoutput591 _147_/Y vssd vssd vccd vccd la_data_in_mprj[0] sky130_fd_sc_hd__buf_8
Xwire2012 wire2012/A vssd vssd vccd vccd wire2012/X sky130_fd_sc_hd__buf_6
XFILLER_27_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2023 wire2024/X vssd vssd vccd vccd _614_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2034 wire2034/A vssd vssd vccd vccd wire2034/X sky130_fd_sc_hd__buf_6
Xwire1300 wire1301/X vssd vssd vccd vccd wire1300/X sky130_fd_sc_hd__buf_6
Xwire2045 wire2046/X vssd vssd vccd vccd _606_/B sky130_fd_sc_hd__buf_6
Xwire1311 wire1312/X vssd vssd vccd vccd wire1311/X sky130_fd_sc_hd__buf_8
Xwire2056 wire2057/X vssd vssd vccd vccd _601_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2067 wire2067/A vssd vssd vccd vccd wire2067/X sky130_fd_sc_hd__buf_6
Xwire1322 _362_/X vssd vssd vccd vccd wire1322/X sky130_fd_sc_hd__buf_6
Xwire2078 wire2079/X vssd vssd vccd vccd _592_/B sky130_fd_sc_hd__buf_6
XANTENNA_input233_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1333 _359_/X vssd vssd vccd vccd wire1333/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2248_A wire2248/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1344 wire1345/X vssd vssd vccd vccd wire1344/X sky130_fd_sc_hd__buf_6
XFILLER_5_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2089 wire2089/A vssd vssd vccd vccd wire2089/X sky130_fd_sc_hd__buf_6
Xwire1355 wire1356/X vssd vssd vccd vccd wire1355/X sky130_fd_sc_hd__buf_6
XFILLER_38_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__558__A _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1366 _348_/X vssd vssd vccd vccd wire1366/X sky130_fd_sc_hd__buf_6
Xwire1377 wire1378/X vssd vssd vccd vccd wire1377/X sky130_fd_sc_hd__buf_6
Xwire1388 wire1389/X vssd vssd vccd vccd wire1388/X sky130_fd_sc_hd__buf_6
XFILLER_35_809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1399 _327_/X vssd vssd vccd vccd wire1399/X sky130_fd_sc_hd__buf_6
XANTENNA_input400_A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__277__B _277_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__293__A _293_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_305_ _305_/A _305_/B vssd vssd vccd vccd _305_/X sky130_fd_sc_hd__and2_4
XFILLER_15_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_236_ _236_/A _236_/B vssd vssd vccd vccd _236_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_167_ _167_/A _167_/B vssd vssd vccd vccd _167_/X sky130_fd_sc_hd__and2_1
XFILLER_10_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_098_ _098_/A vssd vssd vccd vccd _098_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1083_A wire1084/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output717_A _082_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1250_A _412_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1348_A _354_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__187__B _187_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1884_A wire1884/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire968_A wire969/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput308 la_oenb_mprj[28] vssd vssd vccd vccd _525_/A sky130_fd_sc_hd__buf_4
XFILLER_29_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput319 la_oenb_mprj[38] vssd vssd vccd vccd _535_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1103 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_021_ _021_/A vssd vssd vccd vccd _021_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input183_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2198_A wire2199/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__B _560_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input350_A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input448_A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input44_A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1130 wire1130/A vssd vssd vccd vccd _068_/A sky130_fd_sc_hd__buf_6
XFILLER_40_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1141 wire1141/A vssd vssd vccd vccd _104_/A sky130_fd_sc_hd__buf_6
XANTENNA__288__A _288_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1152 _554_/X vssd vssd vccd vccd wire1152/X sky130_fd_sc_hd__buf_6
XFILLER_38_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1163 _546_/X vssd vssd vccd vccd wire1163/X sky130_fd_sc_hd__buf_6
XFILLER_19_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1174 _523_/X vssd vssd vccd vccd wire1174/X sky130_fd_sc_hd__buf_6
XFILLER_21_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1185 _512_/X vssd vssd vccd vccd wire1185/X sky130_fd_sc_hd__buf_6
XFILLER_34_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1196 _501_/X vssd vssd vccd vccd wire1196/X sky130_fd_sc_hd__buf_6
XFILLER_35_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__454__C _454_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_219_ _219_/A _219_/B vssd vssd vccd vccd _219_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__B _470_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output834_A wire1147/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1465_A _258_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] wire1478/X vssd vssd vccd vccd wire1134/A
+ sky130_fd_sc_hd__nand2_8
XTAP_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__198__A _198_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_138 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3546 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2747 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__430__A_N _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__380__B _380_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_749 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput105 la_data_out_mprj[76] vssd vssd vccd vccd _445_/C sky130_fd_sc_hd__buf_4
Xinput116 la_data_out_mprj[86] vssd vssd vccd vccd wire1747/A sky130_fd_sc_hd__buf_6
XFILLER_44_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput127 la_data_out_mprj[96] vssd vssd vccd vccd _465_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 la_iena_mprj[105] vssd vssd vccd vccd _268_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput149 la_iena_mprj[115] vssd vssd vccd vccd _278_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[15\]_B load_slew1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_570_ _570_/A _570_/B vssd vssd vccd vccd _570_/X sky130_fd_sc_hd__and2_4
XTAP_3958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2024 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__555__B _555_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2113_A wire2114/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input398_A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__571__A _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_004_ _004_/A vssd vssd vccd vccd _004_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__B _290_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__449__C _449_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1046_A wire1047/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3833 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__465__B _465_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1213_A _471_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__453__A_N _581_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output784_A _540_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output951_A wire1838/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1582_A wire1583/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1847_A wire1848/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__375__B _375_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_max_length1714_A _416_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2063_A wire2063/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input146_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_622_ _622_/A _622_/B vssd vssd vccd vccd _622_/X sky130_fd_sc_hd__and2_4
XTAP_4478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2230_A wire2231/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2464 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input313_A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__476__A_N _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__566__A _566_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_553_ _553_/A _553_/B vssd vssd vccd vccd _553_/X sky130_fd_sc_hd__and2_2
XTAP_3788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__285__B _285_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_484_ _612_/A _484_/B _484_/C vssd vssd vccd vccd _484_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2098 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output532_A wire1246/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1428_A wire1429/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] _207_/X vssd vssd vccd vccd _027_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_35_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__195__B _195_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1797_A wire1797/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput910 wire1081/X vssd vssd vccd vccd mprj_dat_i_core[7] sky130_fd_sc_hd__buf_8
Xoutput921 wire1346/X vssd vssd vccd vccd mprj_dat_o_user[17] sky130_fd_sc_hd__buf_8
Xoutput932 wire1311/X vssd vssd vccd vccd mprj_dat_o_user[27] sky130_fd_sc_hd__buf_8
Xoutput943 wire1373/X vssd vssd vccd vccd mprj_dat_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_47_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] _169_/X vssd vssd vccd vccd _153_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_25_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput954 output954/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_45_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1707 wire1707/A vssd vssd vccd vccd _562_/A sky130_fd_sc_hd__buf_6
XTAP_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1718 wire1718/A vssd vssd vccd vccd _532_/A sky130_fd_sc_hd__buf_6
XTAP_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3380 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1729 wire1729/A vssd vssd vccd vccd _615_/A sky130_fd_sc_hd__buf_6
XTAP_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input263_A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2180_A wire2181/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2278_A wire2278/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input430_A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__296__A _296_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_605_ _605_/A _605_/B vssd vssd vccd vccd _605_/X sky130_fd_sc_hd__and2_4
XFILLER_45_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_536_ _536_/A _536_/B vssd vssd vccd vccd _536_/X sky130_fd_sc_hd__and2_4
XFILLER_15_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_467_ _595_/A _467_/B _467_/C vssd vssd vccd vccd _467_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_398_ _526_/A _398_/B _398_/C vssd vssd vccd vccd _398_/X sky130_fd_sc_hd__and3b_2
XANTENNA_output482_A _486_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1009_A wire1010/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output747_A _622_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1280_A _383_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output914_A wire1367/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire998_A wire999/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__372__C _372_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput740 _616_/X vssd vssd vccd vccd la_oenb_core[119] sky130_fd_sc_hd__buf_8
XFILLER_5_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput751 wire1187/X vssd vssd vccd vccd la_oenb_core[13] sky130_fd_sc_hd__buf_8
XFILLER_47_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput762 wire1177/X vssd vssd vccd vccd la_oenb_core[23] sky130_fd_sc_hd__buf_8
XFILLER_25_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput773 wire1172/X vssd vssd vccd vccd la_oenb_core[33] sky130_fd_sc_hd__buf_8
XFILLER_9_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput784 _540_/X vssd vssd vccd vccd la_oenb_core[43] sky130_fd_sc_hd__buf_8
XFILLER_40_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2205 wire2205/A vssd vssd vccd vccd wire2205/X sky130_fd_sc_hd__buf_6
Xoutput795 wire1156/X vssd vssd vccd vccd la_oenb_core[53] sky130_fd_sc_hd__buf_8
Xwire2216 wire2217/X vssd vssd vccd vccd wire2216/X sky130_fd_sc_hd__buf_6
Xwire2227 wire2227/A vssd vssd vccd vccd wire2227/X sky130_fd_sc_hd__buf_6
XFILLER_43_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2238 wire2238/A vssd vssd vccd vccd wire2238/X sky130_fd_sc_hd__buf_6
Xwire1504 wire1504/A vssd vssd vccd vccd wire1504/X sky130_fd_sc_hd__buf_6
Xwire2249 wire2249/A vssd vssd vccd vccd _460_/B sky130_fd_sc_hd__buf_6
Xwire1515 wire1515/A vssd vssd vccd vccd _366_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1526 wire1527/X vssd vssd vccd vccd wire1526/X sky130_fd_sc_hd__buf_6
XTAP_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1537 wire1537/A vssd vssd vccd vccd wire1537/X sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[7\]_B _170_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1548 wire1548/A vssd vssd vccd vccd wire1548/X sky130_fd_sc_hd__buf_6
Xwire1559 wire1559/A vssd vssd vccd vccd wire1559/X sky130_fd_sc_hd__buf_6
XFILLER_41_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2026_A wire2027/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input109_A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ _321_/A _321_/B vssd vssd vccd vccd _321_/X sky130_fd_sc_hd__and2_2
XTAP_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_252_ _252_/A _252_/B vssd vssd vccd vccd _252_/X sky130_fd_sc_hd__and2_4
XANTENNA__563__B _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3711 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_402 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_183_ _183_/A _183_/B vssd vssd vccd vccd _183_/X sky130_fd_sc_hd__and2_2
XANTENNA_input380_A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input74_A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__457__C _457_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3644 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_519_ _519_/A _519_/B vssd vssd vccd vccd _519_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__473__B _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output864_A _329_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1495_A wire1496/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1662_A wire1662/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] _281_/X vssd vssd vccd vccd _101_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_3_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__383__B _383_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput570 _450_/X vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__buf_8
XFILLER_44_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput581 wire1222/X vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__buf_8
XFILLER_47_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2002 wire2003/X vssd vssd vccd vccd wire2002/X sky130_fd_sc_hd__buf_6
XFILLER_40_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput592 _083_/Y vssd vssd vccd vccd la_data_in_mprj[100] sky130_fd_sc_hd__buf_8
XFILLER_5_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2013 wire2014/X vssd vssd vccd vccd _617_/B sky130_fd_sc_hd__buf_6
Xwire2024 wire2025/X vssd vssd vccd vccd wire2024/X sky130_fd_sc_hd__buf_6
XFILLER_43_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2035 wire2036/X vssd vssd vccd vccd _610_/B sky130_fd_sc_hd__buf_6
Xwire1301 wire1302/X vssd vssd vccd vccd wire1301/X sky130_fd_sc_hd__buf_6
XFILLER_8_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2046 wire2046/A vssd vssd vccd vccd wire2046/X sky130_fd_sc_hd__buf_6
XFILLER_21_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1312 wire1313/X vssd vssd vccd vccd wire1312/X sky130_fd_sc_hd__buf_6
XFILLER_25_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2057 wire2057/A vssd vssd vccd vccd wire2057/X sky130_fd_sc_hd__buf_6
XFILLER_21_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1323 wire1324/X vssd vssd vccd vccd wire1323/X sky130_fd_sc_hd__buf_8
Xwire2068 wire2069/X vssd vssd vccd vccd _595_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1334 wire1335/X vssd vssd vccd vccd wire1334/X sky130_fd_sc_hd__buf_6
XFILLER_43_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2079 wire2079/A vssd vssd vccd vccd wire2079/X sky130_fd_sc_hd__buf_6
XFILLER_8_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1345 _355_/X vssd vssd vccd vccd wire1345/X sky130_fd_sc_hd__buf_6
Xwire1356 wire1357/X vssd vssd vccd vccd wire1356/X sky130_fd_sc_hd__buf_6
XANTENNA__558__B _558_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1367 wire1368/X vssd vssd vccd vccd wire1367/X sky130_fd_sc_hd__buf_6
XFILLER_38_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input226_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2143_A wire2143/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1378 _344_/X vssd vssd vccd vccd wire1378/X sky130_fd_sc_hd__buf_6
Xwire1389 wire1390/X vssd vssd vccd vccd wire1389/X sky130_fd_sc_hd__buf_6
XFILLER_34_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__574__A _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_51_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_304_ _304_/A _304_/B vssd vssd vccd vccd _304_/X sky130_fd_sc_hd__and2_4
XANTENNA__293__B _293_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_235_ _235_/A _235_/B vssd vssd vccd vccd _235_/X sky130_fd_sc_hd__and2_4
XFILLER_50_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_166_ _166_/A _166_/B vssd vssd vccd vccd _166_/X sky130_fd_sc_hd__and2_1
XFILLER_49_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_097_ _097_/A vssd vssd vccd vccd _097_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_26_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1076_A wire1077/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__468__B _468_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1243_A _419_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1890 wire1890/A vssd vssd vccd vccd _270_/A sky130_fd_sc_hd__buf_6
XFILLER_37_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_629 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1410_A wire1411/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1508_A wire1508/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_15_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_190 _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1877_A wire1878/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput309 la_oenb_mprj[29] vssd vssd vccd vccd wire1722/A sky130_fd_sc_hd__buf_6
XFILLER_29_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__B _378_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_51_150 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_020_ _020_/A vssd vssd vccd vccd _020_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input176_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2093_A wire2094/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2260_A wire2260/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input343_A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__569__A _569_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input37_A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1120 _114_/Y vssd vssd vccd vccd wire1120/X sky130_fd_sc_hd__buf_6
XFILLER_1_3038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1131 wire1131/A vssd vssd vccd vccd _067_/A sky130_fd_sc_hd__buf_6
XANTENNA__288__B _288_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1142 wire1142/A vssd vssd vccd vccd _103_/A sky130_fd_sc_hd__buf_6
Xwire1153 wire1154/X vssd vssd vccd vccd wire1153/X sky130_fd_sc_hd__buf_6
XFILLER_40_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1164 _542_/X vssd vssd vccd vccd wire1164/X sky130_fd_sc_hd__buf_6
XFILLER_38_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1175 _522_/X vssd vssd vccd vccd wire1175/X sky130_fd_sc_hd__buf_6
Xwire1186 _511_/X vssd vssd vccd vccd wire1186/X sky130_fd_sc_hd__buf_6
XFILLER_1_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1197 _500_/X vssd vssd vccd vccd wire1197/X sky130_fd_sc_hd__buf_6
XFILLER_34_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_218_ _218_/A _218_/B vssd vssd vccd vccd _218_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output562_A _443_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_149_ _149_/A vssd vssd vccd vccd _149_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__C _470_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output827_A _579_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1360_A _350_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] _237_/X vssd vssd vccd vccd _057_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1625_A wire1626/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1994_A wire1994/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire980_A wire981/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2467 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput106 la_data_out_mprj[77] vssd vssd vccd vccd _446_/C sky130_fd_sc_hd__buf_4
XFILLER_6_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4048 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput117 la_data_out_mprj[87] vssd vssd vccd vccd wire1746/A sky130_fd_sc_hd__buf_6
XFILLER_48_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput128 la_data_out_mprj[97] vssd vssd vccd vccd _466_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput139 la_iena_mprj[106] vssd vssd vccd vccd _269_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2106_A wire2106/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1546 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input293_A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__571__B _571_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_90 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_003_ _003_/A vssd vssd vccd vccd _003_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input460_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__299__A _299_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3812 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1039_A wire1040/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__465__C _465_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output777_A _534_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__481__B _481_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output944_A wire1370/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1575_A wire1576/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__002__A _002_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] _263_/X vssd vssd vccd vccd _083_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__375__C _375_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_632 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__391__B _391_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3534 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input139_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2056_A wire2057/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_621_ _621_/A _621_/B vssd vssd vccd vccd _621_/X sky130_fd_sc_hd__and2_4
XFILLER_22_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1742 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_552_ _552_/A _552_/B vssd vssd vccd vccd _552_/X sky130_fd_sc_hd__and2_4
XANTENNA__566__B _566_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2223_A wire2223/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input306_A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_483_ _611_/A _483_/B _483_/C vssd vssd vccd vccd _483_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__582__A _582_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output525_A wire1253/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1156_A wire1157/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__420__A_N _548_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__476__B _476_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1323_A wire1324/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_779 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output894_A wire1011/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] _200_/X vssd vssd vccd vccd _020_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput900 wire982/X vssd vssd vccd vccd mprj_dat_i_core[27] sky130_fd_sc_hd__buf_8
XFILLER_47_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput911 wire1076/X vssd vssd vccd vccd mprj_dat_i_core[8] sky130_fd_sc_hd__buf_8
XFILLER_9_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput922 wire1343/X vssd vssd vccd vccd mprj_dat_o_user[18] sky130_fd_sc_hd__buf_8
Xoutput933 wire1307/X vssd vssd vccd vccd mprj_dat_o_user[28] sky130_fd_sc_hd__buf_8
Xoutput944 wire1370/X vssd vssd vccd vccd mprj_dat_o_user[9] sky130_fd_sc_hd__buf_8
XFILLER_28_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput955 wire1453/X vssd vssd vccd vccd user_clock sky130_fd_sc_hd__buf_8
XFILLER_45_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1708 wire1708/A vssd vssd vccd vccd _561_/A sky130_fd_sc_hd__buf_6
XTAP_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1719 wire1719/A vssd vssd vccd vccd _529_/A sky130_fd_sc_hd__buf_6
XFILLER_45_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__386__B _386_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_B _260_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_823 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2173_A wire2173/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input256_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__443__A_N _571_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input423_A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__577__A _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_604_ _604_/A _604_/B vssd vssd vccd vccd _604_/X sky130_fd_sc_hd__and2_4
XTAP_4298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_535_ _535_/A _535_/B vssd vssd vccd vccd _535_/X sky130_fd_sc_hd__and2_4
XFILLER_33_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[88\]_B wire1471/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_466_ _594_/A _466_/B _466_/C vssd vssd vccd vccd _466_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_397_ _525_/A _397_/B _397_/C vssd vssd vccd vccd _397_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output475_A _479_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output642_A _013_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1273_A _390_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_B _175_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output907_A wire1096/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1440_A wire1441/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1538_A wire1539/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B wire1480/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__466__A_N _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput730 wire1190/X vssd vssd vccd vccd la_oenb_core[10] sky130_fd_sc_hd__buf_8
Xoutput741 wire1189/X vssd vssd vccd vccd la_oenb_core[11] sky130_fd_sc_hd__buf_8
Xoutput752 wire1186/X vssd vssd vccd vccd la_oenb_core[14] sky130_fd_sc_hd__buf_8
XFILLER_47_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput763 wire1176/X vssd vssd vccd vccd la_oenb_core[24] sky130_fd_sc_hd__buf_8
XFILLER_21_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput774 wire1171/X vssd vssd vccd vccd la_oenb_core[34] sky130_fd_sc_hd__buf_8
XFILLER_25_4199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput785 wire1165/X vssd vssd vccd vccd la_oenb_core[44] sky130_fd_sc_hd__buf_8
XFILLER_5_3537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2206 wire2207/X vssd vssd vccd vccd _483_/B sky130_fd_sc_hd__buf_6
Xoutput796 _551_/X vssd vssd vccd vccd la_oenb_core[54] sky130_fd_sc_hd__buf_8
XFILLER_48_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2217 wire2217/A vssd vssd vccd vccd wire2217/X sky130_fd_sc_hd__buf_6
Xwire2228 wire2229/X vssd vssd vccd vccd _474_/B sky130_fd_sc_hd__buf_6
Xwire2239 wire2239/A vssd vssd vccd vccd _468_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1505 wire1506/X vssd vssd vccd vccd _342_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1516 wire1516/A vssd vssd vccd vccd _365_/B sky130_fd_sc_hd__buf_6
Xwire1527 wire1527/A vssd vssd vccd vccd wire1527/X sky130_fd_sc_hd__buf_6
XTAP_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1538 wire1539/X vssd vssd vccd vccd _350_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1549 wire1550/X vssd vssd vccd vccd _298_/B sky130_fd_sc_hd__buf_6
XFILLER_38_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ _320_/A _320_/B vssd vssd vccd vccd _320_/X sky130_fd_sc_hd__and2_4
XFILLER_42_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_251_ _251_/A _251_/B vssd vssd vccd vccd _251_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_182_ _182_/A _182_/B vssd vssd vccd vccd _182_/X sky130_fd_sc_hd__and2_2
XFILLER_49_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input373_A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input67_A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__100__A _100_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_518_ _518_/A _518_/B vssd vssd vccd vccd _518_/X sky130_fd_sc_hd__and2_4
XTAP_2682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1021_A wire1022/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output592_A _083_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1119_A wire1120/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__473__C _473_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_449_ _577_/A _449_/B _449_/C vssd vssd vccd vccd _449_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__489__A_N _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output857_A wire1403/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1655_A wire1656/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1822_A wire1823/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__383__C _383_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput560 _441_/X vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__buf_8
XFILLER_40_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput571 _451_/X vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__buf_8
XFILLER_43_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput582 wire1221/X vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__buf_8
XFILLER_44_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2003 wire2003/A vssd vssd vccd vccd wire2003/X sky130_fd_sc_hd__buf_6
Xoutput593 _084_/Y vssd vssd vccd vccd la_data_in_mprj[101] sky130_fd_sc_hd__buf_8
XFILLER_8_1011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2014 wire2015/X vssd vssd vccd vccd wire2014/X sky130_fd_sc_hd__buf_6
XFILLER_40_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2025 wire2025/A vssd vssd vccd vccd wire2025/X sky130_fd_sc_hd__buf_6
Xwire2036 wire2037/X vssd vssd vccd vccd wire2036/X sky130_fd_sc_hd__buf_6
XFILLER_43_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2047 wire2048/X vssd vssd vccd vccd _605_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1302 _367_/X vssd vssd vccd vccd wire1302/X sky130_fd_sc_hd__buf_6
Xwire2058 wire2059/X vssd vssd vccd vccd _600_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1055 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1313 wire1314/X vssd vssd vccd vccd wire1313/X sky130_fd_sc_hd__buf_6
Xwire1324 wire1325/X vssd vssd vccd vccd wire1324/X sky130_fd_sc_hd__buf_6
Xwire2069 wire2069/A vssd vssd vccd vccd wire2069/X sky130_fd_sc_hd__buf_6
XFILLER_25_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1335 wire1336/X vssd vssd vccd vccd wire1335/X sky130_fd_sc_hd__buf_6
Xwire1346 wire1347/X vssd vssd vccd vccd wire1346/X sky130_fd_sc_hd__buf_6
XFILLER_1_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1357 _351_/X vssd vssd vccd vccd wire1357/X sky130_fd_sc_hd__buf_6
Xwire1368 wire1369/X vssd vssd vccd vccd wire1368/X sky130_fd_sc_hd__buf_6
Xwire1379 wire1380/X vssd vssd vccd vccd wire1379/X sky130_fd_sc_hd__buf_6
XFILLER_28_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input121_A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input219_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__574__B _574_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2303_A wire2304/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_303_ _303_/A _303_/B vssd vssd vccd vccd _303_/X sky130_fd_sc_hd__and2_2
XTAP_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_234_ _234_/A _234_/B vssd vssd vccd vccd _234_/X sky130_fd_sc_hd__and2_4
XFILLER_7_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__590__A _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_165_ _165_/A _165_/B vssd vssd vccd vccd _165_/X sky130_fd_sc_hd__and2_1
XFILLER_6_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] max_cap1456/X vssd vssd vccd vccd _116_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_096_ _096_/A vssd vssd vccd vccd _096_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_powergood_check_mprj_vdd_logic1 output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1069_A wire1070/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__468__C _468_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1880 wire1880/A vssd vssd vccd vccd wire1880/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1236_A wire1237/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1891 wire1892/X vssd vssd vccd vccd _269_/A sky130_fd_sc_hd__buf_6
XFILLER_0_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__484__B _484_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_B _281_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_180 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_191 _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1772_A wire1773/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4158 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[27\]_A mprj_dat_i_user[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__C _378_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3206 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__B _394_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[109\]_B _272_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2086_A wire2086/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input169_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__569__B _569_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2253_A wire2254/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input336_A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[18\]_A mprj_dat_i_user[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1110 _116_/Y vssd vssd vccd vccd wire1110/X sky130_fd_sc_hd__buf_6
Xwire1121 wire1121/A vssd vssd vccd vccd _082_/A sky130_fd_sc_hd__buf_6
Xwire1132 wire1132/A vssd vssd vccd vccd _066_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1143 _624_/X vssd vssd vccd vccd wire1143/X sky130_fd_sc_hd__buf_6
Xwire1154 _553_/X vssd vssd vccd vccd wire1154/X sky130_fd_sc_hd__buf_6
XFILLER_43_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1165 _541_/X vssd vssd vccd vccd wire1165/X sky130_fd_sc_hd__buf_6
Xwire1176 _521_/X vssd vssd vccd vccd wire1176/X sky130_fd_sc_hd__buf_6
XFILLER_19_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1187 _510_/X vssd vssd vccd vccd wire1187/X sky130_fd_sc_hd__buf_6
XFILLER_5_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1198 _499_/X vssd vssd vccd vccd wire1198/X sky130_fd_sc_hd__buf_6
XFILLER_53_3907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__585__A _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_217_ _217_/A _217_/B vssd vssd vccd vccd _217_/X sky130_fd_sc_hd__and2_2
XFILLER_51_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_148_ _148_/A vssd vssd vccd vccd _148_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_079_ _079_/A vssd vssd vccd vccd _079_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wire1186_A _511_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output722_A _599_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__479__B _479_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1353_A wire1354/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] _230_/X vssd vssd vccd vccd _050_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1520_A wire1520/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1618_A wire1619/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_170 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3439 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1987_A wire1987/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire973_A _144_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3519 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput107 la_data_out_mprj[78] vssd vssd vccd vccd _447_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput118 la_data_out_mprj[88] vssd vssd vccd vccd wire1745/A sky130_fd_sc_hd__buf_6
XANTENNA__389__B _389_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput129 la_data_out_mprj[98] vssd vssd vccd vccd _467_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3050 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2001_A wire2002/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input286_A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_80 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_002_ _002_/A vssd vssd vccd vccd _002_/Y sky130_fd_sc_hd__inv_2
XANTENNA_91 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input453_A mprj_iena_wb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__299__B _299_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1101_A wire1102/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__481__C _481_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output937_A wire1295/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1470_A _252_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1568_A wire1569/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__391__C _391_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_620_ _620_/A _620_/B vssd vssd vccd vccd _620_/X sky130_fd_sc_hd__and2_4
XTAP_4458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2049_A wire2049/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_551_ _551_/A _551_/B vssd vssd vccd vccd _551_/X sky130_fd_sc_hd__and2_4
XTAP_3768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input201_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_482_ _610_/A _482_/B _482_/C vssd vssd vccd vccd _482_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2216_A wire2217/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__372__A_N _500_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__582__B _582_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input97_A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__103__A _103_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output518_A wire1259/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput460 user_irq_ena[0] vssd vssd vccd vccd _291_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1051_A wire1052/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1149_A _557_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_202 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__476__C _476_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1316_A wire1317/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output887_A wire1041/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__492__B _492_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1685_A wire1685/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput901 wire978/X vssd vssd vccd vccd mprj_dat_i_core[28] sky130_fd_sc_hd__buf_8
Xoutput912 wire1071/X vssd vssd vccd vccd mprj_dat_i_core[9] sky130_fd_sc_hd__buf_8
XANTENNA_wire1852_A wire1852/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput923 wire1340/X vssd vssd vccd vccd mprj_dat_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_9_3844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput934 wire1303/X vssd vssd vccd vccd mprj_dat_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_47_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput945 wire1440/X vssd vssd vccd vccd mprj_sel_o_user[0] sky130_fd_sc_hd__buf_8
Xoutput956 _297_/X vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__buf_8
XFILLER_9_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__013__A _013_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1709 wire1709/A vssd vssd vccd vccd _560_/A sky130_fd_sc_hd__buf_6
XTAP_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__395__A_N _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input151_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2166_A wire2166/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input249_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__577__B _577_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input416_A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_603_ _603_/A _603_/B vssd vssd vccd vccd _603_/X sky130_fd_sc_hd__and2_4
XTAP_4288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_534_ _534_/A _534_/B vssd vssd vccd vccd _534_/X sky130_fd_sc_hd__and2_4
XTAP_2842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__593__A _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ _593_/A _465_/B _465_/C vssd vssd vccd vccd _465_/X sky130_fd_sc_hd__and3b_1
XTAP_2897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_396_ _524_/A _396_/B _396_/C vssd vssd vccd vccd _396_/X sky130_fd_sc_hd__and3b_4
XFILLER_9_423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xmax_cap1456 split4/A vssd vssd vccd vccd max_cap1456/X sky130_fd_sc_hd__buf_8
XFILLER_9_3107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output468_A wire1211/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1099_A wire1100/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3923 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1266_A _396_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output802_A wire1195/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__487__B _487_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1433_A wire1434/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput290 la_oenb_mprj[127] vssd vssd vccd vccd _624_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1600_A wire1601/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput720 _597_/X vssd vssd vccd vccd la_oenb_core[100] sky130_fd_sc_hd__buf_8
XFILLER_47_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput731 _607_/X vssd vssd vccd vccd la_oenb_core[110] sky130_fd_sc_hd__buf_8
XFILLER_9_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput742 _617_/X vssd vssd vccd vccd la_oenb_core[120] sky130_fd_sc_hd__buf_8
Xoutput753 wire1185/X vssd vssd vccd vccd la_oenb_core[15] sky130_fd_sc_hd__buf_8
XFILLER_25_3433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput764 wire1175/X vssd vssd vccd vccd la_oenb_core[25] sky130_fd_sc_hd__buf_8
XFILLER_47_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput775 _532_/X vssd vssd vccd vccd la_oenb_core[35] sky130_fd_sc_hd__buf_8
XFILLER_5_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput786 wire1164/X vssd vssd vccd vccd la_oenb_core[45] sky130_fd_sc_hd__buf_8
Xwire2207 wire2208/X vssd vssd vccd vccd wire2207/X sky130_fd_sc_hd__buf_6
Xoutput797 wire1155/X vssd vssd vccd vccd la_oenb_core[55] sky130_fd_sc_hd__buf_8
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2218 wire2219/X vssd vssd vccd vccd _479_/B sky130_fd_sc_hd__buf_6
Xwire2229 wire2229/A vssd vssd vccd vccd wire2229/X sky130_fd_sc_hd__buf_6
XFILLER_5_2837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1506 wire1506/A vssd vssd vccd vccd wire1506/X sky130_fd_sc_hd__buf_6
XFILLER_3_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1517 wire1517/A vssd vssd vccd vccd _364_/B sky130_fd_sc_hd__buf_6
XFILLER_47_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1528 wire1528/A vssd vssd vccd vccd _356_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1539 wire1539/A vssd vssd vccd vccd wire1539/X sky130_fd_sc_hd__buf_6
XANTENNA__397__B _397_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_250_ _250_/A _250_/B vssd vssd vccd vccd _250_/X sky130_fd_sc_hd__and2_4
XFILLER_36_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_181_ _181_/A _181_/B vssd vssd vccd vccd _181_/X sky130_fd_sc_hd__and2_4
XFILLER_52_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input199_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__A_N _538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input366_A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2283_A wire2283/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_irq_gates\[1\] user_irq_core[1] _292_/X vssd vssd vccd vccd _112_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__588__A _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_517_ _517_/A _517_/B vssd vssd vccd vccd _517_/X sky130_fd_sc_hd__and2_4
XTAP_2672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1334 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ _576_/A _448_/B _448_/C vssd vssd vccd vccd _448_/X sky130_fd_sc_hd__and3b_4
XTAP_1982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1014_A wire1015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output585_A wire1218/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_379_ _507_/A _379_/B _379_/C vssd vssd vccd vccd _379_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output752_A wire1186/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1383_A wire1384/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] _260_/X vssd vssd vccd vccd wire1123/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_42_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1550_A wire1551/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1648_A wire1649/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__498__A _498_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1579 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1815_A wire1815/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__433__A_N _561_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput550 _432_/X vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__buf_8
Xoutput561 _442_/X vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__buf_8
Xoutput572 _452_/X vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__buf_8
XFILLER_5_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput583 wire1220/X vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__buf_8
Xwire2004 wire2005/X vssd vssd vccd vccd _620_/B sky130_fd_sc_hd__buf_6
Xoutput594 _085_/Y vssd vssd vccd vccd la_data_in_mprj[102] sky130_fd_sc_hd__buf_8
XFILLER_5_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2015 wire2015/A vssd vssd vccd vccd wire2015/X sky130_fd_sc_hd__buf_6
XFILLER_8_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2026 wire2027/X vssd vssd vccd vccd _613_/B sky130_fd_sc_hd__buf_6
Xwire2037 wire2037/A vssd vssd vccd vccd wire2037/X sky130_fd_sc_hd__buf_6
Xwire1303 wire1304/X vssd vssd vccd vccd wire1303/X sky130_fd_sc_hd__buf_8
XFILLER_5_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2048 wire2049/X vssd vssd vccd vccd wire2048/X sky130_fd_sc_hd__buf_6
XFILLER_43_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2059 wire2059/A vssd vssd vccd vccd wire2059/X sky130_fd_sc_hd__buf_6
XANTENNA__201__A _201_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1314 _364_/X vssd vssd vccd vccd wire1314/X sky130_fd_sc_hd__buf_6
Xwire1325 wire1326/X vssd vssd vccd vccd wire1325/X sky130_fd_sc_hd__buf_6
XFILLER_47_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1336 _358_/X vssd vssd vccd vccd wire1336/X sky130_fd_sc_hd__buf_6
Xwire1347 wire1348/X vssd vssd vccd vccd wire1347/X sky130_fd_sc_hd__buf_6
XFILLER_3_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1358 wire1359/X vssd vssd vccd vccd wire1358/X sky130_fd_sc_hd__buf_6
XFILLER_5_1955 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1369 _347_/X vssd vssd vccd vccd wire1369/X sky130_fd_sc_hd__buf_6
XFILLER_38_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2031_A wire2031/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input114_A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2129_A wire2129/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _302_/A _302_/B vssd vssd vccd vccd _302_/X sky130_fd_sc_hd__and2_4
XFILLER_51_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_233_ _233_/A _233_/B vssd vssd vccd vccd _233_/X sky130_fd_sc_hd__and2_2
XFILLER_50_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__590__B _590_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_164_ _164_/A _164_/B vssd vssd vccd vccd _164_/X sky130_fd_sc_hd__and2_1
XFILLER_7_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_095_ _095_/A vssd vssd vccd vccd _095_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1898 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1870 wire1871/X vssd vssd vccd vccd _283_/A sky130_fd_sc_hd__buf_6
XANTENNA_output500_A wire1276/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1881 wire1882/X vssd vssd vccd vccd _278_/A sky130_fd_sc_hd__buf_6
XFILLER_37_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1892 wire1892/A vssd vssd vccd vccd wire1892/X sky130_fd_sc_hd__buf_6
XFILLER_34_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1131_A wire1131/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1229_A wire1230/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__456__A_N _584_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__484__C _484_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_170 wire2304/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_181 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_192 _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] _175_/X vssd vssd vccd vccd _159_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] split5/A vssd vssd vccd vccd _139_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_50_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1598_A wire1599/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1765_A wire1765/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[27\]_B split5/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] _286_/X vssd vssd vccd vccd wire1139/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_29_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__394__C _394_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_rebuffer2_A split4/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2079_A wire2079/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1100 _118_/Y vssd vssd vccd vccd wire1100/X sky130_fd_sc_hd__buf_6
XANTENNA_user_wb_dat_gates\[18\]_B load_slew1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1111 wire1112/X vssd vssd vccd vccd wire1111/X sky130_fd_sc_hd__buf_6
Xwire1122 wire1122/A vssd vssd vccd vccd _081_/A sky130_fd_sc_hd__buf_6
XFILLER_43_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input231_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1133 wire1133/A vssd vssd vccd vccd _065_/A sky130_fd_sc_hd__buf_6
XANTENNA_wire2246_A wire2246/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input329_A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__479__A_N _607_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1144 _623_/X vssd vssd vccd vccd wire1144/X sky130_fd_sc_hd__buf_6
Xwire1155 _552_/X vssd vssd vccd vccd wire1155/X sky130_fd_sc_hd__buf_6
XFILLER_47_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1166 _539_/X vssd vssd vccd vccd wire1166/X sky130_fd_sc_hd__buf_6
Xwire1177 _520_/X vssd vssd vccd vccd wire1177/X sky130_fd_sc_hd__buf_6
XFILLER_5_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1188 _509_/X vssd vssd vccd vccd wire1188/X sky130_fd_sc_hd__buf_6
Xwire1199 _498_/X vssd vssd vccd vccd wire1199/X sky130_fd_sc_hd__buf_6
XFILLER_38_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__585__B _585_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3064 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_216_ _216_/A _216_/B vssd vssd vccd vccd _216_/X sky130_fd_sc_hd__and2_2
XFILLER_11_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__106__A _106_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_147_ _147_/A vssd vssd vccd vccd _147_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1083 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_078_ _078_/A vssd vssd vccd vccd _078_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output548_A wire1226/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1081_A wire1082/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3734 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1179_A _518_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__479__C _479_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output715_A _080_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1346_A wire1347/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__495__B _495_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1513_A wire1514/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_182 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire966_A wire967/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__016__A _016_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1746 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2988 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput108 la_data_out_mprj[79] vssd vssd vccd vccd _448_/C sky130_fd_sc_hd__buf_4
XFILLER_44_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput119 la_data_out_mprj[89] vssd vssd vccd vccd _458_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2690 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_70 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_001_ _001_/A vssd vssd vccd vccd _001_/Y sky130_fd_sc_hd__inv_2
XANTENNA_81 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_92 _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input181_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input279_A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2196_A wire2196/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input446_A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input42_A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1858 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__596__A _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output498_A wire1278/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1296_A wire1297/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output832_A _584_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1630_A wire1631/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput90 la_data_out_mprj[62] vssd vssd vccd vccd _431_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_550_ _550_/A _550_/B vssd vssd vccd vccd _550_/X sky130_fd_sc_hd__and2_2
XTAP_3758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_481_ _609_/A _481_/B _481_/C vssd vssd vccd vccd _481_/X sky130_fd_sc_hd__and3b_4
XFILLER_2_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2111_A wire2112/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3700 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2209_A wire2210/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input396_A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput450 mprj_dat_o_core[7] vssd vssd vccd vccd wire1502/A sky130_fd_sc_hd__buf_6
XFILLER_23_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput461 user_irq_ena[1] vssd vssd vccd vccd _292_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1044_A wire1045/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output782_A wire1167/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1309_A wire1310/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__492__C _492_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1580_A wire1581/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1678_A wire1679/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput902 wire974/X vssd vssd vccd vccd mprj_dat_i_core[29] sky130_fd_sc_hd__buf_8
XFILLER_29_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput913 wire1395/X vssd vssd vccd vccd mprj_dat_o_user[0] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput924 wire1393/X vssd vssd vccd vccd mprj_dat_o_user[1] sky130_fd_sc_hd__buf_8
Xoutput935 wire1391/X vssd vssd vccd vccd mprj_dat_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_25_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput946 wire1435/X vssd vssd vccd vccd mprj_sel_o_user[1] sky130_fd_sc_hd__buf_8
XFILLER_8_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput957 _111_/Y vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__buf_8
XANTENNA_wire1845_A wire1846/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__204__A _204_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1870 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input144_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2061_A wire2061/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2159_A wire2159/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_602_ _602_/A _602_/B vssd vssd vccd vccd _602_/X sky130_fd_sc_hd__and2_4
XTAP_4278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input311_A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input409_A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_533_ _533_/A _533_/B vssd vssd vccd vccd _533_/X sky130_fd_sc_hd__and2_4
XTAP_2843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__593__B _593_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_464_ _592_/A _464_/B _464_/C vssd vssd vccd vccd _464_/X sky130_fd_sc_hd__and3b_4
XTAP_2898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_395_ _523_/A _395_/B _395_/C vssd vssd vccd vccd _395_/X sky130_fd_sc_hd__and3b_2
XFILLER_35_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output530_A wire1248/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output628_A _001_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1161_A _547_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1259_A _403_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__487__C _487_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput280 la_oenb_mprj[118] vssd vssd vccd vccd wire1729/A sky130_fd_sc_hd__buf_6
XFILLER_23_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput291 la_oenb_mprj[12] vssd vssd vccd vccd _509_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1426_A wire1427/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] _205_/X vssd vssd vccd vccd _025_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_4055 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1962_A wire1962/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput710 _075_/Y vssd vssd vccd vccd la_data_in_mprj[92] sky130_fd_sc_hd__buf_8
Xoutput721 _598_/X vssd vssd vccd vccd la_oenb_core[101] sky130_fd_sc_hd__buf_8
XANTENNA__024__A _024_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput732 _608_/X vssd vssd vccd vccd la_oenb_core[111] sky130_fd_sc_hd__buf_8
XFILLER_47_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput743 _618_/X vssd vssd vccd vccd la_oenb_core[121] sky130_fd_sc_hd__buf_8
XFILLER_9_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput754 wire1184/X vssd vssd vccd vccd la_oenb_core[16] sky130_fd_sc_hd__buf_8
Xoutput765 wire1174/X vssd vssd vccd vccd la_oenb_core[26] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] _167_/X vssd vssd vccd vccd _151_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_9_3686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput776 _533_/X vssd vssd vccd vccd la_oenb_core[36] sky130_fd_sc_hd__buf_8
XFILLER_28_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput787 _543_/X vssd vssd vccd vccd la_oenb_core[46] sky130_fd_sc_hd__buf_8
Xwire2208 wire2208/A vssd vssd vccd vccd wire2208/X sky130_fd_sc_hd__buf_6
Xoutput798 wire1153/X vssd vssd vccd vccd la_oenb_core[56] sky130_fd_sc_hd__buf_8
Xwire2219 wire2219/A vssd vssd vccd vccd wire2219/X sky130_fd_sc_hd__buf_6
XFILLER_25_2755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1507 wire1508/X vssd vssd vccd vccd _341_/B sky130_fd_sc_hd__buf_6
XTAP_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1518 wire1518/A vssd vssd vccd vccd _363_/B sky130_fd_sc_hd__buf_6
XFILLER_38_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1529 wire1529/A vssd vssd vccd vccd _355_/B sky130_fd_sc_hd__buf_6
XTAP_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__397__C _397_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_180_ _180_/A _180_/B vssd vssd vccd vccd _180_/X sky130_fd_sc_hd__and2_2
XFILLER_17_2294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input261_A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2276_A wire2276/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input359_A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__588__B _588_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_516_ _516_/A _516_/B vssd vssd vccd vccd _516_/X sky130_fd_sc_hd__and2_4
XTAP_2673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__109__A _109_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_447_ _447_/A_N _447_/B _447_/C vssd vssd vccd vccd _447_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1346 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3360 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1007_A wire1008/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_378_ _506_/A _378_/B _378_/C vssd vssd vccd vccd _378_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output480_A _484_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output578_A wire1224/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output745_A _620_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__385__A_N _513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1376_A wire1377/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output912_A wire1071/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__498__B _498_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1808_A wire1809/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput540 wire1236/X vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__buf_8
XFILLER_25_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput551 _433_/X vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__buf_8
XFILLER_9_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput562 _443_/X vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__buf_8
Xoutput573 _453_/X vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__buf_8
XFILLER_43_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput584 wire1219/X vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__buf_8
Xwire2005 wire2006/X vssd vssd vccd vccd wire2005/X sky130_fd_sc_hd__buf_6
Xoutput595 _086_/Y vssd vssd vccd vccd la_data_in_mprj[103] sky130_fd_sc_hd__buf_8
XFILLER_21_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2016 wire2017/X vssd vssd vccd vccd _616_/B sky130_fd_sc_hd__buf_6
Xwire2027 wire2028/X vssd vssd vccd vccd wire2027/X sky130_fd_sc_hd__buf_6
Xwire2038 wire2039/X vssd vssd vccd vccd _609_/B sky130_fd_sc_hd__buf_6
Xwire1304 wire1305/X vssd vssd vccd vccd wire1304/X sky130_fd_sc_hd__buf_6
Xwire2049 wire2049/A vssd vssd vccd vccd wire2049/X sky130_fd_sc_hd__buf_6
Xwire1315 wire1316/X vssd vssd vccd vccd wire1315/X sky130_fd_sc_hd__buf_8
XFILLER_5_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1326 _361_/X vssd vssd vccd vccd wire1326/X sky130_fd_sc_hd__buf_6
Xwire1337 wire1338/X vssd vssd vccd vccd wire1337/X sky130_fd_sc_hd__buf_6
XFILLER_19_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1348 _354_/X vssd vssd vccd vccd wire1348/X sky130_fd_sc_hd__buf_6
Xwire1359 wire1360/X vssd vssd vccd vccd wire1359/X sky130_fd_sc_hd__buf_6
XFILLER_5_1967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2024_A wire2025/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input107_A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_301_ _301_/A _301_/B vssd vssd vccd vccd _301_/X sky130_fd_sc_hd__and2_4
XTAP_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_232_ _232_/A _232_/B vssd vssd vccd vccd _232_/X sky130_fd_sc_hd__and2_2
XFILLER_24_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_163_ _163_/A vssd vssd vccd vccd _163_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input72_A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_094_ _094_/A vssd vssd vccd vccd _094_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__599__A _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1860 wire1860/A vssd vssd vccd vccd wire1860/X sky130_fd_sc_hd__buf_6
Xwire1871 wire1872/X vssd vssd vccd vccd wire1871/X sky130_fd_sc_hd__buf_6
XFILLER_20_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1882 wire1882/A vssd vssd vccd vccd wire1882/X sky130_fd_sc_hd__buf_6
XFILLER_4_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1893 wire1894/X vssd vssd vccd vccd _268_/A sky130_fd_sc_hd__buf_6
XTAP_3160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_171 _398_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_182 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output862_A wire1398/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] load_slew1458/X vssd vssd vccd vccd _132_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_31_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1660_A wire1661/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1758_A wire1758/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__302__A _302_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] _279_/X vssd vssd vccd vccd _099_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__400__A_N _400_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_378 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3842 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__212__A _212_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1101 wire1102/X vssd vssd vccd vccd wire1101/X sky130_fd_sc_hd__buf_8
XFILLER_0_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1112 wire1113/X vssd vssd vccd vccd wire1112/X sky130_fd_sc_hd__buf_8
XFILLER_5_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1123 wire1123/A vssd vssd vccd vccd _080_/A sky130_fd_sc_hd__buf_6
XFILLER_5_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1134 wire1134/A vssd vssd vccd vccd _064_/A sky130_fd_sc_hd__buf_6
XFILLER_43_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1145 _588_/X vssd vssd vccd vccd wire1145/X sky130_fd_sc_hd__buf_6
Xwire1156 wire1157/X vssd vssd vccd vccd wire1156/X sky130_fd_sc_hd__buf_6
Xwire1167 wire1168/X vssd vssd vccd vccd wire1167/X sky130_fd_sc_hd__buf_6
XANTENNA_input224_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2141_A wire2141/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1178 _519_/X vssd vssd vccd vccd wire1178/X sky130_fd_sc_hd__buf_6
XFILLER_1_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2239_A wire2239/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1189 _508_/X vssd vssd vccd vccd wire1189/X sky130_fd_sc_hd__buf_6
XFILLER_28_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3076 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_215_ _215_/A _215_/B vssd vssd vccd vccd _215_/X sky130_fd_sc_hd__and2_2
XFILLER_32_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_146_ _146_/A vssd vssd vccd vccd _146_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_3396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_077_ _077_/A vssd vssd vccd vccd _077_/Y sky130_fd_sc_hd__inv_4
XFILLER_45_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1074_A wire1075/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__423__A_N _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output610_A _100_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output708_A _073_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1339_A _357_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1690 wire1690/A vssd vssd vccd vccd _579_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3506 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1506_A wire1506/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1875_A wire1876/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__032__A _032_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput109 la_data_out_mprj[7] vssd vssd vccd vccd _376_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_6_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2206 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__207__A _207_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_60 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_000_ _000_/A vssd vssd vccd vccd _000_/Y sky130_fd_sc_hd__inv_2
XANTENNA_71 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_82 _269_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_93 _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2091_A wire2091/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input174_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2189_A wire2190/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__446__A_N _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3178 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input341_A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1815 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input439_A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input35_A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__596__B _596_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__117__A _117_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output560_A _441_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output658_A _028_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_129_ _129_/A vssd vssd vccd vccd _129_/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_wire1191_A _506_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[42\]_B _205_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1289_A _374_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output825_A _577_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3554 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] _235_/X vssd vssd vccd vccd _055_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1623_A wire1624/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4059 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1992_A wire1993/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__027__A _027_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__469__A_N _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput80 la_data_out_mprj[53] vssd vssd vccd vccd _422_/C sky130_fd_sc_hd__buf_4
Xinput91 la_data_out_mprj[63] vssd vssd vccd vccd input91/X sky130_fd_sc_hd__buf_6
XFILLER_43_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[33\]_B _196_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1618 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_480_ _608_/A _480_/B _480_/C vssd vssd vccd vccd _480_/X sky130_fd_sc_hd__and3b_4
XFILLER_17_4560 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2104_A wire2104/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1302 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input291_A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input389_A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3924 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput440 mprj_dat_o_core[27] vssd vssd vccd vccd wire1517/A sky130_fd_sc_hd__buf_6
Xinput451 mprj_dat_o_core[8] vssd vssd vccd vccd wire1500/A sky130_fd_sc_hd__buf_6
Xinput462 user_irq_ena[2] vssd vssd vccd vccd _293_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1037_A wire1038/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output775_A _532_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output942_A wire1376/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1573_A wire1574/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput903 wire1106/X vssd vssd vccd vccd mprj_dat_i_core[2] sky130_fd_sc_hd__buf_8
Xoutput914 wire1367/X vssd vssd vccd vccd mprj_dat_o_user[10] sky130_fd_sc_hd__buf_8
Xoutput925 wire1337/X vssd vssd vccd vccd mprj_dat_o_user[20] sky130_fd_sc_hd__buf_8
XFILLER_47_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput936 wire1299/X vssd vssd vccd vccd mprj_dat_o_user[30] sky130_fd_sc_hd__buf_8
XFILLER_9_3857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput947 wire1430/X vssd vssd vccd vccd mprj_sel_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_9_3868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput958 _112_/Y vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__buf_8
XFILLER_23_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1838_A wire1839/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__310__A _310_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2054_A wire2055/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input137_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_601_ _601_/A _601_/B vssd vssd vccd vccd _601_/X sky130_fd_sc_hd__and2_4
XTAP_4268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_532_ _532_/A _532_/B vssd vssd vccd vccd _532_/X sky130_fd_sc_hd__and2_4
XTAP_2822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2221_A wire2221/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input304_A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_463_ _591_/A _463_/B _463_/C vssd vssd vccd vccd _463_/X sky130_fd_sc_hd__and3b_4
XTAP_2877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_394_ _522_/A _394_/B _394_/C vssd vssd vccd vccd _394_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4298 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output523_A wire1254/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput270 la_oenb_mprj[109] vssd vssd vccd vccd _606_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_49_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput281 la_oenb_mprj[119] vssd vssd vccd vccd wire1728/A sky130_fd_sc_hd__buf_6
XFILLER_7_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput292 la_oenb_mprj[13] vssd vssd vccd vccd _510_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1321_A wire1322/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_568 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output892_A wire1111/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1419_A _315_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] _198_/X vssd vssd vccd vccd _018_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_14_3306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1690_A wire1690/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1788_A wire1789/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__305__A _305_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput700 _066_/Y vssd vssd vccd vccd la_data_in_mprj[83] sky130_fd_sc_hd__buf_8
XFILLER_9_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput711 _076_/Y vssd vssd vccd vccd la_data_in_mprj[93] sky130_fd_sc_hd__buf_8
Xoutput722 _599_/X vssd vssd vccd vccd la_oenb_core[102] sky130_fd_sc_hd__buf_8
Xoutput733 _609_/X vssd vssd vccd vccd la_oenb_core[112] sky130_fd_sc_hd__buf_8
Xoutput744 _619_/X vssd vssd vccd vccd la_oenb_core[122] sky130_fd_sc_hd__buf_8
Xoutput755 wire1183/X vssd vssd vccd vccd la_oenb_core[17] sky130_fd_sc_hd__buf_8
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput766 _524_/X vssd vssd vccd vccd la_oenb_core[27] sky130_fd_sc_hd__buf_8
Xoutput777 _534_/X vssd vssd vccd vccd la_oenb_core[37] sky130_fd_sc_hd__buf_8
XFILLER_5_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput788 _544_/X vssd vssd vccd vccd la_oenb_core[47] sky130_fd_sc_hd__buf_8
Xoutput799 wire1152/X vssd vssd vccd vccd la_oenb_core[57] sky130_fd_sc_hd__buf_8
Xwire2209 wire2210/X vssd vssd vccd vccd _482_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1508 wire1508/A vssd vssd vccd vccd wire1508/X sky130_fd_sc_hd__buf_6
XFILLER_28_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1519 wire1519/A vssd vssd vccd vccd _362_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__215__A _215_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_656 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2171_A wire2172/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input254_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2269_A wire2270/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input421_A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_515_ _515_/A _515_/B vssd vssd vccd vccd _515_/X sky130_fd_sc_hd__and2_4
XTAP_2652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_446_ _574_/A _446_/B _446_/C vssd vssd vccd vccd _446_/X sky130_fd_sc_hd__and3b_4
XTAP_1962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_377_ _505_/A _377_/B _377_/C vssd vssd vccd vccd _377_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output473_A _478_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output640_A _012_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output738_A _614_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3755 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1271_A _392_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1369_A _347_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output905_A wire966/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1536_A wire1537/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1703_A wire1703/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire989_A wire990/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__035__A _035_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput530 wire1248/X vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__buf_8
Xoutput541 wire1234/X vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__buf_8
Xoutput552 _434_/X vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__buf_8
XFILLER_25_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput563 _444_/X vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__buf_8
XFILLER_47_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput574 _454_/X vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__buf_8
Xoutput585 wire1218/X vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__buf_8
Xwire2006 wire2006/A vssd vssd vccd vccd wire2006/X sky130_fd_sc_hd__buf_6
XFILLER_25_2531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput596 _087_/Y vssd vssd vccd vccd la_data_in_mprj[104] sky130_fd_sc_hd__buf_8
Xwire2017 wire2018/X vssd vssd vccd vccd wire2017/X sky130_fd_sc_hd__buf_6
XFILLER_5_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2028 wire2028/A vssd vssd vccd vccd wire2028/X sky130_fd_sc_hd__buf_6
XFILLER_21_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2039 wire2039/A vssd vssd vccd vccd wire2039/X sky130_fd_sc_hd__buf_6
Xwire1305 wire1306/X vssd vssd vccd vccd wire1305/X sky130_fd_sc_hd__buf_6
Xwire1316 wire1317/X vssd vssd vccd vccd wire1316/X sky130_fd_sc_hd__buf_6
Xwire1327 wire1328/X vssd vssd vccd vccd wire1327/X sky130_fd_sc_hd__buf_8
Xwire1338 wire1339/X vssd vssd vccd vccd wire1338/X sky130_fd_sc_hd__buf_6
XFILLER_5_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1349 wire1350/X vssd vssd vccd vccd wire1349/X sky130_fd_sc_hd__buf_6
XFILLER_41_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ _300_/A _300_/B vssd vssd vccd vccd _300_/X sky130_fd_sc_hd__and2_4
XFILLER_42_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2017_A wire2018/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_231_ _231_/A _231_/B vssd vssd vccd vccd _231_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_162_ _162_/A vssd vssd vccd vccd _162_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_3556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_093_ _093_/A vssd vssd vccd vccd _093_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input371_A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input65_A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__599__B _599_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_load_slew1459_A wire1460/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1850 wire1851/X vssd vssd vccd vccd _290_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1861 wire1862/X vssd vssd vccd vccd _286_/A sky130_fd_sc_hd__buf_6
XFILLER_1_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1872 wire1872/A vssd vssd vccd vccd wire1872/X sky130_fd_sc_hd__buf_6
Xwire1883 wire1883/A vssd vssd vccd vccd _277_/A sky130_fd_sc_hd__buf_6
Xwire1894 wire1894/A vssd vssd vccd vccd wire1894/X sky130_fd_sc_hd__buf_6
XTAP_3150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_150 _504_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_161 _474_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 wire1761/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_183 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output590_A wire1285/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1117_A wire1118/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_194 _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output688_A _055_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_429_ _557_/A _429_/B _429_/C vssd vssd vccd vccd _429_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output855_A wire1406/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1653_A wire1654/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__302__B _302_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[0\]_A mprj_dat_i_user[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1820_A wire1821/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1918_A wire1918/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput1 caravel_clk vssd vssd vccd vccd _296_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] _272_/X vssd vssd vccd vccd _092_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_20_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__212__B _212_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3178 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1102 wire1103/X vssd vssd vccd vccd wire1102/X sky130_fd_sc_hd__buf_6
XFILLER_44_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1113 wire1114/X vssd vssd vccd vccd wire1113/X sky130_fd_sc_hd__buf_6
XFILLER_25_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1124 wire1124/A vssd vssd vccd vccd _078_/A sky130_fd_sc_hd__buf_6
XFILLER_19_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1135 wire1135/A vssd vssd vccd vccd _063_/A sky130_fd_sc_hd__buf_6
Xwire1146 _587_/X vssd vssd vccd vccd wire1146/X sky130_fd_sc_hd__buf_6
XFILLER_22_3994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1157 _550_/X vssd vssd vccd vccd wire1157/X sky130_fd_sc_hd__buf_6
XFILLER_47_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1168 _538_/X vssd vssd vccd vccd wire1168/X sky130_fd_sc_hd__buf_6
Xwire1179 _518_/X vssd vssd vccd vccd wire1179/X sky130_fd_sc_hd__buf_6
XFILLER_19_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input217_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__375__A_N _503_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2301_A wire2301/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_214_ _214_/A _214_/B vssd vssd vccd vccd _214_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_4076 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_145_ _145_/A vssd vssd vccd vccd _145_/Y sky130_fd_sc_hd__inv_12
XFILLER_32_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] max_cap1456/X vssd vssd vccd vccd _114_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_49_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_076_ _076_/A vssd vssd vccd vccd _076_/Y sky130_fd_sc_hd__inv_4
XFILLER_23_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1067_A wire1068/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1680 wire1680/A vssd vssd vccd vccd _596_/A sky130_fd_sc_hd__buf_6
XFILLER_39_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1234_A wire1235/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1691 wire1691/A vssd vssd vccd vccd _578_/A sky130_fd_sc_hd__buf_8
XFILLER_19_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1818 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] split5/X vssd vssd vccd vccd _144_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_33_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1770_A wire1771/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1868_A wire1869/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__313__A _313_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__398__A_N _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__207__B _207_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_50 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_61 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_72 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_83 _264_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_94 _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2084_A wire2085/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input167_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2251_A wire2251/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input334_A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input28_A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_128_ _128_/A vssd vssd vccd vccd _128_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_29_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output553_A _435_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__133__A _133_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_059_ _059_/A vssd vssd vccd vccd _059_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wire1184_A _513_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output720_A _597_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output818_A _571_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3566 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2990 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1351_A _353_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1449_A wire1450/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] _228_/X vssd vssd vccd vccd _048_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_40_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1616_A wire1616/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__308__A _308_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1985_A wire1985/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire971_A wire972/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput70 la_data_out_mprj[44] vssd vssd vccd vccd _413_/C sky130_fd_sc_hd__clkbuf_4
Xinput81 la_data_out_mprj[54] vssd vssd vccd vccd _423_/C sky130_fd_sc_hd__buf_4
Xinput92 la_data_out_mprj[64] vssd vssd vccd vccd input92/X sky130_fd_sc_hd__buf_6
XFILLER_45_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__218__A _218_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1314 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__413__A_N _541_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input284_A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2299_A wire2299/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input451_A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput430 mprj_dat_o_core[18] vssd vssd vccd vccd wire1529/A sky130_fd_sc_hd__buf_6
XFILLER_23_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput441 mprj_dat_o_core[28] vssd vssd vccd vccd wire1516/A sky130_fd_sc_hd__buf_6
XANTENNA__400__B _400_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput452 mprj_dat_o_core[9] vssd vssd vccd vccd wire1498/A sky130_fd_sc_hd__buf_6
XFILLER_2_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output768_A _526_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1399_A _327_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output935_A wire1391/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput904 wire970/X vssd vssd vccd vccd mprj_dat_i_core[30] sky130_fd_sc_hd__buf_8
Xoutput915 wire1364/X vssd vssd vccd vccd mprj_dat_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_28_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput926 wire1334/X vssd vssd vccd vccd mprj_dat_o_user[21] sky130_fd_sc_hd__buf_8
Xoutput937 wire1295/X vssd vssd vccd vccd mprj_dat_o_user[31] sky130_fd_sc_hd__buf_8
XFILLER_47_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput948 wire1426/X vssd vssd vccd vccd mprj_sel_o_user[3] sky130_fd_sc_hd__buf_8
XFILLER_25_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput959 _113_/Y vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__buf_8
XFILLER_25_2905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__310__B _310_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2302 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__A_N _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__038__A _038_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_600_ _600_/A _600_/B vssd vssd vccd vccd _600_/X sky130_fd_sc_hd__and2_4
XTAP_4258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2047_A wire2048/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_531_ _531_/A _531_/B vssd vssd vccd vccd _531_/X sky130_fd_sc_hd__and2_4
XTAP_2812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_462_ _590_/A _462_/B _462_/C vssd vssd vccd vccd _462_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2214_A wire2214/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_393_ _521_/A _393_/B _393_/C vssd vssd vccd vccd _393_/X sky130_fd_sc_hd__and3b_4
XFILLER_25_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input95_A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output516_A wire1261/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput260 la_oenb_mprj[0] vssd vssd vccd vccd _497_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput271 la_oenb_mprj[10] vssd vssd vccd vccd _507_/A sky130_fd_sc_hd__buf_4
XFILLER_49_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput282 la_oenb_mprj[11] vssd vssd vccd vccd _508_/A sky130_fd_sc_hd__buf_4
XFILLER_53_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput293 la_oenb_mprj[14] vssd vssd vccd vccd _511_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__459__A_N _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1147_A _586_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output885_A wire1051/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] _191_/X vssd vssd vccd vccd _011_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_982 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__305__B _305_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput701 _067_/Y vssd vssd vccd vccd la_data_in_mprj[84] sky130_fd_sc_hd__buf_8
Xoutput712 _077_/Y vssd vssd vccd vccd la_data_in_mprj[94] sky130_fd_sc_hd__buf_8
XANTENNA_wire1850_A wire1851/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput723 _600_/X vssd vssd vccd vccd la_oenb_core[103] sky130_fd_sc_hd__buf_8
XANTENNA_wire1948_A wire1948/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput734 _610_/X vssd vssd vccd vccd la_oenb_core[113] sky130_fd_sc_hd__buf_8
XFILLER_29_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput745 _620_/X vssd vssd vccd vccd la_oenb_core[123] sky130_fd_sc_hd__buf_8
Xoutput756 wire1182/X vssd vssd vccd vccd la_oenb_core[18] sky130_fd_sc_hd__buf_8
XFILLER_42_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput767 wire1173/X vssd vssd vccd vccd la_oenb_core[28] sky130_fd_sc_hd__buf_8
Xoutput778 wire1170/X vssd vssd vccd vccd la_oenb_core[38] sky130_fd_sc_hd__buf_8
XFILLER_29_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput789 _545_/X vssd vssd vccd vccd la_oenb_core[48] sky130_fd_sc_hd__buf_8
XANTENNA_powergood_check_mprj2_vdd_logic1 output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__321__A _321_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2818 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1509 wire1510/X vssd vssd vccd vccd _340_/B sky130_fd_sc_hd__buf_6
XTAP_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__215__B _215_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__231__A _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input247_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2164_A wire2164/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_split5_A split5/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input414_A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_514_ _514_/A _514_/B vssd vssd vccd vccd _514_/X sky130_fd_sc_hd__and2_2
XTAP_2653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_445_ _573_/A _445_/B _445_/C vssd vssd vccd vccd _445_/X sky130_fd_sc_hd__and3b_4
XTAP_1963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ _504_/A _376_/B _376_/C vssd vssd vccd vccd _376_/X sky130_fd_sc_hd__and3b_4
XFILLER_9_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_952 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output466_A wire1213/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_996 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1097_A wire1098/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output633_A _005_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3767 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__141__A _141_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output800_A wire1150/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1431_A wire1432/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1529_A wire1529/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__316__A _316_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput520 wire1257/X vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__buf_8
Xoutput531 wire1247/X vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__buf_8
XFILLER_44_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput542 wire1232/X vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__buf_8
Xoutput553 _435_/X vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__buf_8
XFILLER_43_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput564 _445_/X vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__buf_8
XFILLER_25_3244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput575 _455_/X vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__buf_8
XFILLER_47_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__051__A _051_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput586 wire1217/X vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__buf_8
Xwire2007 wire2008/X vssd vssd vccd vccd _619_/B sky130_fd_sc_hd__buf_6
Xoutput597 _088_/Y vssd vssd vccd vccd la_data_in_mprj[105] sky130_fd_sc_hd__buf_8
Xwire2018 wire2019/X vssd vssd vccd vccd wire2018/X sky130_fd_sc_hd__buf_6
Xwire2029 wire2030/X vssd vssd vccd vccd _612_/B sky130_fd_sc_hd__buf_6
Xwire1306 _366_/X vssd vssd vccd vccd wire1306/X sky130_fd_sc_hd__buf_6
XFILLER_5_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input2_A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1317 wire1318/X vssd vssd vccd vccd wire1317/X sky130_fd_sc_hd__buf_6
XFILLER_47_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1328 wire1329/X vssd vssd vccd vccd wire1328/X sky130_fd_sc_hd__buf_6
XFILLER_41_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1339 _357_/X vssd vssd vccd vccd wire1339/X sky130_fd_sc_hd__buf_6
XFILLER_38_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2372 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_230_ _230_/A _230_/B vssd vssd vccd vccd _230_/X sky130_fd_sc_hd__and2_2
XFILLER_14_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__226__A _226_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_161_ _161_/A vssd vssd vccd vccd _161_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_52_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input197_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_092_ _092_/A vssd vssd vccd vccd _092_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2281_A wire2281/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input364_A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input58_A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_966 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_454 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1840 wire1840/A vssd vssd vccd vccd wire1840/X sky130_fd_sc_hd__buf_6
Xwire1851 wire1852/X vssd vssd vccd vccd wire1851/X sky130_fd_sc_hd__buf_6
XFILLER_20_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1862 wire1863/X vssd vssd vccd vccd wire1862/X sky130_fd_sc_hd__buf_6
XFILLER_1_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1873 wire1874/X vssd vssd vccd vccd _282_/A sky130_fd_sc_hd__buf_6
XFILLER_18_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1884 wire1884/A vssd vssd vccd vccd _276_/A sky130_fd_sc_hd__buf_6
XTAP_3140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1895 wire1896/X vssd vssd vccd vccd _267_/A sky130_fd_sc_hd__buf_6
XTAP_3151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_151 _494_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _474_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 wire1760/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_184 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_428_ _556_/A _428_/B _428_/C vssd vssd vccd vccd _428_/X sky130_fd_sc_hd__and3b_4
XANTENNA_wire1012_A wire1013/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output583_A wire1220/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_359_ _359_/A _359_/B vssd vssd vccd vccd _359_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output750_A wire1188/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output848_A _305_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1479_A _243_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] wire1465/X vssd vssd vccd vccd wire1124/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_44_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1646_A wire1647/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[0\]_B max_cap1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1813_A wire1813/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput2 caravel_clk2 vssd vssd vccd vccd _297_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__046__A _046_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3282 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1103 wire1104/X vssd vssd vccd vccd wire1103/X sky130_fd_sc_hd__buf_6
XFILLER_48_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1114 wire1115/X vssd vssd vccd vccd wire1114/X sky130_fd_sc_hd__buf_6
XFILLER_48_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1125 wire1125/A vssd vssd vccd vccd _075_/A sky130_fd_sc_hd__buf_6
XFILLER_47_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1136 wire1136/A vssd vssd vccd vccd _062_/A sky130_fd_sc_hd__buf_6
Xwire1147 _586_/X vssd vssd vccd vccd wire1147/X sky130_fd_sc_hd__buf_6
Xwire1158 wire1159/X vssd vssd vccd vccd wire1158/X sky130_fd_sc_hd__buf_6
XFILLER_0_4470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1169 _536_/X vssd vssd vccd vccd wire1169/X sky130_fd_sc_hd__buf_6
XFILLER_38_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input112_A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2127_A wire2127/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_358 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_213_ _213_/A _213_/B vssd vssd vccd vccd _213_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_144_ _144_/A vssd vssd vccd vccd _144_/Y sky130_fd_sc_hd__inv_12
XFILLER_13_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_075_ _075_/A vssd vssd vccd vccd _075_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_13_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__403__B _403_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3895 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1670 wire1670/A vssd vssd vccd vccd wire1670/X sky130_fd_sc_hd__buf_6
Xwire1681 wire1681/A vssd vssd vccd vccd _595_/A sky130_fd_sc_hd__buf_6
Xwire1692 wire1692/A vssd vssd vccd vccd _577_/A sky130_fd_sc_hd__buf_8
XFILLER_18_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1227_A _429_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output798_A wire1153/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] rebuffer3/X vssd vssd vccd vccd _137_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_15_2553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] _173_/X vssd vssd vccd vccd _157_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_50_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1596_A wire1596/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1763_A wire1763/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__313__B _313_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1930_A wire1930/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] _284_/X vssd vssd vccd vccd wire1141/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_39_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_40 _321_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_51 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_62 _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_73 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_84 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_95 _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__504__A _504_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2077_A wire2077/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input327_A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2244_A wire2244/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3719 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_954 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__492__A_N _620_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_49_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_127_ _127_/A vssd vssd vccd vccd _127_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_29_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_058_ _058_/A vssd vssd vccd vccd _058_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output546_A wire1289/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1177_A _520_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output713_A _078_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1344_A wire1345/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2190 wire2190/A vssd vssd vccd vccd wire2190/X sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] _221_/X vssd vssd vccd vccd _041_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1511_A wire1511/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3316 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1609_A wire1610/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__308__B _308_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1978_A wire1978/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire964_A wire965/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_11_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput60 la_data_out_mprj[35] vssd vssd vccd vccd _404_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput71 la_data_out_mprj[45] vssd vssd vccd vccd _414_/C sky130_fd_sc_hd__clkbuf_4
Xinput82 la_data_out_mprj[55] vssd vssd vccd vccd _424_/C sky130_fd_sc_hd__buf_4
XFILLER_28_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput93 la_data_out_mprj[65] vssd vssd vccd vccd input93/X sky130_fd_sc_hd__buf_6
XFILLER_8_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1758 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__234__A _234_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2194_A wire2195/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input277_A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input444_A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input40_A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput420 mprj_cyc_o_core vssd vssd vccd vccd wire1552/A sky130_fd_sc_hd__buf_6
Xinput431 mprj_dat_o_core[19] vssd vssd vccd vccd wire1528/A sky130_fd_sc_hd__buf_6
XFILLER_40_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput442 mprj_dat_o_core[29] vssd vssd vccd vccd wire1515/A sky130_fd_sc_hd__buf_6
XANTENNA__400__C _400_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput453 mprj_iena_wb vssd vssd vccd vccd wire1496/A sky130_fd_sc_hd__buf_6
XFILLER_48_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output496_A wire1280/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__144__A _144_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__388__A_N _516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1294_A _369_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput905 wire966/X vssd vssd vccd vccd mprj_dat_i_core[31] sky130_fd_sc_hd__buf_8
XFILLER_49_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput916 wire1361/X vssd vssd vccd vccd mprj_dat_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_7_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output830_A _582_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput927 wire1331/X vssd vssd vccd vccd mprj_dat_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_28_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput938 wire1388/X vssd vssd vccd vccd mprj_dat_o_user[3] sky130_fd_sc_hd__buf_8
XANTENNA_output928_A wire1327/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput949 wire1449/X vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__buf_8
XFILLER_45_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1559_A wire1559/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3160 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__054__A _054_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__501__B _501_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_530_ _530_/A _530_/B vssd vssd vccd vccd _530_/X sky130_fd_sc_hd__and2_4
XTAP_3558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__229__A _229_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_461_ _589_/A _461_/B _461_/C vssd vssd vccd vccd _461_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_392_ _520_/A _392_/B _392_/C vssd vssd vccd vccd _392_/X sky130_fd_sc_hd__and3b_4
XFILLER_52_3571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2207_A wire2208/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input394_A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input88_A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__411__B _411_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput250 la_iena_mprj[91] vssd vssd vccd vccd _254_/B sky130_fd_sc_hd__clkbuf_4
Xinput261 la_oenb_mprj[100] vssd vssd vccd vccd wire1736/A sky130_fd_sc_hd__buf_6
Xinput272 la_oenb_mprj[110] vssd vssd vccd vccd _607_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_23_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput283 la_oenb_mprj[120] vssd vssd vccd vccd wire1727/A sky130_fd_sc_hd__buf_6
XFILLER_18_4101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output509_A wire1267/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput294 la_oenb_mprj[15] vssd vssd vccd vccd _512_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_18_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1042_A wire1043/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3466 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output780_A wire1197/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1307_A wire1308/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output878_A wire1422/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1676_A wire1677/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput702 _068_/Y vssd vssd vccd vccd la_data_in_mprj[85] sky130_fd_sc_hd__buf_8
XFILLER_9_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput713 _078_/Y vssd vssd vccd vccd la_data_in_mprj[95] sky130_fd_sc_hd__buf_8
Xoutput724 _601_/X vssd vssd vccd vccd la_oenb_core[104] sky130_fd_sc_hd__buf_8
XFILLER_25_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput735 _611_/X vssd vssd vccd vccd la_oenb_core[114] sky130_fd_sc_hd__buf_8
XANTENNA__602__A _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput746 _621_/X vssd vssd vccd vccd la_oenb_core[124] sky130_fd_sc_hd__buf_8
Xoutput757 wire1181/X vssd vssd vccd vccd la_oenb_core[19] sky130_fd_sc_hd__buf_8
XFILLER_47_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1843_A wire1843/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput768 _526_/X vssd vssd vccd vccd la_oenb_core[29] sky130_fd_sc_hd__buf_8
Xoutput779 wire1169/X vssd vssd vccd vccd la_oenb_core[39] sky130_fd_sc_hd__buf_8
XANTENNA__321__B _321_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__403__A_N _531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__049__A _049_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__512__A _512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__231__B _231_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input142_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2157_A wire2157/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input407_A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_513_ _513_/A _513_/B vssd vssd vccd vccd _513_/X sky130_fd_sc_hd__and2_2
XFILLER_22_1291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_444_ _572_/A _444_/B _444_/C vssd vssd vccd vccd _444_/X sky130_fd_sc_hd__and3b_4
XTAP_2687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_375_ _503_/A _375_/B _375_/C vssd vssd vccd vccd _375_/X sky130_fd_sc_hd__and3b_4
XTAP_1997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_964 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__426__A_N _554_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1257_A _405_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1424_A wire1425/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] _203_/X vssd vssd vccd vccd _023_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_20_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1793_A wire1794/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__316__B _316_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[90\]_B wire1469/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput510 wire1266/X vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__buf_8
XANTENNA__332__A _332_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput521 wire1256/X vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__buf_8
Xoutput532 wire1246/X vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__buf_8
XFILLER_44_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput543 wire1231/X vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__buf_8
XFILLER_9_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput554 _436_/X vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] _165_/X vssd vssd vccd vccd _149_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput565 _446_/X vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__buf_8
XFILLER_5_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput576 _456_/X vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__buf_8
Xoutput587 _466_/X vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__buf_8
Xwire2008 wire2009/X vssd vssd vccd vccd wire2008/X sky130_fd_sc_hd__buf_6
XFILLER_25_3267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput598 _089_/Y vssd vssd vccd vccd la_data_in_mprj[106] sky130_fd_sc_hd__buf_8
Xwire2019 wire2019/A vssd vssd vccd vccd wire2019/X sky130_fd_sc_hd__buf_6
XFILLER_5_2616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1307 wire1308/X vssd vssd vccd vccd wire1307/X sky130_fd_sc_hd__buf_8
XFILLER_21_2419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1318 _363_/X vssd vssd vccd vccd wire1318/X sky130_fd_sc_hd__buf_6
XFILLER_3_3052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1329 wire1330/X vssd vssd vccd vccd wire1329/X sky130_fd_sc_hd__buf_6
XFILLER_20_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__507__A _507_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_160_ _160_/A vssd vssd vccd vccd _160_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__226__B _226_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_091_ _091_/A vssd vssd vccd vccd _091_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[81\]_B wire1478/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__449__A_N _577_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__242__A _242_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2274_A wire2274/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input357_A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1830 wire1830/A vssd vssd vccd vccd _356_/A sky130_fd_sc_hd__buf_6
XFILLER_19_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1841 wire1842/X vssd vssd vccd vccd _293_/A sky130_fd_sc_hd__buf_6
XFILLER_18_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1852 wire1852/A vssd vssd vccd vccd wire1852/X sky130_fd_sc_hd__buf_6
XFILLER_19_835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1863 wire1863/A vssd vssd vccd vccd wire1863/X sky130_fd_sc_hd__buf_6
Xwire1874 wire1874/A vssd vssd vccd vccd wire1874/X sky130_fd_sc_hd__buf_6
XFILLER_37_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1885 wire1885/A vssd vssd vccd vccd _275_/A sky130_fd_sc_hd__buf_6
XTAP_3141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1896 wire1896/A vssd vssd vccd vccd wire1896/X sky130_fd_sc_hd__buf_6
XTAP_3152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 _494_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_163 _474_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 wire1758/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_196 _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_427_ _555_/A _427_/B _427_/C vssd vssd vccd vccd _427_/X sky130_fd_sc_hd__and3b_4
XTAP_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_358_ _358_/A _358_/B vssd vssd vccd vccd _358_/X sky130_fd_sc_hd__and2_4
XFILLER_31_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1005_A _137_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output576_A _456_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_289_ _289_/A _289_/B vssd vssd vccd vccd _289_/X sky130_fd_sc_hd__and2_1
XFILLER_31_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[72\]_B _235_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output743_A _618_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1374_A wire1375/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output910_A wire1081/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] wire1471/X vssd vssd vccd vccd wire1127/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_26_3587 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1639_A wire1639/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput3 caravel_rstn vssd vssd vccd vccd input3/X sky130_fd_sc_hd__buf_6
XFILLER_37_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1806_A wire1807/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire994_A wire995/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__327__A _327_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4019 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__062__A _062_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2639 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1104 wire1105/X vssd vssd vccd vccd wire1104/X sky130_fd_sc_hd__buf_6
XFILLER_44_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1115 _115_/Y vssd vssd vccd vccd wire1115/X sky130_fd_sc_hd__buf_6
XFILLER_22_3974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1126 wire1126/A vssd vssd vccd vccd _074_/A sky130_fd_sc_hd__buf_6
XFILLER_38_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1137 wire1137/A vssd vssd vccd vccd _061_/A sky130_fd_sc_hd__buf_6
XFILLER_47_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1148 _558_/X vssd vssd vccd vccd wire1148/X sky130_fd_sc_hd__buf_6
XFILLER_21_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1159 _549_/X vssd vssd vccd vccd wire1159/X sky130_fd_sc_hd__buf_6
XFILLER_0_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2022_A wire2022/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__237__A _237_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_370 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_690 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_212_ _212_/A _212_/B vssd vssd vccd vccd _212_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_143_ _143_/A vssd vssd vccd vccd _143_/Y sky130_fd_sc_hd__inv_12
XFILLER_11_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[54\]_B _217_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input70_A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_074_ _074_/A vssd vssd vccd vccd _074_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__403__C _403_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_230 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_4257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1660 wire1661/X vssd vssd vccd vccd wire1660/X sky130_fd_sc_hd__buf_6
Xwire1671 wire1672/X vssd vssd vccd vccd _316_/B sky130_fd_sc_hd__buf_6
XFILLER_19_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1682 wire1682/A vssd vssd vccd vccd _594_/A sky130_fd_sc_hd__buf_6
Xwire1693 wire1693/A vssd vssd vccd vccd _576_/A sky130_fd_sc_hd__buf_8
XFILLER_18_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1122_A wire1122/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output693_A _060_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output860_A wire1400/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] load_slew1458/X vssd vssd vccd vccd _130_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1491_A wire1491/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1589_A wire1590/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1728 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire990 wire991/X vssd vssd vccd vccd wire990/X sky130_fd_sc_hd__buf_6
XFILLER_41_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1756_A wire1757/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__610__A _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] _277_/X vssd vssd vccd vccd _097_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__057__A _057_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_30 _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_41 _321_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_52 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_63 _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_74 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_85 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_96 _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__504__B _504_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_B _283_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__520__A _520_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1902 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input222_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2237_A wire2238/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_4189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_126_ _126_/A vssd vssd vccd vccd _126_/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__414__B _414_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B _274_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_057_ _057_/A vssd vssd vccd vccd _057_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3671 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output539_A wire1238/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1072_A wire1073/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output706_A _072_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2180 wire2181/X vssd vssd vccd vccd wire2180/X sky130_fd_sc_hd__buf_6
XFILLER_43_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2191 wire2192/X vssd vssd vccd vccd _488_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire1337_A wire1338/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1490 input91/X vssd vssd vccd vccd _432_/C sky130_fd_sc_hd__buf_6
XFILLER_17_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1504_A wire1504/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[20\]_A mprj_dat_i_user[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__605__A _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1873_A wire1874/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__324__B _324_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_B _265_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput50 la_data_out_mprj[26] vssd vssd vccd vccd _395_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput61 la_data_out_mprj[36] vssd vssd vccd vccd _405_/C sky130_fd_sc_hd__clkbuf_4
Xinput72 la_data_out_mprj[46] vssd vssd vccd vccd _415_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput83 la_data_out_mprj[56] vssd vssd vccd vccd _425_/C sky130_fd_sc_hd__buf_4
XFILLER_28_2701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput94 la_data_out_mprj[66] vssd vssd vccd vccd input94/X sky130_fd_sc_hd__buf_6
XFILLER_28_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__340__A _340_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_900 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[11\]_A mprj_dat_i_user[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__515__A _515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__234__B _234_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input172_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2187_A wire2187/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__250__A _250_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_4341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input437_A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput410 mprj_adr_o_core[2] vssd vssd vccd vccd wire1596/A sky130_fd_sc_hd__buf_6
XFILLER_7_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput421 mprj_dat_o_core[0] vssd vssd vccd vccd wire1548/A sky130_fd_sc_hd__buf_6
XFILLER_24_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input33_A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput432 mprj_dat_o_core[1] vssd vssd vccd vccd wire1527/A sky130_fd_sc_hd__buf_6
XFILLER_0_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput443 mprj_dat_o_core[2] vssd vssd vccd vccd wire1514/A sky130_fd_sc_hd__buf_6
XFILLER_40_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput454 mprj_sel_o_core[0] vssd vssd vccd vccd _301_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3590 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__409__B _409_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output489_A wire1205/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output656_A _026_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_109_ _109_/A vssd vssd vccd vccd _109_/Y sky130_fd_sc_hd__inv_2
Xoutput906 wire1101/X vssd vssd vccd vccd mprj_dat_i_core[3] sky130_fd_sc_hd__buf_8
Xoutput917 wire1358/X vssd vssd vccd vccd mprj_dat_o_user[13] sky130_fd_sc_hd__buf_8
XFILLER_45_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput928 wire1327/X vssd vssd vccd vccd mprj_dat_o_user[23] sky130_fd_sc_hd__buf_8
XFILLER_7_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1287_A _376_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput939 wire1385/X vssd vssd vccd vccd mprj_dat_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_45_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output823_A _576_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__160__A _160_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1454_A wire1455/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] _233_/X vssd vssd vccd vccd _053_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1621_A wire1621/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__319__B _319_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1990_A wire1991/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__335__A _335_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__482__A_N _610_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__070__A _070_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_460_ _588_/A _460_/B _460_/C vssd vssd vccd vccd _460_/X sky130_fd_sc_hd__and3b_4
XANTENNA__229__B _229_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_391_ _519_/A _391_/B _391_/C vssd vssd vccd vccd _391_/X sky130_fd_sc_hd__and3b_4
XFILLER_53_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2102_A wire2102/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__245__A _245_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input387_A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput240 la_iena_mprj[82] vssd vssd vccd vccd _245_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput251 la_iena_mprj[92] vssd vssd vccd vccd _255_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput262 la_oenb_mprj[101] vssd vssd vccd vccd _598_/A sky130_fd_sc_hd__buf_4
Xinput273 la_oenb_mprj[111] vssd vssd vccd vccd _608_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_23_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput284 la_oenb_mprj[121] vssd vssd vccd vccd wire1726/A sky130_fd_sc_hd__buf_6
XFILLER_18_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput295 la_oenb_mprj[16] vssd vssd vccd vccd _513_/A sky130_fd_sc_hd__buf_4
XFILLER_18_3401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1035_A _131_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_3347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_589_ _589_/A _589_/B vssd vssd vccd vccd _589_/X sky130_fd_sc_hd__and2_4
XFILLER_32_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1202_A _495_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output773_A wire1172/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__155__A _155_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output940_A wire1382/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput703 _069_/Y vssd vssd vccd vccd la_data_in_mprj[86] sky130_fd_sc_hd__buf_8
XANTENNA_wire1571_A wire1571/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1669_A wire1670/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput714 _079_/Y vssd vssd vccd vccd la_data_in_mprj[96] sky130_fd_sc_hd__buf_8
Xoutput725 _602_/X vssd vssd vccd vccd la_oenb_core[105] sky130_fd_sc_hd__buf_8
XFILLER_47_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput736 _612_/X vssd vssd vccd vccd la_oenb_core[115] sky130_fd_sc_hd__buf_8
XANTENNA__602__B _602_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput747 _622_/X vssd vssd vccd vccd la_oenb_core[125] sky130_fd_sc_hd__buf_8
Xoutput758 wire1199/X vssd vssd vccd vccd la_oenb_core[1] sky130_fd_sc_hd__buf_8
XFILLER_42_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput769 wire1198/X vssd vssd vccd vccd la_oenb_core[2] sky130_fd_sc_hd__buf_8
XFILLER_47_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__065__A _065_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__512__B _512_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3983 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3994 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2052_A wire2053/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__378__A_N _506_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_512_ _512_/A _512_/B vssd vssd vccd vccd _512_/X sky130_fd_sc_hd__and2_2
XTAP_2622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input302_A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ _571_/A _443_/B _443_/C vssd vssd vccd vccd _443_/X sky130_fd_sc_hd__and3b_4
XTAP_2677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ _502_/A _374_/B _374_/C vssd vssd vccd vccd _374_/X sky130_fd_sc_hd__and3b_4
XTAP_1987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__406__C _406_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__422__B _422_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output521_A wire1256/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output619_A _108_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1417_A wire1418/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output890_A wire1026/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] _196_/X vssd vssd vccd vccd _016_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_14_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2730 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1786_A wire1787/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__613__A _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1953_A wire1953/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput500 wire1276/X vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__buf_8
Xoutput511 wire1265/X vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__buf_8
XFILLER_9_3432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput522 wire1255/X vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__buf_8
XANTENNA__332__B _332_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput533 wire1245/X vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__buf_8
XFILLER_47_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput544 wire1229/X vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__buf_8
Xoutput555 _437_/X vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__buf_8
Xoutput566 _447_/X vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_A mprj_dat_i_user[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput577 _457_/X vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__buf_8
XFILLER_5_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput588 _467_/X vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__buf_8
Xwire2009 wire2009/A vssd vssd vccd vccd wire2009/X sky130_fd_sc_hd__buf_6
XFILLER_25_2534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput599 _090_/Y vssd vssd vccd vccd la_data_in_mprj[107] sky130_fd_sc_hd__buf_8
XFILLER_29_1991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1308 wire1309/X vssd vssd vccd vccd wire1308/X sky130_fd_sc_hd__buf_6
XFILLER_5_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1319 wire1320/X vssd vssd vccd vccd wire1319/X sky130_fd_sc_hd__buf_8
XFILLER_41_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__507__B _507_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_090_ _090_/A vssd vssd vccd vccd _090_/Y sky130_fd_sc_hd__inv_2
XANTENNA__523__A _523_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__242__B _242_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input252_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1820 wire1821/X vssd vssd vccd vccd _364_/A sky130_fd_sc_hd__buf_6
XFILLER_8_1573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1831 wire1831/A vssd vssd vccd vccd _355_/A sky130_fd_sc_hd__buf_6
XFILLER_1_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1842 wire1843/X vssd vssd vccd vccd wire1842/X sky130_fd_sc_hd__buf_6
Xwire1853 wire1854/X vssd vssd vccd vccd _289_/A sky130_fd_sc_hd__buf_6
Xwire1864 wire1865/X vssd vssd vccd vccd _285_/A sky130_fd_sc_hd__buf_6
XTAP_3120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1875 wire1876/X vssd vssd vccd vccd _281_/A sky130_fd_sc_hd__buf_6
XTAP_3131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1886 wire1886/A vssd vssd vccd vccd _274_/A sky130_fd_sc_hd__buf_6
XFILLER_19_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1897 wire1898/X vssd vssd vccd vccd _266_/A sky130_fd_sc_hd__buf_6
XTAP_3153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_142 _512_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _494_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_164 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_175 _489_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_426_ _554_/A _426_/B _426_/C vssd vssd vccd vccd _426_/X sky130_fd_sc_hd__and3b_4
XTAP_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _342_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__417__B _417_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _357_/A _357_/B vssd vssd vccd vccd _357_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_288_ _288_/A _288_/B vssd vssd vccd vccd _288_/X sky130_fd_sc_hd__and2_2
XANTENNA_output471_A wire1208/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output569_A _449_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output736_A _612_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1367_A wire1368/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output903_A wire1106/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1534_A wire1535/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput4 la_data_out_mprj[0] vssd vssd vccd vccd _369_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_20_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__608__A _608_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__327__B _327_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire987_A wire988/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3868 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__343__A _343_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2607 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1105 _117_/Y vssd vssd vccd vccd wire1105/X sky130_fd_sc_hd__buf_6
XFILLER_40_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1116 wire1117/X vssd vssd vccd vccd wire1116/X sky130_fd_sc_hd__buf_6
Xwire1127 wire1127/A vssd vssd vccd vccd _071_/A sky130_fd_sc_hd__buf_6
XFILLER_5_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1138 wire1138/A vssd vssd vccd vccd _060_/A sky130_fd_sc_hd__buf_6
Xwire1149 _557_/X vssd vssd vccd vccd wire1149/X sky130_fd_sc_hd__buf_6
XFILLER_38_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__A _518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__237__B _237_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__416__A_N _416_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2015_A wire2015/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_211_ _211_/A _211_/B vssd vssd vccd vccd _211_/X sky130_fd_sc_hd__and2_4
XFILLER_49_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_142_ _142_/A vssd vssd vccd vccd _142_/Y sky130_fd_sc_hd__inv_12
XFILLER_32_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2611 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_1191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__253__A _253_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_073_ _073_/A vssd vssd vccd vccd _073_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input63_A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_286 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_load_slew1457_A load_slew1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1650 wire1651/X vssd vssd vccd vccd wire1650/X sky130_fd_sc_hd__buf_6
XFILLER_1_2812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1661 wire1662/X vssd vssd vccd vccd wire1661/X sky130_fd_sc_hd__buf_6
XFILLER_21_3496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1672 wire1672/A vssd vssd vccd vccd wire1672/X sky130_fd_sc_hd__buf_6
XFILLER_18_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1683 wire1683/A vssd vssd vccd vccd _593_/A sky130_fd_sc_hd__buf_6
XFILLER_20_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1694 _447_/A_N vssd vssd vccd vccd _575_/A sky130_fd_sc_hd__buf_6
XFILLER_20_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1115_A _115_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output686_A _053_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_409_ _409_/A_N _409_/B _409_/C vssd vssd vccd vccd _409_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output853_A wire1408/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__163__A _163_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire980 wire981/X vssd vssd vccd vccd wire980/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1484_A input97/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire991 _140_/Y vssd vssd vccd vccd wire991/X sky130_fd_sc_hd__buf_6
XFILLER_6_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1651_A wire1651/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1749_A wire1749/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__610__B _610_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2322 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] _270_/X vssd vssd vccd vccd _090_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_53_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__439__A_N _567_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__338__A _338_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_20 _222_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_31 _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_42 _321_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_53 _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_64 _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_75 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__073__A _073_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_86 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_97 _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__520__B _520_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1914 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input215_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__248__A _248_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_125_ _125_/A vssd vssd vccd vccd _125_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__414__C _414_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_056_ _056_/A vssd vssd vccd vccd _056_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_27_4373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__430__B _430_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1065_A _125_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2170 wire2170/A vssd vssd vccd vccd wire2170/X sky130_fd_sc_hd__buf_6
XFILLER_21_3271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2181 wire2181/A vssd vssd vccd vccd wire2181/X sky130_fd_sc_hd__buf_6
Xwire2192 wire2193/X vssd vssd vccd vccd wire2192/X sky130_fd_sc_hd__buf_6
XFILLER_43_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1480 _242_/X vssd vssd vccd vccd wire1480/X sky130_fd_sc_hd__buf_6
XFILLER_1_3398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1491 wire1491/A vssd vssd vccd vccd _300_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire1232_A wire1233/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__158__A _158_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_B load_slew1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__605__B _605_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1504 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput40 la_data_out_mprj[17] vssd vssd vccd vccd _386_/C sky130_fd_sc_hd__clkbuf_4
Xinput51 la_data_out_mprj[27] vssd vssd vccd vccd _396_/C sky130_fd_sc_hd__clkbuf_4
Xinput62 la_data_out_mprj[37] vssd vssd vccd vccd _406_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput73 la_data_out_mprj[47] vssd vssd vccd vccd _416_/C sky130_fd_sc_hd__clkbuf_4
Xinput84 la_data_out_mprj[57] vssd vssd vccd vccd _426_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_7_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput95 la_data_out_mprj[67] vssd vssd vccd vccd input95/X sky130_fd_sc_hd__buf_6
XFILLER_45_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__621__A _621_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__340__B _340_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_912 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__068__A _068_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__515__B _515_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__531__A _531_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input165_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2082_A wire2082/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput400 mprj_adr_o_core[20] vssd vssd vccd vccd wire1639/A sky130_fd_sc_hd__buf_6
Xinput411 mprj_adr_o_core[30] vssd vssd vccd vccd wire1591/A sky130_fd_sc_hd__buf_6
XFILLER_2_4353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput422 mprj_dat_o_core[10] vssd vssd vccd vccd wire1545/A sky130_fd_sc_hd__buf_6
XFILLER_7_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input332_A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput433 mprj_dat_o_core[20] vssd vssd vccd vccd wire1524/A sky130_fd_sc_hd__buf_6
XFILLER_48_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput444 mprj_dat_o_core[30] vssd vssd vccd vccd wire1512/A sky130_fd_sc_hd__buf_6
XFILLER_0_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput455 mprj_sel_o_core[1] vssd vssd vccd vccd _302_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input26_A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__409__C _409_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__425__B _425_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4446 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_108_ _108_/A vssd vssd vccd vccd _108_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput907 wire1096/X vssd vssd vccd vccd mprj_dat_i_core[4] sky130_fd_sc_hd__buf_8
XFILLER_49_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output551_A _433_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput918 wire1355/X vssd vssd vccd vccd mprj_dat_o_user[14] sky130_fd_sc_hd__buf_8
Xoutput929 wire1323/X vssd vssd vccd vccd mprj_dat_o_user[24] sky130_fd_sc_hd__buf_8
XFILLER_7_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_039_ _039_/A vssd vssd vccd vccd _039_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1182_A _515_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output816_A _569_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1447_A wire1448/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] _226_/X vssd vssd vccd vccd _046_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_27_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1614_A wire1615/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__616__A _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__335__B _335_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__351__A _351_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_390_ _518_/A _390_/B _390_/C vssd vssd vccd vccd _390_/X sky130_fd_sc_hd__and3b_4
XFILLER_52_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__526__A _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input282_A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2297_A wire2297/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__261__A _261_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput230 la_iena_mprj[73] vssd vssd vccd vccd _236_/B sky130_fd_sc_hd__clkbuf_4
Xinput241 la_iena_mprj[83] vssd vssd vccd vccd _246_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput252 la_iena_mprj[93] vssd vssd vccd vccd _256_/B sky130_fd_sc_hd__clkbuf_4
Xinput263 la_oenb_mprj[102] vssd vssd vccd vccd _599_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_40_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput274 la_oenb_mprj[112] vssd vssd vccd vccd wire1735/A sky130_fd_sc_hd__buf_6
XFILLER_2_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput285 la_oenb_mprj[122] vssd vssd vccd vccd _619_/A sky130_fd_sc_hd__buf_4
XFILLER_53_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput296 la_oenb_mprj[17] vssd vssd vccd vccd _514_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_4027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_588_ _588_/A _588_/B vssd vssd vccd vccd _588_/X sky130_fd_sc_hd__and2_1
XANTENNA_wire1028_A wire1029/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output599_A _090_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output766_A _524_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1397_A _328_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output933_A wire1307/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput704 _070_/Y vssd vssd vccd vccd la_data_in_mprj[87] sky130_fd_sc_hd__buf_8
XFILLER_29_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput715 _080_/Y vssd vssd vccd vccd la_data_in_mprj[97] sky130_fd_sc_hd__buf_8
XANTENNA__171__A _171_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput726 _603_/X vssd vssd vccd vccd la_oenb_core[106] sky130_fd_sc_hd__buf_8
XFILLER_42_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput737 _613_/X vssd vssd vccd vccd la_oenb_core[116] sky130_fd_sc_hd__buf_8
XFILLER_47_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1564_A wire1565/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput748 wire1144/X vssd vssd vccd vccd la_oenb_core[126] sky130_fd_sc_hd__buf_8
XFILLER_7_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput759 wire1180/X vssd vssd vccd vccd la_oenb_core[20] sky130_fd_sc_hd__buf_8
XFILLER_42_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1731_A wire1731/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1829_A wire1829/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2556 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__346__A _346_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__081__A _081_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input128_A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2045_A wire2046/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ _511_/A _511_/B vssd vssd vccd vccd _511_/X sky130_fd_sc_hd__and2_4
XTAP_3368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _570_/A _442_/B _442_/C vssd vssd vccd vccd _442_/X sky130_fd_sc_hd__and3b_4
XANTENNA_wire2212_A wire2213/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__256__A _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_373_ _501_/A _373_/B _373_/C vssd vssd vccd vccd _373_/X sky130_fd_sc_hd__and3b_4
XTAP_1988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input93_A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] max_cap1456/X vssd vssd vccd vccd _123_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_4427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__422__C _422_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output514_A wire1263/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1312_A wire1313/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output883_A wire1061/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__472__A_N _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_3118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__166__A _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] _189_/X vssd vssd vccd vccd _009_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1779_A wire1779/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__613__B _613_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput501 wire1275/X vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__buf_8
Xoutput512 wire1264/X vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__buf_8
XFILLER_29_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput523 wire1254/X vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__buf_8
XFILLER_9_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput534 wire1244/X vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__buf_8
XFILLER_44_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1946_A wire1947/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput545 wire1228/X vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__buf_8
XFILLER_47_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput556 _438_/X vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_B max_cap1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput567 _448_/X vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__buf_8
XFILLER_5_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput578 wire1224/X vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__buf_8
Xoutput589 wire1216/X vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__buf_8
XFILLER_47_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1309 wire1310/X vssd vssd vccd vccd wire1309/X sky130_fd_sc_hd__buf_6
XFILLER_25_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_4391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__076__A _076_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__523__B _523_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2162_A wire2162/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input245_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1810 wire1811/X vssd vssd vccd vccd _368_/A sky130_fd_sc_hd__buf_6
XFILLER_41_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1821 wire1821/A vssd vssd vccd vccd wire1821/X sky130_fd_sc_hd__buf_6
XFILLER_8_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1832 wire1832/A vssd vssd vccd vccd _300_/A sky130_fd_sc_hd__buf_6
XFILLER_46_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1843 wire1843/A vssd vssd vccd vccd wire1843/X sky130_fd_sc_hd__buf_6
XFILLER_1_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1854 wire1855/X vssd vssd vccd vccd wire1854/X sky130_fd_sc_hd__buf_6
XTAP_3110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1865 wire1866/X vssd vssd vccd vccd wire1865/X sky130_fd_sc_hd__buf_6
XTAP_3121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input412_A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1876 wire1876/A vssd vssd vccd vccd wire1876/X sky130_fd_sc_hd__buf_6
XFILLER_46_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__495__A_N _623_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1887 wire1887/A vssd vssd vccd vccd _273_/A sky130_fd_sc_hd__buf_6
XTAP_3143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1898 wire1898/A vssd vssd vccd vccd wire1898/X sky130_fd_sc_hd__buf_6
XFILLER_37_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_110 _192_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _512_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_154 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _558_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_425_ _553_/A _425_/B _425_/C vssd vssd vccd vccd _425_/X sky130_fd_sc_hd__and3b_2
XANTENNA_187 _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _340_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__417__C _417_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_356_ _356_/A _356_/B vssd vssd vccd vccd _356_/X sky130_fd_sc_hd__and2_4
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_287_ _287_/A _287_/B vssd vssd vccd vccd _287_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__433__B _433_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_741 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output464_A wire1215/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output631_A _003_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output729_A _606_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2888 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput5 la_data_out_mprj[100] vssd vssd vccd vccd _469_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1527_A wire1527/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3188 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__608__B _608_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3994 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__624__A _624_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__343__B _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1106 wire1107/X vssd vssd vccd vccd wire1106/X sky130_fd_sc_hd__buf_6
Xwire1117 wire1118/X vssd vssd vccd vccd wire1117/X sky130_fd_sc_hd__buf_6
Xwire1128 wire1128/A vssd vssd vccd vccd _070_/A sky130_fd_sc_hd__buf_6
XFILLER_38_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1139 wire1139/A vssd vssd vccd vccd _106_/A sky130_fd_sc_hd__buf_6
XFILLER_19_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3998 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__518__B _518_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_210_ _210_/A _210_/B vssd vssd vccd vccd _210_/X sky130_fd_sc_hd__and2_4
XFILLER_51_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2008_A wire2009/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__534__A _534_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
X_141_ _141_/A vssd vssd vccd vccd _141_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_32_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input195_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2623 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_072_ _072_/A vssd vssd vccd vccd _072_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1679 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input362_A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input56_A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1640 wire1641/X vssd vssd vccd vccd _306_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2824 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1651 wire1651/A vssd vssd vccd vccd wire1651/X sky130_fd_sc_hd__buf_6
Xwire1662 wire1662/A vssd vssd vccd vccd wire1662/X sky130_fd_sc_hd__buf_6
Xwire1673 wire1674/X vssd vssd vccd vccd _315_/B sky130_fd_sc_hd__buf_6
XFILLER_19_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1684 wire1684/A vssd vssd vccd vccd _585_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1695 wire1695/A vssd vssd vccd vccd _574_/A sky130_fd_sc_hd__buf_8
XFILLER_46_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__428__B _428_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_408_ _536_/A _408_/B _408_/C vssd vssd vccd vccd _408_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output581_A wire1222/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1108_A wire1109/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output679_A _047_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_339_ _339_/A _339_/B vssd vssd vccd vccd _339_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire970 wire971/X vssd vssd vccd vccd wire970/X sky130_fd_sc_hd__buf_6
XANTENNA_output846_A wire1191/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire981 _142_/Y vssd vssd vccd vccd wire981/X sky130_fd_sc_hd__buf_6
Xwire992 wire993/X vssd vssd vccd vccd wire992/X sky130_fd_sc_hd__buf_6
XFILLER_31_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1477_A _245_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] wire1466/X vssd vssd vccd vccd _076_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_41_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1644_A wire1644/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1168 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3182 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1811_A wire1811/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1909_A wire1910/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__619__A _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__338__B _338_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_10 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_21 _223_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_32 _588_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__354__A _354_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_43 _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_54 _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_65 _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3092 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_76 _290_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_87 _243_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_98 _231_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3784 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__529__A _529_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input110_A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input208_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1243 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__264__A _264_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_124_ _124_/A vssd vssd vccd vccd _124_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_49_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_055_ _055_/A vssd vssd vccd vccd _055_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_49_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__430__C _430_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2160 wire2160/A vssd vssd vccd vccd _501_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2171 wire2172/X vssd vssd vccd vccd _495_/B sky130_fd_sc_hd__buf_6
XFILLER_1_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2182 wire2183/X vssd vssd vccd vccd _491_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2193 wire2193/A vssd vssd vccd vccd wire2193/X sky130_fd_sc_hd__buf_6
XFILLER_21_3283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1058_A wire1059/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1470 _252_/X vssd vssd vccd vccd wire1470/X sky130_fd_sc_hd__buf_8
XFILLER_53_209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1481 _241_/X vssd vssd vccd vccd wire1481/X sky130_fd_sc_hd__buf_6
Xwire1492 wire1493/X vssd vssd vccd vccd _299_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output796_A _551_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__174__A _174_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] load_slew1458/X vssd vssd vccd vccd _135_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_15_2375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1594_A wire1595/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput30 la_data_out_mprj[123] vssd vssd vccd vccd _492_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput41 la_data_out_mprj[18] vssd vssd vccd vccd _387_/C sky130_fd_sc_hd__clkbuf_4
Xinput52 la_data_out_mprj[28] vssd vssd vccd vccd _397_/C sky130_fd_sc_hd__clkbuf_4
Xinput63 la_data_out_mprj[38] vssd vssd vccd vccd _407_/C sky130_fd_sc_hd__clkbuf_4
Xinput74 la_data_out_mprj[48] vssd vssd vccd vccd _417_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1761_A wire1761/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput85 la_data_out_mprj[58] vssd vssd vccd vccd _427_/C sky130_fd_sc_hd__buf_4
XFILLER_41_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput96 la_data_out_mprj[68] vssd vssd vccd vccd input96/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1859_A wire1860/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__621__B _621_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__406__A_N _406_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__349__A _349_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4401 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__084__A _084_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1004 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__531__B _531_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2075_A wire2075/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input158_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput401 mprj_adr_o_core[21] vssd vssd vccd vccd wire1636/A sky130_fd_sc_hd__buf_6
Xinput412 mprj_adr_o_core[31] vssd vssd vccd vccd wire1586/A sky130_fd_sc_hd__buf_6
XFILLER_22_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput423 mprj_dat_o_core[11] vssd vssd vccd vccd wire1543/A sky130_fd_sc_hd__buf_6
XFILLER_40_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput434 mprj_dat_o_core[21] vssd vssd vccd vccd wire1523/A sky130_fd_sc_hd__buf_6
XFILLER_40_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput445 mprj_dat_o_core[31] vssd vssd vccd vccd wire1511/A sky130_fd_sc_hd__buf_6
XFILLER_2_4387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput456 mprj_sel_o_core[2] vssd vssd vccd vccd _303_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire2242_A wire2243/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input325_A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__259__A _259_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input19_A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__425__C _425_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4458 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_107_ _107_/A vssd vssd vccd vccd _107_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput908 wire1091/X vssd vssd vccd vccd mprj_dat_i_core[5] sky130_fd_sc_hd__buf_8
Xoutput919 wire1352/X vssd vssd vccd vccd mprj_dat_o_user[15] sky130_fd_sc_hd__buf_8
XFILLER_45_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__429__A_N _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_038_ _038_/A vssd vssd vccd vccd _038_/Y sky130_fd_sc_hd__inv_2
XANTENNA__441__B _441_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output544_A wire1229/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1022 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output711_A _076_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1342_A _356_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__169__A _169_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] _219_/X vssd vssd vccd vccd _039_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_35_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1607_A wire1608/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__616__B _616_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3750 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1976_A wire1976/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire962_A wire963/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2036 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__351__B _351_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2616 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__079__A _079_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__526__B _526_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__542__A _542_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2192_A wire2193/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input275_A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__261__B _261_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input442_A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput220 la_iena_mprj[64] vssd vssd vccd vccd _227_/B sky130_fd_sc_hd__buf_4
XFILLER_1_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput231 la_iena_mprj[74] vssd vssd vccd vccd _237_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput242 la_iena_mprj[84] vssd vssd vccd vccd _247_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput253 la_iena_mprj[94] vssd vssd vccd vccd _257_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput264 la_oenb_mprj[103] vssd vssd vccd vccd _600_/A sky130_fd_sc_hd__clkbuf_8
Xinput275 la_oenb_mprj[113] vssd vssd vccd vccd wire1734/A sky130_fd_sc_hd__buf_6
XFILLER_2_3483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput286 la_oenb_mprj[123] vssd vssd vccd vccd _620_/A sky130_fd_sc_hd__buf_4
Xinput297 la_oenb_mprj[18] vssd vssd vccd vccd _515_/A sky130_fd_sc_hd__buf_4
XFILLER_48_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_587_ _587_/A _587_/B vssd vssd vccd vccd _587_/X sky130_fd_sc_hd__and2_2
XFILLER_32_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__B _436_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output494_A wire1282/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output661_A _031_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output759_A wire1180/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1292_A _371_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput705 _071_/Y vssd vssd vccd vccd la_data_in_mprj[88] sky130_fd_sc_hd__buf_8
Xoutput716 _081_/Y vssd vssd vccd vccd la_data_in_mprj[98] sky130_fd_sc_hd__buf_8
XFILLER_29_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput727 _604_/X vssd vssd vccd vccd la_oenb_core[107] sky130_fd_sc_hd__buf_8
Xoutput738 _614_/X vssd vssd vccd vccd la_oenb_core[117] sky130_fd_sc_hd__buf_8
XFILLER_42_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput749 wire1143/X vssd vssd vccd vccd la_oenb_core[127] sky130_fd_sc_hd__buf_8
XANTENNA_output926_A wire1334/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1557_A wire1558/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1724_A wire1725/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__346__B _346_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[93\]_B wire1466/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__362__A _362_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_518 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_510_ _510_/A _510_/B vssd vssd vccd vccd _510_/X sky130_fd_sc_hd__and2_4
XFILLER_22_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2078 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2038_A wire2039/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_441_ _569_/A _441_/B _441_/C vssd vssd vccd vccd _441_/X sky130_fd_sc_hd__and3b_4
XTAP_1912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__537__A _537_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_372_ _500_/A _372_/B _372_/C vssd vssd vccd vccd _372_/X sky130_fd_sc_hd__and3b_4
XTAP_1967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2205_A wire2205/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_4056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input392_A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2632 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[84\]_B wire1475/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input86_A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__272__A _272_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_934 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3451 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2811 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output507_A wire1270/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1040_A _130_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1305_A wire1306/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output876_A wire1424/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] _182_/X vssd vssd vccd vccd _002_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_32_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[75\]_B _238_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__182__A _182_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1674_A wire1674/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput502 wire1293/X vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__buf_8
XFILLER_44_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput513 wire1292/X vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__buf_8
XFILLER_48_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput524 wire1291/X vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__buf_8
XFILLER_9_2700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput535 wire1290/X vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__buf_8
XFILLER_9_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput546 wire1289/X vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__buf_8
XFILLER_44_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput557 wire1288/X vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__buf_8
XANTENNA_wire1841_A wire1842/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput568 wire1287/X vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__buf_8
XFILLER_47_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1939_A wire1939/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput579 wire1286/X vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__buf_8
XFILLER_5_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__357__A _357_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1806 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__092__A _092_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1800 wire1801/X vssd vssd vccd vccd _373_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input140_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1811 wire1811/A vssd vssd vccd vccd wire1811/X sky130_fd_sc_hd__buf_6
XFILLER_24_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1822 wire1823/X vssd vssd vccd vccd _363_/A sky130_fd_sc_hd__buf_6
XANTENNA_input238_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1833 wire1833/A vssd vssd vccd vccd _354_/A sky130_fd_sc_hd__buf_6
Xwire1844 wire1845/X vssd vssd vccd vccd _292_/A sky130_fd_sc_hd__buf_6
XFILLER_46_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1855 wire1855/A vssd vssd vccd vccd wire1855/X sky130_fd_sc_hd__buf_6
XTAP_3100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1866 wire1866/A vssd vssd vccd vccd wire1866/X sky130_fd_sc_hd__buf_6
XTAP_3122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1877 wire1878/X vssd vssd vccd vccd _280_/A sky130_fd_sc_hd__buf_6
XTAP_3133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1888 wire1888/A vssd vssd vccd vccd _272_/A sky130_fd_sc_hd__buf_6
XFILLER_41_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1899 wire1900/X vssd vssd vccd vccd _265_/A sky130_fd_sc_hd__buf_6
XTAP_3155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input405_A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_100 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__267__A _267_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _512_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_155 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _473_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_424_ _552_/A _424_/B _424_/C vssd vssd vccd vccd _424_/X sky130_fd_sc_hd__and3b_2
XTAP_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_177 wire995/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _340_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _355_/A _355_/B vssd vssd vccd vccd _355_/X sky130_fd_sc_hd__and2_4
XFILLER_50_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_B _220_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_286_ _286_/A _286_/B vssd vssd vccd vccd _286_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__433__C _433_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4247 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1088_A wire1089/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1255_A _407_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput6 la_data_out_mprj[101] vssd vssd vccd vccd _470_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1422_A _313_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__177__A _177_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1791_A wire1792/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[48\]_B _211_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1889_A wire1889/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__624__B _624_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] _625_/X vssd vssd vccd vccd _147_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_40_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1107 wire1108/X vssd vssd vccd vccd wire1107/X sky130_fd_sc_hd__buf_6
XFILLER_29_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1118 wire1119/X vssd vssd vccd vccd wire1118/X sky130_fd_sc_hd__buf_6
Xwire1129 wire1129/A vssd vssd vccd vccd _069_/A sky130_fd_sc_hd__buf_6
XFILLER_20_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__087__A _087_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[39\]_B _202_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_140_ _140_/A vssd vssd vccd vccd _140_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__534__B _534_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_B _286_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_071_ _071_/A vssd vssd vccd vccd _071_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_3369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2635 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input188_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__550__A _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input355_A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2272_A wire2272/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__A_N _590_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input49_A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1630 wire1631/X vssd vssd vccd vccd _327_/B sky130_fd_sc_hd__buf_6
Xwire1641 wire1642/X vssd vssd vccd vccd wire1641/X sky130_fd_sc_hd__buf_6
XFILLER_47_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1652 wire1653/X vssd vssd vccd vccd _322_/B sky130_fd_sc_hd__buf_6
XFILLER_19_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1663 wire1664/X vssd vssd vccd vccd _319_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1674 wire1674/A vssd vssd vccd vccd wire1674/X sky130_fd_sc_hd__buf_6
Xwire1685 wire1685/A vssd vssd vccd vccd _584_/A sky130_fd_sc_hd__buf_6
XFILLER_19_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1696 wire1696/A vssd vssd vccd vccd _573_/A sky130_fd_sc_hd__buf_8
XFILLER_34_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__428__C _428_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ _535_/A _407_/B _407_/C vssd vssd vccd vccd _407_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_3258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__444__B _444_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_B _277_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_338_ _338_/A _338_/B vssd vssd vccd vccd _338_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1003_A wire1004/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output574_A _454_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_269_ _269_/A _269_/B vssd vssd vccd vccd _269_/X sky130_fd_sc_hd__and2_2
Xwire971 wire972/X vssd vssd vccd vccd wire971/X sky130_fd_sc_hd__buf_6
XFILLER_48_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire982 wire983/X vssd vssd vccd vccd wire982/X sky130_fd_sc_hd__buf_6
Xwire993 wire994/X vssd vssd vccd vccd wire993/X sky130_fd_sc_hd__buf_6
XANTENNA_output741_A wire1189/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output839_A _590_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1372_A _346_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] wire1473/X vssd vssd vccd vccd wire1129/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_3387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1637_A wire1638/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3194 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__619__B _619_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1804_A wire1805/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[23\]_A mprj_dat_i_user[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire992_A wire993/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_11 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_22 _223_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_B wire1463/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__354__B _354_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_33 _361_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_44 _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_55 _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_66 _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_77 _288_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_88 _243_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_99 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__485__A_N _613_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2439 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3796 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_A mprj_dat_i_user[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2020_A wire2021/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input103_A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2118_A wire2118/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3567 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__545__A _545_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__264__B _264_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_123_ _123_/A vssd vssd vccd vccd _123_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_054_ _054_/A vssd vssd vccd vccd _054_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__280__A _280_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2150 wire2150/A vssd vssd vccd vccd wire2150/X sky130_fd_sc_hd__buf_6
XFILLER_1_4068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2161 wire2162/X vssd vssd vccd vccd _500_/B sky130_fd_sc_hd__buf_6
XFILLER_40_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2172 wire2173/X vssd vssd vccd vccd wire2172/X sky130_fd_sc_hd__buf_6
XFILLER_8_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2183 wire2184/X vssd vssd vccd vccd wire2183/X sky130_fd_sc_hd__buf_6
XFILLER_5_2780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2194 wire2195/X vssd vssd vccd vccd _487_/B sky130_fd_sc_hd__buf_6
XFILLER_19_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1460 wire1461/X vssd vssd vccd vccd wire1460/X sky130_fd_sc_hd__buf_8
XFILLER_1_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__439__B _439_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1471 _251_/X vssd vssd vccd vccd wire1471/X sky130_fd_sc_hd__buf_6
XFILLER_1_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1482 _240_/X vssd vssd vccd vccd wire1482/X sky130_fd_sc_hd__buf_6
XFILLER_21_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1493 wire1493/A vssd vssd vccd vccd wire1493/X sky130_fd_sc_hd__buf_6
XFILLER_1_2666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1120_A _114_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1218_A _464_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output691_A _058_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output789_A _545_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__174__B _174_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output956_A _297_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] split4/X vssd vssd vccd vccd _128_/A
+ sky130_fd_sc_hd__nand2_8
Xinput20 la_data_out_mprj[114] vssd vssd vccd vccd input20/X sky130_fd_sc_hd__buf_6
XFILLER_28_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput31 la_data_out_mprj[124] vssd vssd vccd vccd _493_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1587_A wire1588/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput42 la_data_out_mprj[19] vssd vssd vccd vccd _388_/C sky130_fd_sc_hd__clkbuf_4
Xinput53 la_data_out_mprj[29] vssd vssd vccd vccd _398_/C sky130_fd_sc_hd__clkbuf_4
Xinput64 la_data_out_mprj[39] vssd vssd vccd vccd _408_/C sky130_fd_sc_hd__clkbuf_4
Xinput75 la_data_out_mprj[49] vssd vssd vccd vccd _418_/C sky130_fd_sc_hd__clkbuf_4
Xinput86 la_data_out_mprj[59] vssd vssd vccd vccd _428_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__A _190_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput97 la_data_out_mprj[69] vssd vssd vccd vccd input97/X sky130_fd_sc_hd__buf_6
XFILLER_44_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] _275_/X vssd vssd vccd vccd _095_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA__349__B _349_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__365__A _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1016 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput402 mprj_adr_o_core[22] vssd vssd vccd vccd wire1632/A sky130_fd_sc_hd__buf_6
XFILLER_2_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput413 mprj_adr_o_core[3] vssd vssd vccd vccd wire1581/A sky130_fd_sc_hd__buf_6
XANTENNA_wire2068_A wire2069/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput424 mprj_dat_o_core[12] vssd vssd vccd vccd wire1541/A sky130_fd_sc_hd__buf_6
Xinput435 mprj_dat_o_core[22] vssd vssd vccd vccd wire1522/A sky130_fd_sc_hd__buf_6
XFILLER_0_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput446 mprj_dat_o_core[3] vssd vssd vccd vccd wire1510/A sky130_fd_sc_hd__buf_6
XFILLER_5_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput457 mprj_sel_o_core[3] vssd vssd vccd vccd _304_/B sky130_fd_sc_hd__buf_4
XFILLER_2_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input220_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input318_A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__275__A _275_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3206 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2554 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_106_ _106_/A vssd vssd vccd vccd _106_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput909 wire1086/X vssd vssd vccd vccd mprj_dat_i_core[6] sky130_fd_sc_hd__buf_8
X_037_ _037_/A vssd vssd vccd vccd _037_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__441__C _441_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output537_A wire1242/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1070_A _124_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1335_A wire1336/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1290 _373_/X vssd vssd vccd vccd wire1290/X sky130_fd_sc_hd__buf_6
XFILLER_39_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] _212_/X vssd vssd vccd vccd _032_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_35_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1502_A wire1502/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__185__A _185_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3762 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1871_A wire1872/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1969_A wire1969/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2628 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3640 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3531 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__095__A _095_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__542__B _542_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input170_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input268_A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2185_A wire2186/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input435_A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput210 la_iena_mprj[55] vssd vssd vccd vccd _218_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input31_A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput221 la_iena_mprj[65] vssd vssd vccd vccd _228_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput232 la_iena_mprj[75] vssd vssd vccd vccd _238_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput243 la_iena_mprj[85] vssd vssd vccd vccd _248_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput254 la_iena_mprj[95] vssd vssd vccd vccd _258_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput265 la_oenb_mprj[104] vssd vssd vccd vccd _601_/A sky130_fd_sc_hd__buf_4
XFILLER_48_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput276 la_oenb_mprj[114] vssd vssd vccd vccd wire1733/A sky130_fd_sc_hd__buf_6
Xinput287 la_oenb_mprj[124] vssd vssd vccd vccd _621_/A sky130_fd_sc_hd__buf_4
XFILLER_18_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput298 la_oenb_mprj[19] vssd vssd vccd vccd _516_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_586_ _586_/A _586_/B vssd vssd vccd vccd _586_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__C _436_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output487_A _490_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__452__B _452_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output654_A _024_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput706 _072_/Y vssd vssd vccd vccd la_data_in_mprj[89] sky130_fd_sc_hd__buf_8
Xoutput717 _082_/Y vssd vssd vccd vccd la_data_in_mprj[99] sky130_fd_sc_hd__buf_8
XFILLER_29_2821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput728 _605_/X vssd vssd vccd vccd la_oenb_core[108] sky130_fd_sc_hd__buf_8
XFILLER_25_3419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1285_A _378_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput739 _615_/X vssd vssd vccd vccd la_oenb_core[118] sky130_fd_sc_hd__buf_8
XFILLER_42_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output821_A _574_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output919_A wire1352/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3226 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1717_A _405_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__362__B _362_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1734 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[6\]_A mprj_dat_i_user[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_440_ _568_/A _440_/B _440_/C vssd vssd vccd vccd _440_/X sky130_fd_sc_hd__and3b_4
XTAP_2658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__419__A_N _547_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_371_ _499_/A _371_/B _371_/C vssd vssd vccd vccd _371_/X sky130_fd_sc_hd__and3b_4
XTAP_1957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4068 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2100_A wire2100/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__553__A _553_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input385_A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input79_A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4028 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3463 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__447__B _447_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1033_A wire1034/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_569_ _569_/A _569_/B vssd vssd vccd vccd _569_/X sky130_fd_sc_hd__and2_4
XFILLER_31_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1200_A _497_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output771_A _528_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output869_A _334_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__182__B _182_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput503 wire1274/X vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__buf_8
Xoutput514 wire1263/X vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__buf_8
XFILLER_44_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1667_A wire1667/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput525 wire1253/X vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__buf_8
XFILLER_48_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput536 wire1243/X vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__buf_8
XFILLER_47_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput547 wire1227/X vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__buf_8
XFILLER_42_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput558 _439_/X vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__buf_8
Xoutput569 _449_/X vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__buf_8
XFILLER_47_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__357__B _357_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1239 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2222 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3980 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3783 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1801 wire1801/A vssd vssd vccd vccd wire1801/X sky130_fd_sc_hd__buf_6
XFILLER_41_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1812 wire1813/X vssd vssd vccd vccd _367_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1823 wire1823/A vssd vssd vccd vccd wire1823/X sky130_fd_sc_hd__buf_6
Xwire1834 wire1834/A vssd vssd vccd vccd _353_/A sky130_fd_sc_hd__buf_6
XFILLER_19_817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1845 wire1846/X vssd vssd vccd vccd wire1845/X sky130_fd_sc_hd__buf_6
XANTENNA_input133_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2050_A wire2051/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1856 wire1857/X vssd vssd vccd vccd _288_/A sky130_fd_sc_hd__buf_6
XTAP_3101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1867 wire1868/X vssd vssd vccd vccd _284_/A sky130_fd_sc_hd__buf_6
XFILLER_45_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__548__A _548_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1878 wire1878/A vssd vssd vccd vccd wire1878/X sky130_fd_sc_hd__buf_6
XTAP_3134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1889 wire1889/A vssd vssd vccd vccd _271_/A sky130_fd_sc_hd__buf_6
XTAP_3145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_101 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_112 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input300_A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_123 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__267__B _267_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1718 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_167 _465_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_423_ _551_/A _423_/B _423_/C vssd vssd vccd vccd _423_/X sky130_fd_sc_hd__and3b_2
XFILLER_35_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_178 wire1094/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__391__A_N _519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_189 _343_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_354_ _354_/A _354_/B vssd vssd vccd vccd _354_/X sky130_fd_sc_hd__and2_4
XTAP_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__283__A _283_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_285_ _285_/A _285_/B vssd vssd vccd vccd _285_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4215 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output617_A _106_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1150_A wire1151/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2592 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1248_A _414_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput7 la_data_out_mprj[102] vssd vssd vccd vccd _471_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__177__B _177_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1415_A wire1416/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] _194_/X vssd vssd vccd vccd _014_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_138 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__193__A _193_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1784_A wire1785/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1951_A wire1951/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1108 wire1109/X vssd vssd vccd vccd wire1108/X sky130_fd_sc_hd__buf_6
XFILLER_5_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1119 wire1120/X vssd vssd vccd vccd wire1119/X sky130_fd_sc_hd__buf_6
XFILLER_9_1874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__368__A _368_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_070_ _070_/A vssd vssd vccd vccd _070_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1924 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2098_A wire2098/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__550__B _550_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input250_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2265_A wire2266/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input348_A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1620 wire1621/X vssd vssd vccd vccd wire1620/X sky130_fd_sc_hd__buf_6
XFILLER_8_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1631 wire1632/X vssd vssd vccd vccd wire1631/X sky130_fd_sc_hd__buf_6
Xwire1642 wire1643/X vssd vssd vccd vccd wire1642/X sky130_fd_sc_hd__buf_6
Xwire1653 wire1654/X vssd vssd vccd vccd wire1653/X sky130_fd_sc_hd__buf_6
XFILLER_5_2984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1664 wire1665/X vssd vssd vccd vccd wire1664/X sky130_fd_sc_hd__buf_6
XFILLER_20_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__278__A _278_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1675 wire1676/X vssd vssd vccd vccd _305_/B sky130_fd_sc_hd__buf_6
XFILLER_46_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1686 wire1686/A vssd vssd vccd vccd _583_/A sky130_fd_sc_hd__buf_6
Xwire1697 wire1697/A vssd vssd vccd vccd _572_/A sky130_fd_sc_hd__buf_8
XFILLER_19_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_406_ _406_/A_N _406_/B _406_/C vssd vssd vccd vccd _406_/X sky130_fd_sc_hd__and3b_4
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_337_ _337_/A _337_/B vssd vssd vccd vccd _337_/X sky130_fd_sc_hd__and2_2
XANTENNA__444__C _444_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_268_ _268_/A _268_/B vssd vssd vccd vccd _268_/X sky130_fd_sc_hd__and2_2
XANTENNA_output567_A _448_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire961 wire962/X vssd vssd vccd vccd wire961/X sky130_fd_sc_hd__buf_6
XFILLER_28_3609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire972 wire973/X vssd vssd vccd vccd wire972/X sky130_fd_sc_hd__buf_6
XFILLER_45_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire983 wire984/X vssd vssd vccd vccd wire983/X sky130_fd_sc_hd__buf_6
XFILLER_31_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire994 wire995/X vssd vssd vccd vccd wire994/X sky130_fd_sc_hd__buf_6
X_199_ _199_/A _199_/B vssd vssd vccd vccd _199_/X sky130_fd_sc_hd__and2_2
XFILLER_6_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1198_A _499_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__460__B _460_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4067 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output734_A _610_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1365_A wire1366/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_790 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output901_A wire978/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] wire1480/X vssd vssd vccd vccd wire1136/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_46_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1532_A wire1533/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__188__A _188_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1999_A wire2000/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire985_A wire986/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_12 _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_23 _285_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_34 _361_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_45 _618_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_56 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_67 _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_78 _288_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_89 _243_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__370__B _370_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__098__A _098_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_B split4/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2013_A wire2014/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input298_A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_122_ _122_/A vssd vssd vccd vccd _122_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_3145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__561__A _561_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_053_ _053_/A vssd vssd vccd vccd _053_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_27_4343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input61_A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2140 wire2140/A vssd vssd vccd vccd _518_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2151 wire2151/A vssd vssd vccd vccd _508_/B sky130_fd_sc_hd__buf_6
XFILLER_43_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2162 wire2162/A vssd vssd vccd vccd wire2162/X sky130_fd_sc_hd__buf_6
Xwire2173 wire2173/A vssd vssd vccd vccd wire2173/X sky130_fd_sc_hd__buf_6
XFILLER_5_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2184 wire2184/A vssd vssd vccd vccd wire2184/X sky130_fd_sc_hd__buf_6
Xwire1450 wire1451/X vssd vssd vccd vccd wire1450/X sky130_fd_sc_hd__buf_6
Xwire2195 wire2196/X vssd vssd vccd vccd wire2195/X sky130_fd_sc_hd__buf_6
XFILLER_5_2792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1461 _294_/X vssd vssd vccd vccd wire1461/X sky130_fd_sc_hd__buf_6
XFILLER_47_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1472 _250_/X vssd vssd vccd vccd wire1472/X sky130_fd_sc_hd__buf_6
XANTENNA__439__C _439_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1483 input99/X vssd vssd vccd vccd _439_/C sky130_fd_sc_hd__buf_6
XFILLER_47_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1494 wire1495/X vssd vssd vccd vccd _294_/B sky130_fd_sc_hd__buf_6
XFILLER_35_926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__455__B _455_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1113_A wire1114/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output684_A _052_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput10 la_data_out_mprj[105] vssd vssd vccd vccd _474_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output851_A wire1412/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput21 la_data_out_mprj[115] vssd vssd vccd vccd input21/X sky130_fd_sc_hd__buf_6
XFILLER_28_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput32 la_data_out_mprj[125] vssd vssd vccd vccd _494_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output949_A wire1449/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput43 la_data_out_mprj[1] vssd vssd vccd vccd _370_/C sky130_fd_sc_hd__clkbuf_4
Xinput54 la_data_out_mprj[2] vssd vssd vccd vccd _371_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput65 la_data_out_mprj[3] vssd vssd vccd vccd _372_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1482_A _240_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput76 la_data_out_mprj[4] vssd vssd vccd vccd _373_/C sky130_fd_sc_hd__clkbuf_4
Xinput87 la_data_out_mprj[5] vssd vssd vccd vccd _374_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__B _190_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput98 la_data_out_mprj[6] vssd vssd vccd vccd _375_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1747_A wire1747/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1719 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] wire1463/X vssd vssd vccd vccd
+ _088_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_2144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj2_logic_high_inst wire2306/A vccd2_uq0 vssd2_uq0 mprj2_logic_high
XFILLER_11_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__365__B _365_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__452__A_N _580_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_4301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2259 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput403 mprj_adr_o_core[23] vssd vssd vccd vccd wire1629/A sky130_fd_sc_hd__buf_6
XFILLER_44_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput414 mprj_adr_o_core[4] vssd vssd vccd vccd wire1576/A sky130_fd_sc_hd__buf_6
XFILLER_22_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput425 mprj_dat_o_core[13] vssd vssd vccd vccd wire1539/A sky130_fd_sc_hd__buf_6
XFILLER_6_3791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput436 mprj_dat_o_core[23] vssd vssd vccd vccd wire1521/A sky130_fd_sc_hd__buf_6
XFILLER_40_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput447 mprj_dat_o_core[4] vssd vssd vccd vccd wire1508/A sky130_fd_sc_hd__buf_6
Xinput458 mprj_stb_o_core vssd vssd vccd vccd wire1493/A sky130_fd_sc_hd__buf_6
XFILLER_5_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2130_A wire2130/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input213_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2228_A wire2229/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__556__A _556_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__275__B _275_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__291__A _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_105_ _105_/A vssd vssd vccd vccd _105_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_036_ _036_/A vssd vssd vccd vccd _036_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1063_A wire1064/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1280 _383_/X vssd vssd vccd vccd wire1280/X sky130_fd_sc_hd__buf_6
Xwire1291 _372_/X vssd vssd vccd vccd wire1291/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1328_A wire1329/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__475__A_N _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output899_A wire987/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__185__B _185_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1864_A wire1865/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1906 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xmprj_logic_high_inst wire2301/A wire2300/A _396_/B _397_/B _398_/B _399_/B _400_/B
+ _401_/B _402_/B _403_/B _404_/B wire2299/A _405_/B _406_/B _407_/B _408_/B _409_/B
+ _410_/B _411_/B _412_/B _413_/B _414_/B wire2298/A _415_/B _416_/B _417_/B _418_/B
+ _419_/B _420_/B _421_/B _422_/B _423_/B _424_/B wire2297/A _425_/B _426_/B _427_/B
+ _428_/B _429_/B _430_/B _431_/B wire2296/A wire2295/A wire2294/A wire2293/A wire2292/A
+ wire2291/A wire2290/A wire2288/A wire2287/A wire2286/A wire2285/A wire2284/A wire2283/A
+ wire2282/A wire2281/A wire2280/A wire2279/A wire2278/A wire2277/A wire2276/A wire2274/A
+ wire2272/A wire2270/A wire2267/A wire2264/A wire2261/A wire2260/A wire2257/A wire2254/A
+ wire2251/A wire2250/A wire2249/A wire2248/A wire2247/A wire2246/A wire2245/A _311_/A
+ wire2244/A wire2243/A wire2241/A wire2239/A wire2238/A wire2236/A wire2235/A wire2233/A
+ wire2231/A wire2229/A _312_/A wire2227/A wire2225/A wire2223/A wire2221/A wire2219/A
+ wire2217/A wire2214/A wire2211/A wire2208/A wire2205/A _313_/A wire2202/A wire2199/A
+ wire2196/A wire2193/A wire2190/A wire2187/A wire2184/A wire2181/A wire2178/A wire2175/A
+ _314_/A _296_/A wire2173/A wire2170/A wire2168/A wire2166/A wire2164/A wire2162/A
+ wire2160/A wire2159/A wire2157/A wire2156/A _315_/A wire2155/A wire2154/A wire2152/A
+ wire2151/A _509_/B wire2150/A wire2148/A wire2146/A wire2145/A wire2144/A _316_/A
+ wire2143/A wire2142/A wire2141/A wire2140/A wire2139/A wire2138/A wire2137/A wire2136/A
+ _523_/B _524_/B _317_/A wire2135/A _526_/B _527_/B _528_/B _529_/B wire2134/A wire2133/A
+ _532_/B _533_/B _534_/B _318_/A _535_/B _536_/B _537_/B wire2132/A _539_/B _540_/B
+ _541_/B _542_/B _543_/B _544_/B _319_/A _545_/B _546_/B _547_/B _548_/B _549_/B
+ _550_/B _551_/B _552_/B _553_/B _554_/B _320_/A _555_/B _556_/B _557_/B _558_/B
+ wire2131/A _560_/B wire2130/A wire2129/A wire2128/A wire2127/A _321_/A wire2126/A
+ wire2125/A wire2123/A wire2122/A wire2120/A wire2118/A wire2117/A wire2116/A wire2114/A
+ wire2112/A _322_/A wire2110/A wire2108/A wire2106/A wire2104/A wire2102/A wire2100/A
+ wire2098/A wire2096/A wire2094/A wire2091/A _323_/A wire2089/A wire2087/A wire2086/A
+ wire2085/A wire2083/A wire2082/A wire2081/A wire2079/A wire2077/A wire2075/A _324_/A
+ wire2073/A wire2069/A wire2067/A wire2065/A wire2063/A wire2061/A wire2059/A wire2057/A
+ wire2055/A wire2053/A wire2051/A _325_/A wire2049/A wire2046/A wire2044/A wire2041/A
+ wire2039/A wire2037/A wire2034/A wire2031/A wire2028/A wire2025/A _326_/A wire2022/A
+ wire2019/A wire2015/A wire2012/A wire2009/A wire2006/A wire2003/A wire2000/A wire1997/A
+ wire1994/A _327_/A wire1991/A wire1989/A wire1987/A wire1985/A wire1983/A wire1981/A
+ wire1979/A wire1978/A wire1976/A wire1975/A _328_/A wire1974/A wire1973/A wire1971/A
+ wire1969/A wire1967/A wire1966/A wire1964/A wire1962/A wire1961/A wire1960/A wire1958/A
+ wire1957/A wire1955/A wire1953/A wire1952/A wire1951/A wire1950/A wire1949/A wire1948/A
+ wire1947/A wire1945/A wire1944/A wire1943/A wire1942/A wire1941/A wire1940/A _197_/A
+ _198_/A _199_/A _200_/A _201_/A _202_/A wire1939/A _203_/A _204_/A _205_/A _206_/A
+ wire1938/A wire1937/A wire1936/A _210_/A _211_/A _212_/A wire1935/A _213_/A _214_/A
+ _215_/A _216_/A _217_/A _218_/A _219_/A _220_/A _221_/A _222_/A wire1934/A _223_/A
+ _224_/A _225_/A _226_/A _227_/A _228_/A _229_/A wire1933/A wire1932/A wire1931/A
+ wire1930/A wire1929/A wire1928/A wire1927/A _235_/A _236_/A _237_/A wire1926/A _239_/A
+ _240_/A _241_/A wire1925/A wire1924/A wire1923/A _244_/A _245_/A _246_/A _247_/A
+ wire1922/A wire1921/A wire1920/A wire1919/A wire1918/A _336_/A wire1917/A wire1916/A
+ wire1915/A wire1914/A wire1913/A wire1912/A wire1911/A wire1910/A wire1908/A wire1906/A
+ _337_/A wire1904/A wire1902/A wire1900/A wire1898/A wire1896/A wire1894/A wire1892/A
+ wire1890/A wire1889/A wire1888/A _338_/A wire1887/A wire1886/A wire1885/A wire1884/A
+ wire1883/A wire1882/A wire1880/A wire1878/A wire1876/A wire1874/A _339_/A wire1872/A
+ wire1869/A wire1866/A wire1863/A wire1860/A wire1858/A wire1855/A wire1852/A wire1849/A
+ wire1846/A _340_/A wire1843/A wire1840/A _294_/A _341_/A _342_/A _343_/A _344_/A
+ _299_/A _345_/A _346_/A _347_/A _348_/A _349_/A wire1837/A wire1836/A wire1835/A
+ wire1834/A wire1833/A wire1832/A wire1831/A wire1830/A wire1829/A wire1828/A wire1827/A
+ wire1826/A wire1825/A wire1824/A wire1823/A wire1821/A wire1819/A wire1817/A wire1815/A
+ wire1813/A wire1811/A wire1809/A wire1807/A wire1805/A wire1803/A wire1801/A wire1799/A
+ wire1797/A wire1795/A wire1792/A wire1789/A wire1787/A wire1785/A wire1783/A wire1781/A
+ wire1779/A wire1777/A wire1775/A wire1773/A wire1771/A wire1769/A wire1767/A wire1765/A
+ wire1763/A wire1761/A wire1760/A wire1759/A wire1758/A wire1757/A wire1755/A vccd1_uq1
+ vssd1_uq1 mprj_logic_high
XTAP_3508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_962 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2080_A wire2081/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input163_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2178_A wire2178/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput200 la_iena_mprj[46] vssd vssd vccd vccd _209_/B sky130_fd_sc_hd__buf_4
XFILLER_24_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput211 la_iena_mprj[56] vssd vssd vccd vccd _219_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput222 la_iena_mprj[66] vssd vssd vccd vccd _229_/B sky130_fd_sc_hd__buf_4
XFILLER_0_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput233 la_iena_mprj[76] vssd vssd vccd vccd _239_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input330_A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput244 la_iena_mprj[86] vssd vssd vccd vccd _249_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_input428_A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput255 la_iena_mprj[96] vssd vssd vccd vccd _259_/B sky130_fd_sc_hd__clkbuf_4
Xinput266 la_oenb_mprj[105] vssd vssd vccd vccd _602_/A sky130_fd_sc_hd__buf_4
XANTENNA_input24_A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput277 la_oenb_mprj[115] vssd vssd vccd vccd wire1732/A sky130_fd_sc_hd__buf_6
XFILLER_40_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput288 la_oenb_mprj[125] vssd vssd vccd vccd _622_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_2740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput299 la_oenb_mprj[1] vssd vssd vccd vccd _498_/A sky130_fd_sc_hd__buf_4
XFILLER_29_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__286__A _286_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_585_ _585_/A _585_/B vssd vssd vccd vccd _585_/X sky130_fd_sc_hd__and2_4
XFILLER_17_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__452__C _452_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput707 _155_/Y vssd vssd vccd vccd la_data_in_mprj[8] sky130_fd_sc_hd__buf_8
Xoutput718 _156_/Y vssd vssd vccd vccd la_data_in_mprj[9] sky130_fd_sc_hd__buf_8
Xoutput729 _606_/X vssd vssd vccd vccd la_oenb_core[109] sky130_fd_sc_hd__buf_8
X_019_ _019_/A vssd vssd vccd vccd _019_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_29_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1180_A _517_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1278_A _385_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1445_A wire1446/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1961 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] _224_/X vssd vssd vccd vccd _044_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_3_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1612_A wire1613/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__196__A _196_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[6\]_B split4/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1747 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _498_/A _370_/B _370_/C vssd vssd vccd vccd _370_/X sky130_fd_sc_hd__and3b_4
XTAP_1947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__553__B _553_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input280_A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2295_A wire2295/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input378_A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__447__C _447_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_568_ _568_/A _568_/B vssd vssd vccd vccd _568_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1026_A wire1027/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output597_A _088_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_499_ _499_/A _499_/B vssd vssd vccd vccd _499_/X sky130_fd_sc_hd__and2_4
XFILLER_32_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__B _463_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output764_A wire1175/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1395_A wire1396/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput504 wire1273/X vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__buf_8
XANTENNA_output931_A wire1315/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput515 wire1262/X vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__buf_8
XFILLER_44_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput526 wire1252/X vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__buf_8
Xoutput537 wire1242/X vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__buf_8
Xoutput548 wire1226/X vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__buf_8
XANTENNA_wire1562_A wire1563/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput559 _440_/X vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__buf_8
XFILLER_42_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1827_A wire1827/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__373__B _373_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2234 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1802 wire1803/X vssd vssd vccd vccd _372_/B sky130_fd_sc_hd__buf_6
Xwire1813 wire1813/A vssd vssd vccd vccd wire1813/X sky130_fd_sc_hd__buf_6
Xwire1824 wire1824/A vssd vssd vccd vccd _362_/A sky130_fd_sc_hd__buf_6
XFILLER_43_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1835 wire1835/A vssd vssd vccd vccd _352_/A sky130_fd_sc_hd__buf_6
Xwire1846 wire1846/A vssd vssd vccd vccd wire1846/X sky130_fd_sc_hd__buf_6
XTAP_3102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1857 wire1858/X vssd vssd vccd vccd wire1857/X sky130_fd_sc_hd__buf_6
XTAP_3113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1868 wire1869/X vssd vssd vccd vccd wire1868/X sky130_fd_sc_hd__buf_6
XFILLER_41_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1879 wire1880/X vssd vssd vccd vccd _279_/A sky130_fd_sc_hd__buf_6
XFILLER_46_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__548__B _548_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2043_A wire2044/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input126_A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_113 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_146 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 wire2208/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_422_ _550_/A _422_/B _422_/C vssd vssd vccd vccd _422_/X sky130_fd_sc_hd__and3b_2
XTAP_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2210_A wire2211/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _465_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_179 wire1107/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__564__A _564_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ _353_/A _353_/B vssd vssd vccd vccd _353_/X sky130_fd_sc_hd__and2_4
XTAP_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__283__B _283_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input91_A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_284_ _284_/A _284_/B vssd vssd vccd vccd _284_/X sky130_fd_sc_hd__and2_4
XFILLER_52_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] rebuffer1/X vssd vssd vccd vccd _121_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_26_4227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2908 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2858 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output512_A wire1264/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput8 la_data_out_mprj[103] vssd vssd vccd vccd _472_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__458__B _458_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1143_A _624_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1310_A _365_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1408_A wire1409/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output881_A wire1116/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] _187_/X vssd vssd vccd vccd _007_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__193__B _193_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1777_A wire1777/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1944_A wire1944/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__409__A_N _409_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1109 wire1110/X vssd vssd vccd vccd wire1109/X sky130_fd_sc_hd__buf_6
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__368__B _368_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3692 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_14_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2300 wire2300/A vssd vssd vccd vccd _395_/B sky130_fd_sc_hd__buf_6
Xoutput890 wire1026/X vssd vssd vccd vccd mprj_dat_i_core[18] sky130_fd_sc_hd__buf_8
XFILLER_43_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2160_A wire2160/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input243_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4168 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2258_A wire2259/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1610 wire1611/X vssd vssd vccd vccd wire1610/X sky130_fd_sc_hd__buf_6
XANTENNA__559__A _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1621 wire1621/A vssd vssd vccd vccd wire1621/X sky130_fd_sc_hd__buf_6
XFILLER_24_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1632 wire1632/A vssd vssd vccd vccd wire1632/X sky130_fd_sc_hd__buf_6
Xwire1643 wire1644/X vssd vssd vccd vccd wire1643/X sky130_fd_sc_hd__buf_6
XFILLER_8_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1654 wire1654/A vssd vssd vccd vccd wire1654/X sky130_fd_sc_hd__buf_6
XFILLER_19_4020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1665 wire1665/A vssd vssd vccd vccd wire1665/X sky130_fd_sc_hd__buf_6
XANTENNA_input410_A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1676 wire1677/X vssd vssd vccd vccd wire1676/X sky130_fd_sc_hd__buf_6
XFILLER_46_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1687 wire1687/A vssd vssd vccd vccd _582_/A sky130_fd_sc_hd__buf_6
Xwire1698 wire1698/A vssd vssd vccd vccd _571_/A sky130_fd_sc_hd__buf_8
XFILLER_18_147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ _405_/A_N _405_/B _405_/C vssd vssd vccd vccd _405_/X sky130_fd_sc_hd__and3b_4
XANTENNA__294__A _294_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_336_ _336_/A _336_/B vssd vssd vccd vccd _336_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_267_ _267_/A _267_/B vssd vssd vccd vccd _267_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire962 wire963/X vssd vssd vccd vccd wire962/X sky130_fd_sc_hd__buf_6
Xwire973 _144_/Y vssd vssd vccd vccd wire973/X sky130_fd_sc_hd__buf_6
Xwire984 wire985/X vssd vssd vccd vccd wire984/X sky130_fd_sc_hd__buf_6
X_198_ _198_/A _198_/B vssd vssd vccd vccd _198_/X sky130_fd_sc_hd__and2_2
XFILLER_45_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire995 wire996/X vssd vssd vccd vccd wire995/X sky130_fd_sc_hd__buf_6
XFILLER_26_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1093_A wire1094/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4079 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output727_A _604_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1358_A wire1359/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__188__B _188_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1525_A wire1526/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_13 _219_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire978_A wire979/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_24 _290_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_35 _361_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_46 _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_57 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_68 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_79 _288_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1379 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__C _370_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__381__A_N _509_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2006_A wire2006/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_121_ _121_/A vssd vssd vccd vccd _121_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input193_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_052_ _052_/A vssd vssd vccd vccd _052_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__561__B _561_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input360_A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input458_A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input54_A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3220 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2130 wire2130/A vssd vssd vccd vccd _561_/B sky130_fd_sc_hd__buf_6
Xwire2141 wire2141/A vssd vssd vccd vccd _517_/B sky130_fd_sc_hd__buf_6
XANTENNA__289__A _289_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2152 wire2152/A vssd vssd vccd vccd _507_/B sky130_fd_sc_hd__buf_6
XFILLER_38_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2163 wire2164/X vssd vssd vccd vccd _499_/B sky130_fd_sc_hd__buf_6
Xwire2174 wire2175/X vssd vssd vccd vccd _494_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1440 wire1441/X vssd vssd vccd vccd wire1440/X sky130_fd_sc_hd__buf_8
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2185 wire2186/X vssd vssd vccd vccd _490_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2196 wire2196/A vssd vssd vccd vccd wire2196/X sky130_fd_sc_hd__buf_6
Xwire1451 _299_/X vssd vssd vccd vccd wire1451/X sky130_fd_sc_hd__buf_6
XFILLER_4_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1462 _269_/X vssd vssd vccd vccd wire1462/X sky130_fd_sc_hd__buf_8
XFILLER_38_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1473 _249_/X vssd vssd vccd vccd wire1473/X sky130_fd_sc_hd__buf_8
Xwire1484 input97/X vssd vssd vccd vccd _438_/C sky130_fd_sc_hd__buf_6
XFILLER_46_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1495 wire1496/X vssd vssd vccd vccd wire1495/X sky130_fd_sc_hd__buf_6
Xpowergood_check vccd vssd vdda1_uq0 vssa1_uq0 vdda2_uq0 vssa2_uq0 output954/A output952/A
+ mgmt_protect_hv
XFILLER_19_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__455__C _455_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1106_A wire1107/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_319_ _319_/A _319_/B vssd vssd vccd vccd _319_/X sky130_fd_sc_hd__and2_2
XFILLER_50_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput11 la_data_out_mprj[106] vssd vssd vccd vccd _475_/C sky130_fd_sc_hd__clkbuf_4
Xinput22 la_data_out_mprj[116] vssd vssd vccd vccd input22/X sky130_fd_sc_hd__buf_6
XFILLER_30_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput33 la_data_out_mprj[126] vssd vssd vccd vccd _495_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__471__B _471_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput44 la_data_out_mprj[20] vssd vssd vccd vccd _389_/C sky130_fd_sc_hd__clkbuf_4
Xinput55 la_data_out_mprj[30] vssd vssd vccd vccd _399_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output844_A _595_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput66 la_data_out_mprj[40] vssd vssd vccd vccd _409_/C sky130_fd_sc_hd__clkbuf_4
Xinput77 la_data_out_mprj[50] vssd vssd vccd vccd _419_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput88 la_data_out_mprj[60] vssd vssd vccd vccd _429_/C sky130_fd_sc_hd__clkbuf_4
Xinput99 la_data_out_mprj[70] vssd vssd vccd vccd input99/X sky130_fd_sc_hd__buf_6
XFILLER_28_2717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1475_A _247_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] wire1468/X vssd vssd vccd vccd wire1126/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_6_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1642_A wire1643/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__199__A _199_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1907_A wire1908/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3725 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__381__B _381_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4252 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput404 mprj_adr_o_core[24] vssd vssd vccd vccd wire1626/A sky130_fd_sc_hd__buf_6
XFILLER_40_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput415 mprj_adr_o_core[5] vssd vssd vccd vccd wire1571/A sky130_fd_sc_hd__buf_6
XFILLER_44_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput426 mprj_dat_o_core[14] vssd vssd vccd vccd wire1537/A sky130_fd_sc_hd__buf_6
XFILLER_6_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput437 mprj_dat_o_core[24] vssd vssd vccd vccd wire1520/A sky130_fd_sc_hd__buf_6
XFILLER_40_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput448 mprj_dat_o_core[5] vssd vssd vccd vccd wire1506/A sky130_fd_sc_hd__buf_6
XFILLER_22_3573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput459 mprj_we_o_core vssd vssd vccd vccd wire1491/A sky130_fd_sc_hd__buf_6
XFILLER_22_3584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__556__B _556_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2123_A wire2123/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input206_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__572__A _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_104_ _104_/A vssd vssd vccd vccd _104_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_8_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__291__B _291_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_035_ _035_/A vssd vssd vccd vccd _035_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4163 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1056_A wire1057/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1270 _393_/X vssd vssd vccd vccd wire1270/X sky130_fd_sc_hd__buf_6
Xwire1281 _382_/X vssd vssd vccd vccd wire1281/X sky130_fd_sc_hd__buf_6
XFILLER_1_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1292 _371_/X vssd vssd vccd vccd wire1292/X sky130_fd_sc_hd__buf_6
XFILLER_1_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__466__B _466_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1223_A _459_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output794_A wire1158/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1592_A wire1593/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1857_A wire1858/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__376__B _376_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B wire1464/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2073_A wire2073/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input156_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput201 la_iena_mprj[47] vssd vssd vccd vccd _210_/B sky130_fd_sc_hd__buf_4
XFILLER_2_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput212 la_iena_mprj[57] vssd vssd vccd vccd _220_/B sky130_fd_sc_hd__clkbuf_4
Xinput223 la_iena_mprj[67] vssd vssd vccd vccd _230_/B sky130_fd_sc_hd__buf_4
XTAP_4700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput234 la_iena_mprj[77] vssd vssd vccd vccd _240_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 la_iena_mprj[87] vssd vssd vccd vccd _250_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput256 la_iena_mprj[97] vssd vssd vccd vccd _260_/B sky130_fd_sc_hd__clkbuf_4
Xinput267 la_oenb_mprj[106] vssd vssd vccd vccd _603_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_input323_A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2240_A wire2241/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput278 la_oenb_mprj[116] vssd vssd vccd vccd wire1731/A sky130_fd_sc_hd__buf_6
Xinput289 la_oenb_mprj[126] vssd vssd vccd vccd _623_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__567__A _567_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input17_A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__286__B _286_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_584_ _584_/A _584_/B vssd vssd vccd vccd _584_/X sky130_fd_sc_hd__and2_4
XFILLER_38_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[87\]_B wire1472/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput708 _073_/Y vssd vssd vccd vccd la_data_in_mprj[90] sky130_fd_sc_hd__buf_8
Xoutput719 wire1200/X vssd vssd vccd vccd la_oenb_core[0] sky130_fd_sc_hd__buf_8
X_018_ _018_/A vssd vssd vccd vccd _018_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output542_A wire1232/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1173_A _525_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[11\]_B _174_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__442__A_N _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output807_A _561_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1340_A wire1341/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1438_A wire1439/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] _217_/X vssd vssd vccd vccd _037_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA__196__B _196_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1605_A wire1606/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[78\]_B wire1481/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1974_A wire1974/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3572 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input9_A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4026 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1002 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input273_A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2288_A wire2288/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__465__A_N _593_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input440_A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__297__A _297_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3236 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1870 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_567_ _567_/A _567_/B vssd vssd vccd vccd _567_/X sky130_fd_sc_hd__and2_2
XFILLER_32_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2459 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_498_ _498_/A _498_/B vssd vssd vccd vccd _498_/X sky130_fd_sc_hd__and2_4
XANTENNA_output492_A wire1202/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1019_A wire1020/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__C _463_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2194 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output757_A wire1181/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1290_A _373_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput505 wire1272/X vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__buf_8
XANTENNA_wire1388_A wire1389/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput516 wire1261/X vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__buf_8
Xoutput527 wire1251/X vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__buf_8
XFILLER_9_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput538 wire1240/X vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__buf_8
XANTENNA_output924_A wire1393/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput549 wire1225/X vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__buf_8
XFILLER_42_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__000__A _000_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1322 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__488__A_N _616_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2246 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1803 wire1803/A vssd vssd vccd vccd wire1803/X sky130_fd_sc_hd__buf_6
Xwire1814 wire1815/X vssd vssd vccd vccd _366_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1825 wire1825/A vssd vssd vccd vccd _361_/A sky130_fd_sc_hd__buf_6
Xwire1836 wire1836/A vssd vssd vccd vccd _351_/A sky130_fd_sc_hd__buf_4
XFILLER_8_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1847 wire1848/X vssd vssd vccd vccd _291_/A sky130_fd_sc_hd__buf_6
XTAP_3103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1858 wire1858/A vssd vssd vccd vccd wire1858/X sky130_fd_sc_hd__buf_6
XTAP_3114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1869 wire1869/A vssd vssd vccd vccd wire1869/X sky130_fd_sc_hd__buf_6
XTAP_3125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2880 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2036_A wire2037/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_421_ _549_/A _421_/B _421_/C vssd vssd vccd vccd _421_/X sky130_fd_sc_hd__and3b_2
XANTENNA_136 _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _506_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 wire2263/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _352_/A _352_/B vssd vssd vccd vccd _352_/X sky130_fd_sc_hd__and2_4
XANTENNA__564__B _564_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2203_A wire2204/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_283_ _283_/A _283_/B vssd vssd vccd vccd _283_/X sky130_fd_sc_hd__and2_2
XFILLER_35_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input390_A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input84_A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__580__A _580_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput9 la_data_out_mprj[104] vssd vssd vccd vccd _473_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__458__C _458_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output505_A wire1272/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1136_A wire1136/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_619_ _619_/A _619_/B vssd vssd vccd vccd _619_/X sky130_fd_sc_hd__and2_4
XFILLER_35_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__B _474_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[117\]_B _280_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1303_A wire1304/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output874_A _309_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] _180_/X vssd vssd vccd vccd _000_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1672_A wire1672/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1937_A wire1937/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1094 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A mprj_dat_i_user[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__B _384_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_B _271_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput880 wire1452/X vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__buf_8
XFILLER_8_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2301 wire2301/A vssd vssd vccd vccd _295_/B sky130_fd_sc_hd__buf_6
Xoutput891 wire1021/X vssd vssd vccd vccd mprj_dat_i_core[19] sky130_fd_sc_hd__buf_8
XFILLER_25_3571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1600 wire1601/X vssd vssd vccd vccd wire1600/X sky130_fd_sc_hd__buf_6
XFILLER_24_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1611 wire1611/A vssd vssd vccd vccd wire1611/X sky130_fd_sc_hd__buf_6
XANTENNA__559__B _559_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input236_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2153_A wire2154/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1622 wire1623/X vssd vssd vccd vccd _329_/B sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[17\]_A mprj_dat_i_user[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1633 wire1634/X vssd vssd vccd vccd _326_/B sky130_fd_sc_hd__buf_6
Xwire1644 wire1644/A vssd vssd vccd vccd wire1644/X sky130_fd_sc_hd__buf_6
XFILLER_46_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1655 wire1656/X vssd vssd vccd vccd _321_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1666 wire1667/X vssd vssd vccd vccd _318_/B sky130_fd_sc_hd__buf_6
XFILLER_19_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1677 wire1678/X vssd vssd vccd vccd wire1677/X sky130_fd_sc_hd__buf_6
Xwire1688 wire1688/A vssd vssd vccd vccd _581_/A sky130_fd_sc_hd__buf_6
XFILLER_18_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1699 wire1699/A vssd vssd vccd vccd _570_/A sky130_fd_sc_hd__buf_8
XANTENNA_input403_A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__575__A _575_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_404_ _532_/A _404_/B _404_/C vssd vssd vccd vccd _404_/X sky130_fd_sc_hd__and3b_2
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__294__B _294_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_335_ _335_/A _335_/B vssd vssd vccd vccd _335_/X sky130_fd_sc_hd__and2_4
XFILLER_30_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_266_ _266_/A _266_/B vssd vssd vccd vccd _266_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire963 wire964/X vssd vssd vccd vccd wire963/X sky130_fd_sc_hd__buf_6
XFILLER_6_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire974 wire975/X vssd vssd vccd vccd wire974/X sky130_fd_sc_hd__buf_6
X_197_ _197_/A _197_/B vssd vssd vccd vccd _197_/X sky130_fd_sc_hd__and2_4
Xwire985 wire986/X vssd vssd vccd vccd wire985/X sky130_fd_sc_hd__buf_6
XFILLER_48_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire996 _139_/Y vssd vssd vccd vccd wire996/X sky130_fd_sc_hd__buf_6
XFILLER_26_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1086_A wire1087/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__469__B _469_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1253_A _409_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1420_A wire1421/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1518_A wire1518/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_14 _219_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_25 _230_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1887_A wire1887/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_36 _349_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_47 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_58 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_69 _291_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__379__B _379_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_120_ _120_/A vssd vssd vccd vccd _120_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_3114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_051_ _051_/A vssd vssd vccd vccd _051_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_49_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input186_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input353_A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1218 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input47_A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2120 wire2120/A vssd vssd vccd vccd wire2120/X sky130_fd_sc_hd__buf_6
XFILLER_27_2998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__289__B _289_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2131 wire2131/A vssd vssd vccd vccd _559_/B sky130_fd_sc_hd__buf_6
XFILLER_43_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2142 wire2142/A vssd vssd vccd vccd _516_/B sky130_fd_sc_hd__buf_6
Xwire2153 wire2154/X vssd vssd vccd vccd _506_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2164 wire2164/A vssd vssd vccd vccd wire2164/X sky130_fd_sc_hd__buf_6
XFILLER_43_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1430 wire1431/X vssd vssd vccd vccd wire1430/X sky130_fd_sc_hd__buf_8
Xwire2175 wire2175/A vssd vssd vccd vccd wire2175/X sky130_fd_sc_hd__buf_6
Xwire1441 wire1442/X vssd vssd vccd vccd wire1441/X sky130_fd_sc_hd__buf_8
XFILLER_1_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2186 wire2187/X vssd vssd vccd vccd wire2186/X sky130_fd_sc_hd__buf_6
Xwire2197 wire2198/X vssd vssd vccd vccd _486_/B sky130_fd_sc_hd__buf_6
Xwire1452 _298_/X vssd vssd vccd vccd wire1452/X sky130_fd_sc_hd__buf_6
XFILLER_46_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1463 _268_/X vssd vssd vccd vccd wire1463/X sky130_fd_sc_hd__buf_8
XFILLER_19_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1474 _248_/X vssd vssd vccd vccd wire1474/X sky130_fd_sc_hd__buf_8
Xwire1485 input96/X vssd vssd vccd vccd _437_/C sky130_fd_sc_hd__buf_6
XFILLER_1_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1496 wire1496/A vssd vssd vccd vccd wire1496/X sky130_fd_sc_hd__buf_6
XFILLER_46_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_318_ _318_/A _318_/B vssd vssd vccd vccd _318_/X sky130_fd_sc_hd__and2_4
XANTENNA_output572_A _452_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput12 la_data_out_mprj[107] vssd vssd vccd vccd _476_/C sky130_fd_sc_hd__clkbuf_4
Xinput23 la_data_out_mprj[117] vssd vssd vccd vccd input23/X sky130_fd_sc_hd__buf_6
Xinput34 la_data_out_mprj[127] vssd vssd vccd vccd _496_/C sky130_fd_sc_hd__clkbuf_4
Xinput45 la_data_out_mprj[21] vssd vssd vccd vccd _390_/C sky130_fd_sc_hd__clkbuf_4
X_249_ _249_/A _249_/B vssd vssd vccd vccd _249_/X sky130_fd_sc_hd__and2_4
XFILLER_45_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput56 la_data_out_mprj[31] vssd vssd vccd vccd _400_/C sky130_fd_sc_hd__clkbuf_4
Xinput67 la_data_out_mprj[41] vssd vssd vccd vccd _410_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput78 la_data_out_mprj[51] vssd vssd vccd vccd _420_/C sky130_fd_sc_hd__clkbuf_4
Xinput89 la_data_out_mprj[61] vssd vssd vccd vccd _430_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_28_2707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output837_A wire1145/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1370_A wire1371/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1468_A _254_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] wire1475/X vssd vssd vccd vccd wire1131/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2486 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1635_A wire1636/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1802_A wire1803/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire990_A wire991/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__381__C _381_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_4325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput405 mprj_adr_o_core[25] vssd vssd vccd vccd wire1621/A sky130_fd_sc_hd__buf_6
XFILLER_6_3760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput416 mprj_adr_o_core[6] vssd vssd vccd vccd wire1566/A sky130_fd_sc_hd__buf_6
XFILLER_2_3624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput427 mprj_dat_o_core[15] vssd vssd vccd vccd wire1535/A sky130_fd_sc_hd__buf_6
XFILLER_44_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput438 mprj_dat_o_core[25] vssd vssd vccd vccd wire1519/A sky130_fd_sc_hd__buf_6
XFILLER_9_1470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_2901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput449 mprj_dat_o_core[6] vssd vssd vccd vccd wire1504/A sky130_fd_sc_hd__buf_6
XFILLER_2_2923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_4002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input101_A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2116_A wire2116/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__572__B _572_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_103_ _103_/A vssd vssd vccd vccd _103_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4131 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_034_ _034_/A vssd vssd vccd vccd _034_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1260 _402_/X vssd vssd vccd vccd wire1260/X sky130_fd_sc_hd__buf_6
XFILLER_1_3178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_2372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1271 _392_/X vssd vssd vccd vccd wire1271/X sky130_fd_sc_hd__buf_6
Xwire1282 _381_/X vssd vssd vccd vccd wire1282/X sky130_fd_sc_hd__buf_6
XFILLER_19_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1293 _370_/X vssd vssd vccd vccd wire1293/X sky130_fd_sc_hd__buf_6
XFILLER_47_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1049_A wire1050/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__466__C _466_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output787_A _543_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3710 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__371__A_N _499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__B _482_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output954_A output954/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] split4/A vssd vssd vccd vccd _126_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_30_1918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1585_A wire1586/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__003__A _003_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] _273_/X vssd vssd vccd vccd _093_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_27_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__376__C _376_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_942 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__392__B _392_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_A mprj_dat_i_user[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1840 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput202 la_iena_mprj[48] vssd vssd vccd vccd _211_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput213 la_iena_mprj[58] vssd vssd vccd vccd _221_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput224 la_iena_mprj[68] vssd vssd vccd vccd _231_/B sky130_fd_sc_hd__buf_4
XTAP_4701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input149_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2066_A wire2067/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput235 la_iena_mprj[78] vssd vssd vccd vccd _241_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput246 la_iena_mprj[88] vssd vssd vccd vccd _251_/B sky130_fd_sc_hd__clkbuf_4
Xinput257 la_iena_mprj[98] vssd vssd vccd vccd _261_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput268 la_oenb_mprj[107] vssd vssd vccd vccd _604_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_40_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput279 la_oenb_mprj[117] vssd vssd vccd vccd wire1730/A sky130_fd_sc_hd__buf_6
XFILLER_29_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__567__B _567_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2233_A wire2233/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input316_A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_583_ _583_/A _583_/B vssd vssd vccd vccd _583_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__A_N _522_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__A _583_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput709 _074_/Y vssd vssd vccd vccd la_data_in_mprj[91] sky130_fd_sc_hd__buf_8
XFILLER_29_2813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_017_ _017_/A vssd vssd vccd vccd _017_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_46_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output535_A wire1290/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1166_A _539_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__477__B _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1333_A _359_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1090 _120_/Y vssd vssd vccd vccd wire1090/X sky130_fd_sc_hd__buf_6
XFILLER_47_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] _210_/X vssd vssd vccd vccd _030_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_14_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_706 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1967_A wire1967/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1748 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] _172_/X vssd vssd vccd vccd _156_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_28_1622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__387__B _387_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1014 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_293 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2183_A wire2184/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input266_A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input433_A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__578__A _578_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_566_ _566_/A _566_/B vssd vssd vccd vccd _566_/X sky130_fd_sc_hd__and2_2
XFILLER_38_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_497_ _497_/A _497_/B vssd vssd vccd vccd _497_/X sky130_fd_sc_hd__and2_4
XFILLER_32_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4572 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output485_A wire1283/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_3405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput506 wire1271/X vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__buf_8
Xoutput517 wire1260/X vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__buf_8
Xoutput528 wire1250/X vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__buf_8
XANTENNA_wire1283_A _380_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput539 wire1238/X vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__buf_8
XFILLER_10_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output917_A wire1358/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1450_A wire1451/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1548_A wire1548/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1715_A _409_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3370 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1804 wire1805/X vssd vssd vccd vccd _371_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1815 wire1815/A vssd vssd vccd vccd wire1815/X sky130_fd_sc_hd__buf_6
XFILLER_41_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1826 wire1826/A vssd vssd vccd vccd _360_/A sky130_fd_sc_hd__buf_6
XTAP_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1837 wire1837/A vssd vssd vccd vccd _350_/A sky130_fd_sc_hd__buf_4
Xwire1848 wire1849/X vssd vssd vccd vccd wire1848/X sky130_fd_sc_hd__buf_6
XTAP_3104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1859 wire1860/X vssd vssd vccd vccd _287_/A sky130_fd_sc_hd__buf_6
XTAP_3115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_104 _209_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_420_ _548_/A _420_/B _420_/C vssd vssd vccd vccd _420_/X sky130_fd_sc_hd__and3b_4
XANTENNA_137 _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _504_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _477_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2029_A wire2030/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_351_ _351_/A _351_/B vssd vssd vccd vccd _351_/X sky130_fd_sc_hd__and2_4
XFILLER_42_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_282_ _282_/A _282_/B vssd vssd vccd vccd _282_/X sky130_fd_sc_hd__and2_4
XANTENNA__432__A_N _560_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input383_A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__580__B _580_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input77_A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4036 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__101__A _101_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ _618_/A _618_/B vssd vssd vccd vccd _618_/X sky130_fd_sc_hd__and2_4
XTAP_3693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1031_A wire1032/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1129_A wire1129/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__474__C _474_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_549_ _549_/A _549_/B vssd vssd vccd vccd _549_/X sky130_fd_sc_hd__and2_2
XFILLER_32_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3808 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output867_A _332_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__B _490_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1665_A wire1665/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3904 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2484 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1832_A wire1832/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[26\]_B split5/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__455__A_N _583_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__C _384_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3815 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput870 _307_/X vssd vssd vccd vccd mprj_adr_o_user[2] sky130_fd_sc_hd__buf_8
XFILLER_5_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput881 wire1116/X vssd vssd vccd vccd mprj_dat_i_core[0] sky130_fd_sc_hd__buf_8
Xwire2302 wire2303/X vssd vssd vccd vccd wire2302/X sky130_fd_sc_hd__buf_6
XFILLER_8_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput892 wire1111/X vssd vssd vccd vccd mprj_dat_i_core[1] sky130_fd_sc_hd__buf_8
XFILLER_5_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1601 wire1601/A vssd vssd vccd vccd wire1601/X sky130_fd_sc_hd__buf_6
XFILLER_21_3447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1612 wire1613/X vssd vssd vccd vccd _331_/B sky130_fd_sc_hd__buf_8
Xwire1623 wire1624/X vssd vssd vccd vccd wire1623/X sky130_fd_sc_hd__buf_6
XFILLER_5_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1634 wire1635/X vssd vssd vccd vccd wire1634/X sky130_fd_sc_hd__buf_6
XFILLER_24_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[17\]_B load_slew1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1645 wire1646/X vssd vssd vccd vccd _324_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1656 wire1657/X vssd vssd vccd vccd wire1656/X sky130_fd_sc_hd__buf_6
XANTENNA_input131_A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1667 wire1667/A vssd vssd vccd vccd wire1667/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2146_A wire2146/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1678 wire1679/X vssd vssd vccd vccd wire1678/X sky130_fd_sc_hd__buf_6
XANTENNA_input229_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1689 wire1689/A vssd vssd vccd vccd _580_/A sky130_fd_sc_hd__buf_6
XFILLER_19_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__575__B _575_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _531_/A _403_/B _403_/C vssd vssd vccd vccd _403_/X sky130_fd_sc_hd__and3b_4
XTAP_2277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_334_ _334_/A _334_/B vssd vssd vccd vccd _334_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__591__A _591_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_265_ _265_/A _265_/B vssd vssd vccd vccd _265_/X sky130_fd_sc_hd__and2_4
XFILLER_13_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire964 wire965/X vssd vssd vccd vccd wire964/X sky130_fd_sc_hd__buf_6
X_196_ _196_/A _196_/B vssd vssd vccd vccd _196_/X sky130_fd_sc_hd__and2_4
Xwire975 wire976/X vssd vssd vccd vccd wire975/X sky130_fd_sc_hd__buf_6
XFILLER_10_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire986 _141_/Y vssd vssd vccd vccd wire986/X sky130_fd_sc_hd__buf_6
Xwire997 wire998/X vssd vssd vccd vccd wire997/X sky130_fd_sc_hd__buf_6
XFILLER_48_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1079_A wire1080/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__469__C _469_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1246_A _416_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__478__A_N _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__485__B _485_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1413_A _317_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_15 _220_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_26 _231_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_37 _312_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_48 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1782_A wire1783/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_59 _365_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__379__C _379_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_970 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__395__B _395_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2414 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_050_ _050_/A vssd vssd vccd vccd _050_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2096_A wire2096/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input179_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2263_A wire2264/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input346_A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2110 wire2110/A vssd vssd vccd vccd wire2110/X sky130_fd_sc_hd__buf_6
Xwire2121 wire2122/X vssd vssd vccd vccd _568_/B sky130_fd_sc_hd__buf_6
Xwire2132 wire2132/A vssd vssd vccd vccd _538_/B sky130_fd_sc_hd__buf_6
XFILLER_1_3305 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2143 wire2143/A vssd vssd vccd vccd _515_/B sky130_fd_sc_hd__buf_6
XFILLER_5_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2154 wire2154/A vssd vssd vccd vccd wire2154/X sky130_fd_sc_hd__buf_6
Xwire1420 wire1421/X vssd vssd vccd vccd wire1420/X sky130_fd_sc_hd__buf_6
Xwire2165 wire2166/X vssd vssd vccd vccd _498_/B sky130_fd_sc_hd__buf_6
Xwire1431 wire1432/X vssd vssd vccd vccd wire1431/X sky130_fd_sc_hd__buf_8
XFILLER_5_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2176 wire2177/X vssd vssd vccd vccd _493_/B sky130_fd_sc_hd__buf_6
Xwire1442 wire1443/X vssd vssd vccd vccd wire1442/X sky130_fd_sc_hd__buf_6
Xwire2187 wire2187/A vssd vssd vccd vccd wire2187/X sky130_fd_sc_hd__buf_6
Xwire1453 wire1454/X vssd vssd vccd vccd wire1453/X sky130_fd_sc_hd__buf_6
Xwire2198 wire2199/X vssd vssd vccd vccd wire2198/X sky130_fd_sc_hd__buf_6
XFILLER_4_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__586__A _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1464 _259_/X vssd vssd vccd vccd wire1464/X sky130_fd_sc_hd__buf_8
XFILLER_46_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1475 _247_/X vssd vssd vccd vccd wire1475/X sky130_fd_sc_hd__buf_8
Xwire1486 input95/X vssd vssd vccd vccd _436_/C sky130_fd_sc_hd__buf_6
XFILLER_21_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1497 wire1498/X vssd vssd vccd vccd _346_/B sky130_fd_sc_hd__buf_6
XFILLER_46_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_317_ _317_/A _317_/B vssd vssd vccd vccd _317_/X sky130_fd_sc_hd__and2_2
XFILLER_50_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput13 la_data_out_mprj[108] vssd vssd vccd vccd _477_/C sky130_fd_sc_hd__clkbuf_4
Xinput24 la_data_out_mprj[118] vssd vssd vccd vccd input24/X sky130_fd_sc_hd__buf_6
XFILLER_10_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_248_ _248_/A _248_/B vssd vssd vccd vccd _248_/X sky130_fd_sc_hd__and2_4
XFILLER_7_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput35 la_data_out_mprj[12] vssd vssd vccd vccd _381_/C sky130_fd_sc_hd__clkbuf_4
Xinput46 la_data_out_mprj[22] vssd vssd vccd vccd _391_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA_output565_A _446_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput57 la_data_out_mprj[32] vssd vssd vccd vccd _401_/C sky130_fd_sc_hd__clkbuf_4
Xinput68 la_data_out_mprj[42] vssd vssd vccd vccd _411_/C sky130_fd_sc_hd__clkbuf_4
Xinput79 la_data_out_mprj[52] vssd vssd vccd vccd _421_/C sky130_fd_sc_hd__buf_4
X_179_ _179_/A _179_/B vssd vssd vccd vccd _179_/X sky130_fd_sc_hd__and2_2
XANTENNA_wire1196_A _501_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output732_A _608_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1363_A _349_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] wire1482/X vssd vssd vccd vccd wire1138/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_38_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1530_A wire1531/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1628_A wire1629/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_726 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1997_A wire1997/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire983_A wire984/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_656 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1270 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput406 mprj_adr_o_core[26] vssd vssd vccd vccd wire1616/A sky130_fd_sc_hd__buf_6
XFILLER_9_2183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput417 mprj_adr_o_core[7] vssd vssd vccd vccd wire1563/A sky130_fd_sc_hd__buf_6
XFILLER_6_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput428 mprj_dat_o_core[16] vssd vssd vccd vccd wire1533/A sky130_fd_sc_hd__buf_6
XFILLER_2_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1230 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput439 mprj_dat_o_core[26] vssd vssd vccd vccd wire1518/A sky130_fd_sc_hd__buf_6
XFILLER_22_3564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2957 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2011_A wire2012/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2109_A wire2110/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input296_A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_102_ _102_/A vssd vssd vccd vccd _102_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_033_ _033_/A vssd vssd vccd vccd _033_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_4_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2857 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1250 _412_/X vssd vssd vccd vccd wire1250/X sky130_fd_sc_hd__buf_6
XFILLER_19_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1261 _401_/X vssd vssd vccd vccd wire1261/X sky130_fd_sc_hd__buf_6
XFILLER_47_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1272 _391_/X vssd vssd vccd vccd wire1272/X sky130_fd_sc_hd__buf_6
XFILLER_47_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1283 _380_/X vssd vssd vccd vccd wire1283/X sky130_fd_sc_hd__buf_6
Xwire1294 _369_/X vssd vssd vccd vccd wire1294/X sky130_fd_sc_hd__buf_6
XFILLER_38_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1111_A wire1112/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output682_A _050_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__C _482_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output947_A wire1430/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1480_A _242_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1578_A wire1579/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1745_A wire1745/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1912_A wire1912/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] _266_/X vssd vssd vccd vccd _086_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_25_203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__392__C _392_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[9\]_B max_cap1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1598 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput203 la_iena_mprj[49] vssd vssd vccd vccd _212_/B sky130_fd_sc_hd__buf_4
XFILLER_2_4145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[9\]_B _172_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput214 la_iena_mprj[59] vssd vssd vccd vccd _222_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput225 la_iena_mprj[69] vssd vssd vccd vccd _232_/B sky130_fd_sc_hd__buf_4
XFILLER_2_4167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 la_iena_mprj[79] vssd vssd vccd vccd _242_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 la_iena_mprj[89] vssd vssd vccd vccd _252_/B sky130_fd_sc_hd__clkbuf_4
Xinput258 la_iena_mprj[99] vssd vssd vccd vccd _262_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput269 la_oenb_mprj[108] vssd vssd vccd vccd _605_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_2_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2059_A wire2059/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input211_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_582_ _582_/A _582_/B vssd vssd vccd vccd _582_/X sky130_fd_sc_hd__and2_4
XFILLER_29_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2226_A wire2227/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input309_A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__B _583_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_958 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_016_ _016_/A vssd vssd vccd vccd _016_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__104__A _104_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output528_A wire1250/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1061_A wire1062/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1159_A _549_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__477__C _477_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1080 _122_/Y vssd vssd vccd vccd wire1080/X sky130_fd_sc_hd__buf_6
XFILLER_53_4523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1091 wire1092/X vssd vssd vccd vccd wire1091/X sky130_fd_sc_hd__buf_6
XANTENNA_output897_A wire997/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__493__B _493_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1862_A wire1863/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__387__C _387_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4011 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4006 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1774 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4135 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input161_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2176_A wire2177/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input259_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__578__B _578_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input426_A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input22_A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3274 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__594__A _594_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_565_ _565_/A _565_/B vssd vssd vccd vccd _565_/X sky130_fd_sc_hd__and2_2
XFILLER_18_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_496_ _624_/A _496_/B _496_/C vssd vssd vccd vccd _496_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3850 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output478_A _482_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput507 wire1270/X vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__buf_8
Xoutput518 wire1259/X vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__buf_8
XFILLER_29_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput529 wire1249/X vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__buf_8
XANTENNA_output645_A _016_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1276_A _387_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__488__B _488_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1443_A wire1444/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3898 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1610_A wire1611/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3750 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3663 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3794 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4072 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__384__A_N _512_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__398__B _398_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1805 wire1805/A vssd vssd vccd vccd wire1805/X sky130_fd_sc_hd__buf_6
XTAP_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1816 wire1817/X vssd vssd vccd vccd _365_/A sky130_fd_sc_hd__buf_6
Xwire1827 wire1827/A vssd vssd vccd vccd _359_/A sky130_fd_sc_hd__buf_6
XTAP_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1838 wire1839/X vssd vssd vccd vccd wire1838/X sky130_fd_sc_hd__buf_6
XFILLER_41_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1849 wire1849/A vssd vssd vccd vccd wire1849/X sky130_fd_sc_hd__buf_6
XTAP_3105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _168_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_127 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_138 _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_149 _504_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _350_/A _350_/B vssd vssd vccd vccd _350_/X sky130_fd_sc_hd__and2_4
XTAP_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_281_ _281_/A _281_/B vssd vssd vccd vccd _281_/X sky130_fd_sc_hd__and2_4
XFILLER_52_3195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input376_A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2293_A wire2293/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4048 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__589__A _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3264 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2552 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_617_ _617_/A _617_/B vssd vssd vccd vccd _617_/X sky130_fd_sc_hd__and2_4
XFILLER_45_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ _548_/A _548_/B vssd vssd vccd vccd _548_/X sky130_fd_sc_hd__and2_4
XTAP_2993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1024_A wire1025/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output595_A _086_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3956 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_479_ _607_/A _479_/B _479_/C vssd vssd vccd vccd _479_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4392 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output762_A wire1177/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__490__C _490_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1393_A wire1394/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1560_A wire1561/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1658_A wire1658/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__499__A _499_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3916 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2496 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1878 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1825_A wire1825/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3827 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput860 wire1400/X vssd vssd vccd vccd mprj_adr_o_user[20] sky130_fd_sc_hd__buf_8
XFILLER_5_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput871 _335_/X vssd vssd vccd vccd mprj_adr_o_user[30] sky130_fd_sc_hd__buf_8
XFILLER_9_3792 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput882 wire1066/X vssd vssd vccd vccd mprj_dat_i_core[10] sky130_fd_sc_hd__buf_8
XFILLER_21_4138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2900 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2303 wire2304/X vssd vssd vccd vccd wire2303/X sky130_fd_sc_hd__buf_6
XFILLER_47_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput893 wire1016/X vssd vssd vccd vccd mprj_dat_i_core[20] sky130_fd_sc_hd__buf_8
XANTENNA__202__A _202_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1602 wire1603/X vssd vssd vccd vccd _333_/B sky130_fd_sc_hd__buf_8
XFILLER_43_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1613 wire1614/X vssd vssd vccd vccd wire1613/X sky130_fd_sc_hd__buf_6
Xwire1624 wire1625/X vssd vssd vccd vccd wire1624/X sky130_fd_sc_hd__buf_6
Xwire1635 wire1636/X vssd vssd vccd vccd wire1635/X sky130_fd_sc_hd__buf_6
Xwire1646 wire1647/X vssd vssd vccd vccd wire1646/X sky130_fd_sc_hd__buf_6
XFILLER_24_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1657 wire1658/X vssd vssd vccd vccd wire1657/X sky130_fd_sc_hd__buf_6
XFILLER_3_3380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1668 wire1669/X vssd vssd vccd vccd _317_/B sky130_fd_sc_hd__buf_6
Xwire1679 wire1679/A vssd vssd vccd vccd wire1679/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2041_A wire2041/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input124_A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2139_A wire2139/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _530_/A _402_/B _402_/C vssd vssd vccd vccd _402_/X sky130_fd_sc_hd__and3b_2
XFILLER_15_3208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3388 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2306_A wire2306/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2676 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_333_ _333_/A _333_/B vssd vssd vccd vccd _333_/X sky130_fd_sc_hd__and2_4
XTAP_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2810 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__591__B _591_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_264_ _264_/A _264_/B vssd vssd vccd vccd _264_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_195_ _195_/A _195_/B vssd vssd vccd vccd _195_/X sky130_fd_sc_hd__and2_4
XFILLER_6_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire965 _146_/Y vssd vssd vccd vccd wire965/X sky130_fd_sc_hd__buf_6
XFILLER_48_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire976 wire977/X vssd vssd vccd vccd wire976/X sky130_fd_sc_hd__buf_6
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] split4/X vssd vssd vccd vccd _119_/A sky130_fd_sc_hd__nand2_4
Xwire987 wire988/X vssd vssd vccd vccd wire987/X sky130_fd_sc_hd__buf_6
Xwire998 wire999/X vssd vssd vccd vccd wire998/X sky130_fd_sc_hd__buf_6
XFILLER_48_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output510_A wire1266/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output608_A _098_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__485__C _485_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1406_A _321_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] _185_/X vssd vssd vccd vccd _005_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_32_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_16 _220_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_27 _233_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_38 _312_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_49 _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1775_A wire1775/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__022__A _022_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__422__A_N _550_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_982 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1274 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__395__C _395_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2089_A wire2089/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2100 wire2100/A vssd vssd vccd vccd wire2100/X sky130_fd_sc_hd__buf_6
Xoutput690 _057_/Y vssd vssd vccd vccd la_data_in_mprj[74] sky130_fd_sc_hd__buf_8
Xwire2111 wire2112/X vssd vssd vccd vccd _574_/B sky130_fd_sc_hd__buf_6
XFILLER_47_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input241_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2122 wire2122/A vssd vssd vccd vccd wire2122/X sky130_fd_sc_hd__buf_6
Xwire2133 wire2133/A vssd vssd vccd vccd _531_/B sky130_fd_sc_hd__buf_6
XANTENNA_input339_A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2144 wire2144/A vssd vssd vccd vccd _514_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire2256_A wire2257/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1410 wire1411/X vssd vssd vccd vccd wire1410/X sky130_fd_sc_hd__buf_6
Xwire2155 wire2155/A vssd vssd vccd vccd _505_/B sky130_fd_sc_hd__buf_6
XFILLER_5_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2166 wire2166/A vssd vssd vccd vccd wire2166/X sky130_fd_sc_hd__buf_6
Xwire1421 _314_/X vssd vssd vccd vccd wire1421/X sky130_fd_sc_hd__buf_6
XFILLER_25_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1432 wire1433/X vssd vssd vccd vccd wire1432/X sky130_fd_sc_hd__buf_6
Xwire2177 wire2178/X vssd vssd vccd vccd wire2177/X sky130_fd_sc_hd__buf_6
XFILLER_38_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2188 wire2189/X vssd vssd vccd vccd _489_/B sky130_fd_sc_hd__buf_6
Xwire1443 wire1444/X vssd vssd vccd vccd wire1443/X sky130_fd_sc_hd__buf_6
Xwire1454 wire1455/X vssd vssd vccd vccd wire1454/X sky130_fd_sc_hd__buf_6
Xwire2199 wire2199/A vssd vssd vccd vccd wire2199/X sky130_fd_sc_hd__buf_6
XFILLER_1_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1465 _258_/X vssd vssd vccd vccd wire1465/X sky130_fd_sc_hd__buf_6
XFILLER_4_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__586__B _586_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1476 _246_/X vssd vssd vccd vccd wire1476/X sky130_fd_sc_hd__buf_8
XFILLER_38_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_908 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1487 input94/X vssd vssd vccd vccd _435_/C sky130_fd_sc_hd__buf_6
Xwire1498 wire1498/A vssd vssd vccd vccd wire1498/X sky130_fd_sc_hd__buf_6
XFILLER_21_2599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3926 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_316_ _316_/A _316_/B vssd vssd vccd vccd _316_/X sky130_fd_sc_hd__and2_2
XFILLER_30_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__107__A _107_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput14 la_data_out_mprj[109] vssd vssd vccd vccd _478_/C sky130_fd_sc_hd__clkbuf_4
X_247_ _247_/A _247_/B vssd vssd vccd vccd _247_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput25 la_data_out_mprj[119] vssd vssd vccd vccd _488_/C sky130_fd_sc_hd__buf_4
Xinput36 la_data_out_mprj[13] vssd vssd vccd vccd _382_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput47 la_data_out_mprj[23] vssd vssd vccd vccd _392_/C sky130_fd_sc_hd__clkbuf_4
Xinput58 la_data_out_mprj[33] vssd vssd vccd vccd _402_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput69 la_data_out_mprj[43] vssd vssd vccd vccd _412_/C sky130_fd_sc_hd__clkbuf_4
X_178_ _178_/A _178_/B vssd vssd vccd vccd _178_/X sky130_fd_sc_hd__and2_4
XFILLER_7_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output558_A _439_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1091_A wire1092/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[41\]_B _204_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1189_A _508_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__445__A_N _573_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output725_A _602_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1356_A wire1357/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__496__B _496_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1523_A wire1523/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire976_A wire977/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__017__A _017_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_B _195_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput407 mprj_adr_o_core[27] vssd vssd vccd vccd wire1611/A sky130_fd_sc_hd__buf_6
Xinput418 mprj_adr_o_core[8] vssd vssd vccd vccd wire1559/A sky130_fd_sc_hd__buf_6
Xinput429 mprj_dat_o_core[17] vssd vssd vccd vccd wire1531/A sky130_fd_sc_hd__buf_6
XFILLER_22_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_B _262_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_996 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2004_A wire2005/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_101_ _101_/A vssd vssd vccd vccd _101_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input191_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input289_A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_032_ _032_/A vssd vssd vccd vccd _032_/Y sky130_fd_sc_hd__inv_2
XANTENNA__468__A_N _596_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3410 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input456_A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input52_A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__597__A _597_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1240 wire1241/X vssd vssd vccd vccd wire1240/X sky130_fd_sc_hd__buf_6
XFILLER_1_2402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1251 _411_/X vssd vssd vccd vccd wire1251/X sky130_fd_sc_hd__buf_6
Xwire1262 _400_/X vssd vssd vccd vccd wire1262/X sky130_fd_sc_hd__buf_6
XFILLER_40_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1273 _390_/X vssd vssd vccd vccd wire1273/X sky130_fd_sc_hd__buf_6
Xwire1284 _379_/X vssd vssd vccd vccd wire1284/X sky130_fd_sc_hd__buf_6
XFILLER_1_2446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1295 wire1296/X vssd vssd vccd vccd wire1295/X sky130_fd_sc_hd__buf_8
XFILLER_47_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_2396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1104_A wire1105/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output842_A _593_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1473_A _249_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B _177_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1640_A wire1641/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1738_A input23/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__300__A _300_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1905_A wire1906/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput204 la_iena_mprj[4] vssd vssd vccd vccd _167_/B sky130_fd_sc_hd__clkbuf_4
Xinput215 la_iena_mprj[5] vssd vssd vccd vccd _168_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput226 la_iena_mprj[6] vssd vssd vccd vccd _169_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 la_iena_mprj[7] vssd vssd vccd vccd _170_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput248 la_iena_mprj[8] vssd vssd vccd vccd _171_/B sky130_fd_sc_hd__clkbuf_4
Xinput259 la_iena_mprj[9] vssd vssd vccd vccd _172_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__210__A _210_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2744 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_581_ _581_/A _581_/B vssd vssd vccd vccd _581_/X sky130_fd_sc_hd__and2_4
XFILLER_44_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input204_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2121_A wire2122/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2219_A wire2219/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1600 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_015_ _015_/A vssd vssd vccd vccd _015_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2583 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__120__A _120_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2469 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1054_A wire1055/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1070 _124_/Y vssd vssd vccd vccd wire1070/X sky130_fd_sc_hd__buf_6
XFILLER_35_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1081 wire1082/X vssd vssd vccd vccd wire1081/X sky130_fd_sc_hd__buf_8
XFILLER_47_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1092 wire1093/X vssd vssd vccd vccd wire1092/X sky130_fd_sc_hd__buf_6
XFILLER_53_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1221_A _461_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output792_A wire1160/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1319_A wire1320/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__493__C _493_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1590_A wire1591/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3586 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1688_A wire1688/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1855_A wire1855/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__030__A _030_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1328 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_321 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_4089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1330 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__205__A _205_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input154_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2071_A wire2072/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2169_A wire2170/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2609 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input321_A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input419_A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__594__B _594_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_564_ _564_/A _564_/B vssd vssd vccd vccd _564_/X sky130_fd_sc_hd__and2_2
XTAP_3898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_495_ _623_/A _495_/B _495_/C vssd vssd vccd vccd _495_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_3406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3862 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1403 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput508 wire1269/X vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__buf_8
Xoutput519 wire1258/X vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__buf_8
XFILLER_49_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output540_A wire1236/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output638_A _010_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1171_A _531_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1269_A _394_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_ack_gate mprj_ack_i_user max_cap1456/X vssd vssd vccd vccd _146_/A sky130_fd_sc_hd__nand2_8
XFILLER_7_3197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__488__C _488_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output805_A _559_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2327 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1436_A wire1437/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] _215_/X vssd vssd vccd vccd _035_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_2040 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1603_A wire1604/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3762 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4084 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1972_A wire1973/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2660 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[29\]_A mprj_dat_i_user[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1806 wire1807/X vssd vssd vccd vccd _370_/B sky130_fd_sc_hd__buf_6
XFILLER_3_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input7_A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__398__C _398_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1817 wire1817/A vssd vssd vccd vccd wire1817/X sky130_fd_sc_hd__buf_6
XTAP_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1828 wire1828/A vssd vssd vccd vccd _358_/A sky130_fd_sc_hd__buf_6
XTAP_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1839 wire1840/X vssd vssd vccd vccd wire1839/X sky130_fd_sc_hd__buf_6
XFILLER_41_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_106 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_128 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_280_ _280_/A _280_/B vssd vssd vccd vccd _280_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3136 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input271_A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2286_A wire2286/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input369_A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__589__B _589_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ _616_/A _616_/B vssd vssd vccd vccd _616_/X sky130_fd_sc_hd__and2_4
XFILLER_17_343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_547_ _547_/A _547_/B vssd vssd vccd vccd _547_/X sky130_fd_sc_hd__and2_2
XFILLER_35_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_478_ _606_/A _478_/B _478_/C vssd vssd vccd vccd _478_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output490_A wire1204/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1017_A wire1018/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output588_A _467_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1812 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output755_A wire1183/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1386_A wire1387/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3248 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output922_A wire1343/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__499__B _499_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1553_A wire1554/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3928 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1720_A _400_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1818_A wire1819/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_4102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3456 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_4231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3839 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput850 wire1414/X vssd vssd vccd vccd mprj_adr_o_user[11] sky130_fd_sc_hd__buf_8
XFILLER_25_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput861 _326_/X vssd vssd vccd vccd mprj_adr_o_user[21] sky130_fd_sc_hd__buf_8
XFILLER_47_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput872 _336_/X vssd vssd vccd vccd mprj_adr_o_user[31] sky130_fd_sc_hd__buf_8
XFILLER_5_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput883 wire1061/X vssd vssd vccd vccd mprj_dat_i_core[11] sky130_fd_sc_hd__buf_8
Xwire2304 wire2305/X vssd vssd vccd vccd wire2304/X sky130_fd_sc_hd__buf_6
Xoutput894 wire1011/X vssd vssd vccd vccd mprj_dat_i_core[21] sky130_fd_sc_hd__buf_8
XFILLER_43_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3416 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1603 wire1604/X vssd vssd vccd vccd wire1603/X sky130_fd_sc_hd__buf_6
XFILLER_43_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1614 wire1615/X vssd vssd vccd vccd wire1614/X sky130_fd_sc_hd__buf_6
XFILLER_8_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1625 wire1626/X vssd vssd vccd vccd wire1625/X sky130_fd_sc_hd__buf_6
XFILLER_3_4093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1636 wire1636/A vssd vssd vccd vccd wire1636/X sky130_fd_sc_hd__buf_6
XTAP_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1647 wire1647/A vssd vssd vccd vccd wire1647/X sky130_fd_sc_hd__buf_6
XFILLER_41_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1658 wire1658/A vssd vssd vccd vccd wire1658/X sky130_fd_sc_hd__buf_6
Xwire1669 wire1670/X vssd vssd vccd vccd wire1669/X sky130_fd_sc_hd__buf_6
XFILLER_3_3392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2034_A wire2034/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_401_ _529_/A _401_/B _401_/C vssd vssd vccd vccd _401_/X sky130_fd_sc_hd__and3b_2
XFILLER_27_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_332_ _332_/A _332_/B vssd vssd vccd vccd _332_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire2201_A wire2202/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_263_ _263_/A _263_/B vssd vssd vccd vccd _263_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input82_A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_194_ _194_/A _194_/B vssd vssd vccd vccd _194_/X sky130_fd_sc_hd__and2_4
Xwire966 wire967/X vssd vssd vccd vccd wire966/X sky130_fd_sc_hd__buf_6
Xwire977 _143_/Y vssd vssd vccd vccd wire977/X sky130_fd_sc_hd__buf_6
XFILLER_6_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire988 wire989/X vssd vssd vccd vccd wire988/X sky130_fd_sc_hd__buf_6
Xwire999 wire999/A vssd vssd vccd vccd wire999/X sky130_fd_sc_hd__buf_6
XFILLER_6_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output503_A wire1274/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1134_A wire1134/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__374__A_N _502_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_4308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1301_A wire1302/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output872_A _336_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_17 _221_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] split5/X vssd vssd vccd vccd _142_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_28 _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] _178_/X vssd vssd vccd vccd _162_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_33_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_39 _312_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1670_A wire1670/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1768_A wire1769/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__303__A _303_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1935_A wire1935/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3736 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] _289_/X vssd vssd vccd vccd _109_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_4244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_994 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_110 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3647 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__213__A _213_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput680 _048_/Y vssd vssd vccd vccd la_data_in_mprj[65] sky130_fd_sc_hd__buf_8
Xwire2101 wire2102/X vssd vssd vccd vccd _579_/B sky130_fd_sc_hd__buf_6
Xoutput691 _058_/Y vssd vssd vccd vccd la_data_in_mprj[75] sky130_fd_sc_hd__buf_8
Xwire2112 wire2112/A vssd vssd vccd vccd wire2112/X sky130_fd_sc_hd__buf_6
XFILLER_43_1513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2123 wire2123/A vssd vssd vccd vccd _567_/B sky130_fd_sc_hd__buf_6
XFILLER_25_3382 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2134 wire2134/A vssd vssd vccd vccd _530_/B sky130_fd_sc_hd__buf_4
XFILLER_47_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1400 wire1401/X vssd vssd vccd vccd wire1400/X sky130_fd_sc_hd__buf_6
XFILLER_5_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire2145 wire2145/A vssd vssd vccd vccd _513_/B sky130_fd_sc_hd__buf_6
Xwire2156 wire2156/A vssd vssd vccd vccd _504_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1411 _318_/X vssd vssd vccd vccd wire1411/X sky130_fd_sc_hd__buf_6
XFILLER_1_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2151_A wire2151/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2167 wire2168/X vssd vssd vccd vccd _497_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1422 _313_/X vssd vssd vccd vccd wire1422/X sky130_fd_sc_hd__buf_6
XFILLER_25_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input234_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2178 wire2178/A vssd vssd vccd vccd wire2178/X sky130_fd_sc_hd__buf_6
Xwire1433 wire1434/X vssd vssd vccd vccd wire1433/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2249_A wire2249/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1444 _301_/X vssd vssd vccd vccd wire1444/X sky130_fd_sc_hd__buf_6
XFILLER_38_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2189 wire2190/X vssd vssd vccd vccd wire2189/X sky130_fd_sc_hd__buf_6
XFILLER_5_2786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1455 _296_/X vssd vssd vccd vccd wire1455/X sky130_fd_sc_hd__buf_6
Xwire1466 _256_/X vssd vssd vccd vccd wire1466/X sky130_fd_sc_hd__buf_6
XFILLER_1_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__397__A_N _525_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1477 _245_/X vssd vssd vccd vccd wire1477/X sky130_fd_sc_hd__buf_8
XFILLER_47_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1488 input93/X vssd vssd vccd vccd _434_/C sky130_fd_sc_hd__buf_6
XFILLER_41_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1499 wire1500/X vssd vssd vccd vccd _345_/B sky130_fd_sc_hd__buf_6
XTAP_2010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input401_A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_315_ _315_/A _315_/B vssd vssd vccd vccd _315_/X sky130_fd_sc_hd__and2_2
XTAP_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_246_ _246_/A _246_/B vssd vssd vccd vccd _246_/X sky130_fd_sc_hd__and2_4
XFILLER_7_821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput15 la_data_out_mprj[10] vssd vssd vccd vccd _379_/C sky130_fd_sc_hd__clkbuf_4
Xinput26 la_data_out_mprj[11] vssd vssd vccd vccd _380_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput37 la_data_out_mprj[14] vssd vssd vccd vccd _383_/C sky130_fd_sc_hd__clkbuf_4
Xinput48 la_data_out_mprj[24] vssd vssd vccd vccd _393_/C sky130_fd_sc_hd__clkbuf_4
Xinput59 la_data_out_mprj[34] vssd vssd vccd vccd _403_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_177_ _177_/A _177_/B vssd vssd vccd vccd _177_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1084_A wire1085/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2467 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output620_A _109_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1251_A _411_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1349_A wire1350/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1516_A wire1516/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_942 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3562 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1103 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1885_A wire1885/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire969_A _145_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__033__A _033_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput408 mprj_adr_o_core[28] vssd vssd vccd vccd wire1606/A sky130_fd_sc_hd__buf_6
XFILLER_44_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput419 mprj_adr_o_core[9] vssd vssd vccd vccd wire1555/A sky130_fd_sc_hd__buf_6
XFILLER_6_3785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4027 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__208__A _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_100_ _100_/A vssd vssd vccd vccd _100_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_51_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_031_ _031_/A vssd vssd vccd vccd _031_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input184_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2199_A wire2199/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_824 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input351_A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input449_A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input45_A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__597__B _597_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1230 _427_/X vssd vssd vccd vccd wire1230/X sky130_fd_sc_hd__buf_6
XFILLER_40_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1241 _421_/X vssd vssd vccd vccd wire1241/X sky130_fd_sc_hd__buf_6
Xwire1252 _410_/X vssd vssd vccd vccd wire1252/X sky130_fd_sc_hd__buf_6
XFILLER_38_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1263 _399_/X vssd vssd vccd vccd wire1263/X sky130_fd_sc_hd__buf_6
XFILLER_5_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1274 _389_/X vssd vssd vccd vccd wire1274/X sky130_fd_sc_hd__buf_6
XFILLER_5_1871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1285 _378_/X vssd vssd vccd vccd wire1285/X sky130_fd_sc_hd__buf_6
Xwire1296 wire1297/X vssd vssd vccd vccd wire1296/X sky130_fd_sc_hd__buf_6
XFILLER_1_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__118__A _118_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__A_N _540_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output570_A _450_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_229_ _229_/A _229_/B vssd vssd vccd vccd _229_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1299_A wire1300/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output835_A wire1192/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1466_A _256_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] wire1477/X vssd vssd vccd vccd wire1133/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1633_A wire1634/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__300__B _300_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1800_A wire1801/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_4216 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2803 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1979 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_411 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__028__A _028_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2916 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput205 la_iena_mprj[50] vssd vssd vccd vccd _213_/B sky130_fd_sc_hd__clkbuf_4
Xinput216 la_iena_mprj[60] vssd vssd vccd vccd _223_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput227 la_iena_mprj[70] vssd vssd vccd vccd _233_/B sky130_fd_sc_hd__buf_4
XTAP_4704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput238 la_iena_mprj[80] vssd vssd vccd vccd _243_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 la_iena_mprj[90] vssd vssd vccd vccd _253_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__210__B _210_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_580_ _580_/A _580_/B vssd vssd vccd vccd _580_/X sky130_fd_sc_hd__and2_4
XFILLER_44_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3003 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2114_A wire2114/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__435__A_N _563_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input399_A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_014_ _014_/A vssd vssd vccd vccd _014_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_2805 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1060 _126_/Y vssd vssd vccd vccd wire1060/X sky130_fd_sc_hd__buf_6
XFILLER_53_4503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1071 wire1072/X vssd vssd vccd vccd wire1071/X sky130_fd_sc_hd__buf_6
Xwire1082 wire1083/X vssd vssd vccd vccd wire1082/X sky130_fd_sc_hd__buf_6
Xwire1093 wire1094/X vssd vssd vccd vccd wire1093/X sky130_fd_sc_hd__buf_6
XFILLER_47_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1047_A wire1048/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output785_A wire1165/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output952_A output952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] max_cap1456/X vssd vssd vccd vccd _124_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_12_3598 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1583_A wire1584/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1750_A wire1750/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1848_A wire1849/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3708 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__458__A_N _586_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2064_A wire2065/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input147_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2520 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2231_A wire2231/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input314_A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3218 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_563_ _563_/A _563_/B vssd vssd vccd vccd _563_/X sky130_fd_sc_hd__and2_2
XTAP_3888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_494_ _622_/A _494_/B _494_/C vssd vssd vccd vccd _494_/X sky130_fd_sc_hd__and3b_2
XFILLER_38_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2110 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2706 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput509 wire1267/X vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__buf_8
XFILLER_5_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output533_A wire1245/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1164_A _542_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3823 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1331_A wire1332/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1429_A _304_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] _208_/X vssd vssd vccd vccd _028_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_4355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_344 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_804 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1798_A wire1799/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__306__A _306_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1965_A wire1966/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] _170_/X vssd vssd vccd vccd _154_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_28_1433 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[29\]_B split5/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1807 wire1807/A vssd vssd vccd vccd wire1807/X sky130_fd_sc_hd__buf_6
Xwire1818 wire1819/X vssd vssd vccd vccd _301_/A sky130_fd_sc_hd__buf_6
XTAP_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1829 wire1829/A vssd vssd vccd vccd _357_/A sky130_fd_sc_hd__buf_6
XTAP_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_107 _208_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_118 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_129 _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__216__A _216_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input264_A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2279_A wire2279/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input431_A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2626 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ _615_/A _615_/B vssd vssd vccd vccd _615_/X sky130_fd_sc_hd__and2_4
XTAP_3663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_546_ _546_/A _546_/B vssd vssd vccd vccd _546_/X sky130_fd_sc_hd__and2_2
XFILLER_45_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_477_ _605_/A _477_/B _477_/C vssd vssd vccd vccd _477_/X sky130_fd_sc_hd__and3b_1
XFILLER_50_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output483_A _487_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1824 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output650_A _021_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output748_A wire1144/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1281_A _382_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2515 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1379_A wire1380/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output915_A wire1364/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1546_A wire1547/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_3861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1713_A wire1713/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1457 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire999_A wire999/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_678 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1112 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__036__A _036_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput840 _591_/X vssd vssd vccd vccd la_oenb_core[94] sky130_fd_sc_hd__buf_8
XFILLER_5_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput851 wire1412/X vssd vssd vccd vccd mprj_adr_o_user[12] sky130_fd_sc_hd__buf_8
XFILLER_43_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput862 wire1398/X vssd vssd vccd vccd mprj_adr_o_user[22] sky130_fd_sc_hd__buf_8
XFILLER_25_4287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput873 _308_/X vssd vssd vccd vccd mprj_adr_o_user[3] sky130_fd_sc_hd__buf_8
XFILLER_25_3553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput884 wire1056/X vssd vssd vccd vccd mprj_dat_i_core[12] sky130_fd_sc_hd__buf_8
Xwire2305 wire2306/X vssd vssd vccd vccd wire2305/X sky130_fd_sc_hd__buf_6
XFILLER_25_3575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput895 wire1006/X vssd vssd vccd vccd mprj_dat_i_core[22] sky130_fd_sc_hd__buf_8
XFILLER_43_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1335 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3428 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1604 wire1605/X vssd vssd vccd vccd wire1604/X sky130_fd_sc_hd__buf_6
XFILLER_28_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1615 wire1616/X vssd vssd vccd vccd wire1615/X sky130_fd_sc_hd__buf_6
XFILLER_41_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1626 wire1626/A vssd vssd vccd vccd wire1626/X sky130_fd_sc_hd__buf_6
Xwire1637 wire1638/X vssd vssd vccd vccd _325_/B sky130_fd_sc_hd__buf_6
XFILLER_19_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1648 wire1649/X vssd vssd vccd vccd _323_/B sky130_fd_sc_hd__buf_6
XTAP_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1659 wire1660/X vssd vssd vccd vccd _320_/B sky130_fd_sc_hd__buf_6
XFILLER_41_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_400_ _400_/A_N _400_/B _400_/C vssd vssd vccd vccd _400_/X sky130_fd_sc_hd__and3b_2
XTAP_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2027_A wire2028/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ _331_/A _331_/B vssd vssd vccd vccd _331_/X sky130_fd_sc_hd__and2_4
XFILLER_32_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_262_ _262_/A _262_/B vssd vssd vccd vccd _262_/X sky130_fd_sc_hd__and2_4
XFILLER_23_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input381_A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_193_ _193_/A _193_/B vssd vssd vccd vccd _193_/X sky130_fd_sc_hd__and2_2
XFILLER_6_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire967 wire968/X vssd vssd vccd vccd wire967/X sky130_fd_sc_hd__buf_6
XFILLER_13_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire978 wire979/X vssd vssd vccd vccd wire978/X sky130_fd_sc_hd__buf_6
XANTENNA_input75_A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire989 wire990/X vssd vssd vccd vccd wire989/X sky130_fd_sc_hd__buf_6
XFILLER_6_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_529_ _529_/A _529_/B vssd vssd vccd vccd _529_/X sky130_fd_sc_hd__and2_4
XTAP_2792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_18 _221_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_29 _604_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output865_A _330_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1663_A wire1664/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__303__B _303_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1830_A wire1830/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] _282_/X vssd vssd vccd vccd _102_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_0_3544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3659 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4051 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__213__B _213_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput670 _039_/Y vssd vssd vccd vccd la_data_in_mprj[56] sky130_fd_sc_hd__buf_8
XFILLER_25_4095 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput681 _049_/Y vssd vssd vccd vccd la_data_in_mprj[66] sky130_fd_sc_hd__buf_8
Xwire2102 wire2102/A vssd vssd vccd vccd wire2102/X sky130_fd_sc_hd__buf_6
XFILLER_5_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput692 _059_/Y vssd vssd vccd vccd la_data_in_mprj[76] sky130_fd_sc_hd__buf_8
XFILLER_40_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2113 wire2114/X vssd vssd vccd vccd _573_/B sky130_fd_sc_hd__buf_6
Xwire2124 wire2125/X vssd vssd vccd vccd _566_/B sky130_fd_sc_hd__buf_6
XFILLER_25_3394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire2135 wire2135/A vssd vssd vccd vccd _525_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2146 wire2146/A vssd vssd vccd vccd _512_/B sky130_fd_sc_hd__buf_6
Xwire1401 _325_/X vssd vssd vccd vccd wire1401/X sky130_fd_sc_hd__buf_6
Xwire1412 wire1413/X vssd vssd vccd vccd wire1412/X sky130_fd_sc_hd__buf_6
Xwire2157 wire2157/A vssd vssd vccd vccd _503_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2168 wire2168/A vssd vssd vccd vccd wire2168/X sky130_fd_sc_hd__buf_6
Xwire1423 _312_/X vssd vssd vccd vccd wire1423/X sky130_fd_sc_hd__buf_6
XFILLER_43_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2179 wire2180/X vssd vssd vccd vccd _492_/B sky130_fd_sc_hd__buf_6
Xwire1434 _303_/X vssd vssd vccd vccd wire1434/X sky130_fd_sc_hd__buf_6
Xwire1445 wire1446/X vssd vssd vccd vccd wire1445/X sky130_fd_sc_hd__buf_8
XFILLER_4_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2144_A wire2144/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1467 _255_/X vssd vssd vccd vccd wire1467/X sky130_fd_sc_hd__buf_6
XANTENNA_input227_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1478 _244_/X vssd vssd vccd vccd wire1478/X sky130_fd_sc_hd__buf_8
Xwire1489 input92/X vssd vssd vccd vccd _433_/C sky130_fd_sc_hd__buf_6
XFILLER_34_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1928 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3906 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_314_ _314_/A _314_/B vssd vssd vccd vccd _314_/X sky130_fd_sc_hd__and2_4
XTAP_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_245_ _245_/A _245_/B vssd vssd vccd vccd _245_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput16 la_data_out_mprj[110] vssd vssd vccd vccd _479_/C sky130_fd_sc_hd__buf_4
Xinput27 la_data_out_mprj[120] vssd vssd vccd vccd _489_/C sky130_fd_sc_hd__buf_4
XFILLER_45_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput38 la_data_out_mprj[15] vssd vssd vccd vccd _384_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput49 la_data_out_mprj[25] vssd vssd vccd vccd _394_/C sky130_fd_sc_hd__clkbuf_4
X_176_ _176_/A _176_/B vssd vssd vccd vccd _176_/X sky130_fd_sc_hd__and2_2
XFILLER_7_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1077_A wire1078/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1244_A _418_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1990 wire1991/X vssd vssd vccd vccd _625_/A sky130_fd_sc_hd__buf_6
XFILLER_53_729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1411_A _318_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1509_A wire1510/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__491__A_N _619_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_290 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_114 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1780_A wire1781/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1878_A wire1878/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_6_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput409 mprj_adr_o_core[29] vssd vssd vccd vccd wire1601/A sky130_fd_sc_hd__buf_6
XFILLER_44_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3330 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1040 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__208__B _208_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_030_ _030_/A vssd vssd vccd vccd _030_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_3972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__224__A _224_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input177_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2094_A wire2094/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input344_A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2261_A wire2261/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input38_A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1220 _462_/X vssd vssd vccd vccd wire1220/X sky130_fd_sc_hd__buf_6
Xwire1231 _426_/X vssd vssd vccd vccd wire1231/X sky130_fd_sc_hd__buf_6
Xwire1242 _420_/X vssd vssd vccd vccd wire1242/X sky130_fd_sc_hd__buf_6
XFILLER_47_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1253 _409_/X vssd vssd vccd vccd wire1253/X sky130_fd_sc_hd__buf_6
XFILLER_19_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1264 _398_/X vssd vssd vccd vccd wire1264/X sky130_fd_sc_hd__buf_6
XFILLER_38_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1275 _388_/X vssd vssd vccd vccd wire1275/X sky130_fd_sc_hd__buf_6
Xwire1286 _377_/X vssd vssd vccd vccd wire1286/X sky130_fd_sc_hd__buf_6
XFILLER_1_2459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1297 wire1298/X vssd vssd vccd vccd wire1297/X sky130_fd_sc_hd__buf_6
XFILLER_35_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_228_ _228_/A _228_/B vssd vssd vccd vccd _228_/X sky130_fd_sc_hd__and2_2
XFILLER_7_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output563_A _444_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3209 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_159_ _159_/A vssd vssd vccd vccd _159_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1194_A _503_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output730_A wire1190/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3016 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output828_A _580_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1361_A wire1362/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] _238_/X vssd vssd vccd vccd _058_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1626_A wire1626/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__309__A _309_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1995_A wire1996/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire981_A _142_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__044__A _044_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__387__A_N _515_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3787 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput206 la_iena_mprj[51] vssd vssd vccd vccd _214_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput217 la_iena_mprj[61] vssd vssd vccd vccd _224_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput228 la_iena_mprj[71] vssd vssd vccd vccd _234_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_6_3594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput239 la_iena_mprj[81] vssd vssd vccd vccd _244_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2882 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2107_A wire2108/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input294_A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_013_ _013_/A vssd vssd vccd vccd _013_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input461_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3106 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1050 _128_/Y vssd vssd vccd vccd wire1050/X sky130_fd_sc_hd__buf_6
XFILLER_48_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1061 wire1062/X vssd vssd vccd vccd wire1061/X sky130_fd_sc_hd__buf_6
XFILLER_2_3981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1072 wire1073/X vssd vssd vccd vccd wire1072/X sky130_fd_sc_hd__buf_6
XFILLER_38_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1083 wire1084/X vssd vssd vccd vccd wire1083/X sky130_fd_sc_hd__buf_6
XFILLER_1_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1094 wire1095/X vssd vssd vccd vccd wire1094/X sky130_fd_sc_hd__buf_6
XFILLER_53_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output778_A wire1170/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output945_A wire1440/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3017 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1576_A wire1576/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3927 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__311__B _311_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] _264_/X vssd vssd vccd vccd _084_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_17_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__039__A _039_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_2618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1933 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__502__A _502_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2057_A wire2057/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__402__A_N _530_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_562_ _562_/A _562_/B vssd vssd vccd vccd _562_/X sky130_fd_sc_hd__and2_2
XTAP_3878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2224_A wire2225/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input307_A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_493_ _621_/A _493_/B _493_/C vssd vssd vccd vccd _493_/X sky130_fd_sc_hd__and3b_2
XFILLER_44_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2718 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2371 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output526_A wire1252/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_2268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1324_A wire1325/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output895_A wire1006/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_356 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_816 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] _201_/X vssd vssd vccd vccd _021_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__306__B _306_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1860_A wire1860/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1958_A wire1958/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4210 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__425__A_N _553_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1808 wire1809/X vssd vssd vccd vccd _369_/B sky130_fd_sc_hd__buf_6
XFILLER_23_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1819 wire1819/A vssd vssd vccd vccd wire1819/X sky130_fd_sc_hd__buf_6
XTAP_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_108 _192_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_119 _166_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_551 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2415 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__216__B _216_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_B wire1479/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__232__A _232_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input257_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2174_A wire2175/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2638 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3041 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input424_A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2419 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_614_ _614_/A _614_/B vssd vssd vccd vccd _614_/X sky130_fd_sc_hd__and2_4
XTAP_4398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_545_ _545_/A _545_/B vssd vssd vccd vccd _545_/X sky130_fd_sc_hd__and2_4
XFILLER_35_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_476_ _604_/A _476_/B _476_/C vssd vssd vccd vccd _476_/X sky130_fd_sc_hd__and3b_2
XFILLER_38_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output476_A _480_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[71\]_B _234_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__448__A_N _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output643_A _014_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__142__A _142_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1274_A _389_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output908_A wire1091/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1441_A wire1442/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput830 _582_/X vssd vssd vccd vccd la_oenb_core[85] sky130_fd_sc_hd__buf_8
XANTENNA__052__A _052_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput841 _592_/X vssd vssd vccd vccd la_oenb_core[95] sky130_fd_sc_hd__buf_8
XFILLER_8_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput852 wire1410/X vssd vssd vccd vccd mprj_adr_o_user[13] sky130_fd_sc_hd__buf_8
XFILLER_47_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput863 wire1397/X vssd vssd vccd vccd mprj_adr_o_user[23] sky130_fd_sc_hd__buf_8
XFILLER_8_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput874 _309_/X vssd vssd vccd vccd mprj_adr_o_user[4] sky130_fd_sc_hd__buf_8
XFILLER_25_4299 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput885 wire1051/X vssd vssd vccd vccd mprj_dat_i_core[13] sky130_fd_sc_hd__buf_8
Xwire2306 wire2306/A vssd vssd vccd vccd wire2306/X sky130_fd_sc_hd__buf_6
Xoutput896 wire1002/X vssd vssd vccd vccd mprj_dat_i_core[23] sky130_fd_sc_hd__buf_8
XFILLER_25_2831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1605 wire1606/X vssd vssd vccd vccd wire1605/X sky130_fd_sc_hd__buf_6
Xwire1616 wire1616/A vssd vssd vccd vccd wire1616/X sky130_fd_sc_hd__buf_6
XTAP_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1627 wire1628/X vssd vssd vccd vccd _328_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_2897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1638 wire1639/X vssd vssd vccd vccd wire1638/X sky130_fd_sc_hd__buf_6
Xwire1649 wire1650/X vssd vssd vccd vccd wire1649/X sky130_fd_sc_hd__buf_6
XFILLER_19_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_330_ _330_/A _330_/B vssd vssd vccd vccd _330_/X sky130_fd_sc_hd__and2_4
XFILLER_26_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__227__A _227_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_261_ _261_/A _261_/B vssd vssd vccd vccd _261_/X sky130_fd_sc_hd__and2_4
XFILLER_17_2370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_192_ _192_/A _192_/B vssd vssd vccd vccd _192_/X sky130_fd_sc_hd__and2_2
XFILLER_48_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire968 wire969/X vssd vssd vccd vccd wire968/X sky130_fd_sc_hd__buf_6
XFILLER_10_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire979 wire980/X vssd vssd vccd vccd wire979/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2291_A wire2291/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input374_A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input68_A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_528_ _528_/A _528_/B vssd vssd vccd vccd _528_/X sky130_fd_sc_hd__and2_4
XFILLER_50_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1022_A wire1023/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output593_A _084_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__137__A _137_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_19 _222_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_459_ _587_/A _459_/B _459_/C vssd vssd vccd vccd _459_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output760_A wire1179/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output858_A wire1402/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1391_A wire1392/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1656_A wire1657/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__600__A _600_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4257 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__047__A _047_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_2510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4317 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[35\]_B _198_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4063 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput660 _030_/Y vssd vssd vccd vccd la_data_in_mprj[47] sky130_fd_sc_hd__buf_8
XFILLER_5_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput671 _040_/Y vssd vssd vccd vccd la_data_in_mprj[57] sky130_fd_sc_hd__buf_8
Xoutput682 _050_/Y vssd vssd vccd vccd la_data_in_mprj[67] sky130_fd_sc_hd__buf_8
Xwire2103 wire2104/X vssd vssd vccd vccd _578_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2700 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput693 _060_/Y vssd vssd vccd vccd la_data_in_mprj[77] sky130_fd_sc_hd__buf_8
Xwire2114 wire2114/A vssd vssd vccd vccd wire2114/X sky130_fd_sc_hd__buf_6
XFILLER_5_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2125 wire2125/A vssd vssd vccd vccd wire2125/X sky130_fd_sc_hd__buf_6
XFILLER_40_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2136 wire2136/A vssd vssd vccd vccd _522_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2147 wire2148/X vssd vssd vccd vccd _511_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1402 _324_/X vssd vssd vccd vccd wire1402/X sky130_fd_sc_hd__buf_6
Xwire2158 wire2159/X vssd vssd vccd vccd _502_/B sky130_fd_sc_hd__buf_6
Xwire1413 _317_/X vssd vssd vccd vccd wire1413/X sky130_fd_sc_hd__buf_6
Xwire1424 wire1425/X vssd vssd vccd vccd wire1424/X sky130_fd_sc_hd__buf_6
Xwire2169 wire2170/X vssd vssd vccd vccd _496_/B sky130_fd_sc_hd__buf_6
Xwire1435 wire1436/X vssd vssd vccd vccd wire1435/X sky130_fd_sc_hd__buf_8
XFILLER_47_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1446 wire1447/X vssd vssd vccd vccd wire1446/X sky130_fd_sc_hd__buf_6
XFILLER_8_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1468 _254_/X vssd vssd vccd vccd wire1468/X sky130_fd_sc_hd__buf_6
Xwire1479 _243_/X vssd vssd vccd vccd wire1479/X sky130_fd_sc_hd__buf_6
XFILLER_38_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_3100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input122_A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2137_A wire2137/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2304_A wire2305/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_313_ _313_/A _313_/B vssd vssd vccd vccd _313_/X sky130_fd_sc_hd__and2_4
XTAP_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_244_ _244_/A _244_/B vssd vssd vccd vccd _244_/X sky130_fd_sc_hd__and2_4
XFILLER_10_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput17 la_data_out_mprj[111] vssd vssd vccd vccd _480_/C sky130_fd_sc_hd__buf_4
XFILLER_10_3642 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput28 la_data_out_mprj[121] vssd vssd vccd vccd _490_/C sky130_fd_sc_hd__buf_4
Xinput39 la_data_out_mprj[16] vssd vssd vccd vccd _385_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_175_ _175_/A _175_/B vssd vssd vccd vccd _175_/X sky130_fd_sc_hd__and2_4
XFILLER_6_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] max_cap1456/X vssd vssd vccd vccd _117_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_7_878 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1363 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[110\]_B _273_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_3126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1980 wire1981/X vssd vssd vccd vccd _168_/A sky130_fd_sc_hd__buf_6
XFILLER_19_963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1991 wire1991/A vssd vssd vccd vccd wire1991/X sky130_fd_sc_hd__buf_6
XFILLER_4_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_985 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1404_A wire1405/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_280 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] _183_/X vssd vssd vccd vccd _003_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_291 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__314__B _314_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_B _264_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1940_A wire1940/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2176 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__330__A _330_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_A mprj_dat_i_user[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__505__A _505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__224__B _224_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2087_A wire2087/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__240__A _240_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput490 wire1204/X vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__buf_8
XFILLER_43_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2254_A wire2254/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input337_A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1210 _474_/X vssd vssd vccd vccd wire1210/X sky130_fd_sc_hd__buf_6
XFILLER_21_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1221 _461_/X vssd vssd vccd vccd wire1221/X sky130_fd_sc_hd__buf_6
Xwire1232 wire1233/X vssd vssd vccd vccd wire1232/X sky130_fd_sc_hd__buf_6
XFILLER_21_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1243 _419_/X vssd vssd vccd vccd wire1243/X sky130_fd_sc_hd__buf_6
XFILLER_5_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1254 _408_/X vssd vssd vccd vccd wire1254/X sky130_fd_sc_hd__buf_6
XFILLER_21_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1265 _397_/X vssd vssd vccd vccd wire1265/X sky130_fd_sc_hd__buf_6
Xwire1276 _387_/X vssd vssd vccd vccd wire1276/X sky130_fd_sc_hd__buf_6
XFILLER_38_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1287 _376_/X vssd vssd vccd vccd wire1287/X sky130_fd_sc_hd__buf_6
Xwire1298 _368_/X vssd vssd vccd vccd wire1298/X sky130_fd_sc_hd__buf_6
XFILLER_5_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_4140 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_227_ _227_/A _227_/B vssd vssd vccd vccd _227_/X sky130_fd_sc_hd__and2_2
XFILLER_10_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_158_ _158_/A vssd vssd vccd vccd _158_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output556_A _438_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_089_ _089_/A vssd vssd vccd vccd _089_/Y sky130_fd_sc_hd__inv_2
XANTENNA_wire1187_A _510_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output723_A _600_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3844 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1354_A _352_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] _231_/X vssd vssd vccd vccd _051_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_22_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1521_A wire1521/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1619_A wire1620/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__309__B _309_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1890_A wire1890/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1988_A wire1989/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire974_A wire975/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1812 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3619 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__060__A _060_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput207 la_iena_mprj[52] vssd vssd vccd vccd _215_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput218 la_iena_mprj[62] vssd vssd vccd vccd _225_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput229 la_iena_mprj[72] vssd vssd vccd vccd _235_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_402 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2002_A wire2003/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__235__A _235_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input287_A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_012_ _012_/A vssd vssd vccd vccd _012_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_11_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input454_A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input50_A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__481__A_N _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3118 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__401__C _401_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1040 _130_/Y vssd vssd vccd vccd wire1040/X sky130_fd_sc_hd__buf_6
Xwire1051 wire1052/X vssd vssd vccd vccd wire1051/X sky130_fd_sc_hd__buf_6
Xwire1062 wire1063/X vssd vssd vccd vccd wire1062/X sky130_fd_sc_hd__buf_6
Xwire1073 wire1074/X vssd vssd vccd vccd wire1073/X sky130_fd_sc_hd__buf_6
XFILLER_2_3993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1084 wire1085/X vssd vssd vccd vccd wire1084/X sky130_fd_sc_hd__buf_6
XFILLER_35_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3902 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1095 _119_/Y vssd vssd vccd vccd wire1095/X sky130_fd_sc_hd__buf_6
XFILLER_53_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3859 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1102_A wire1103/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__145__A _145_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output840_A _591_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output938_A wire1388/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1471_A _251_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1569_A wire1570/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1384 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1903_A wire1904/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_265 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__055__A _055_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_max_cap1456_A split4/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__502__B _502_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1159 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_561_ _561_/A _561_/B vssd vssd vccd vccd _561_/X sky130_fd_sc_hd__and2_4
XTAP_3868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1854 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input202_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_492_ _620_/A _492_/B _492_/C vssd vssd vccd vccd _492_/X sky130_fd_sc_hd__and3b_2
XANTENNA_wire2217_A wire2217/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1411 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input98_A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__B _412_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2383 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_3908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output519_A wire1258/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1052_A wire1053/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__377__A_N _505_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output790_A wire1162/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_828 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1317_A wire1318/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output888_A wire1036/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_891 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1686_A wire1686/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__603__A _603_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1853_A wire1854/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__322__B _322_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3819 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[2\]_A mprj_dat_i_user[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1809 wire1809/A vssd vssd vccd vccd wire1809/X sky130_fd_sc_hd__buf_6
XTAP_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1056 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_109 _192_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_880 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_4133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__513__A _513_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__232__B _232_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input152_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2167_A wire2168/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input417_A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_613_ _613_/A _613_/B vssd vssd vccd vccd _613_/X sky130_fd_sc_hd__and2_4
XTAP_4388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_544_ _544_/A _544_/B vssd vssd vccd vccd _544_/X sky130_fd_sc_hd__and2_4
XTAP_3698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_475_ _603_/A _475_/B _475_/C vssd vssd vccd vccd _475_/X sky130_fd_sc_hd__and3b_1
XFILLER_31_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_585 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1350 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output469_A wire1210/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1267_A wire1268/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output803_A wire1149/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput390 mprj_adr_o_core[11] vssd vssd vccd vccd wire1672/A sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] _213_/X vssd vssd vccd vccd _033_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_35_143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1601_A wire1601/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_3448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__317__B _317_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1970_A wire1971/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__A _333_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput820 _573_/X vssd vssd vccd vccd la_oenb_core[76] sky130_fd_sc_hd__buf_8
XFILLER_47_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput831 _583_/X vssd vssd vccd vccd la_oenb_core[86] sky130_fd_sc_hd__buf_8
XFILLER_9_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput842 _593_/X vssd vssd vccd vccd la_oenb_core[96] sky130_fd_sc_hd__buf_8
Xoutput853 wire1408/X vssd vssd vccd vccd mprj_adr_o_user[14] sky130_fd_sc_hd__buf_8
XFILLER_9_3774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput864 _329_/X vssd vssd vccd vccd mprj_adr_o_user[24] sky130_fd_sc_hd__buf_8
XFILLER_43_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput875 _310_/X vssd vssd vccd vccd mprj_adr_o_user[5] sky130_fd_sc_hd__buf_8
XFILLER_5_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput886 wire1046/X vssd vssd vccd vccd mprj_dat_i_core[14] sky130_fd_sc_hd__buf_8
XFILLER_3_4030 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput897 wire997/X vssd vssd vccd vccd mprj_dat_i_core[24] sky130_fd_sc_hd__buf_8
XFILLER_3_4063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input5_A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1606 wire1606/A vssd vssd vccd vccd wire1606/X sky130_fd_sc_hd__buf_6
XFILLER_24_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1617 wire1618/X vssd vssd vccd vccd _330_/B sky130_fd_sc_hd__buf_8
XFILLER_47_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1628 wire1629/X vssd vssd vccd vccd wire1628/X sky130_fd_sc_hd__buf_6
XTAP_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1639 wire1639/A vssd vssd vccd vccd wire1639/X sky130_fd_sc_hd__buf_6
XTAP_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__508__A _508_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__227__B _227_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_260_ _260_/A _260_/B vssd vssd vccd vccd _260_/X sky130_fd_sc_hd__and2_4
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_191_ _191_/A _191_/B vssd vssd vccd vccd _191_/X sky130_fd_sc_hd__and2_2
XFILLER_22_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire969 _145_/Y vssd vssd vccd vccd wire969/X sky130_fd_sc_hd__buf_6
XFILLER_26_4009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__243__A _243_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2284_A wire2284/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input367_A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_irq_gates\[2\] user_irq_core[2] _293_/X vssd vssd vccd vccd _113_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_765 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2320 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_527_ _527_/A _527_/B vssd vssd vccd vccd _527_/X sky130_fd_sc_hd__and2_2
XFILLER_15_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_458_ _586_/A _458_/B _458_/C vssd vssd vccd vccd _458_/X sky130_fd_sc_hd__and3b_4
XANTENNA_wire1015_A _135_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__415__A_N _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output586_A wire1217/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_389_ _517_/A _389_/B _389_/C vssd vssd vccd vccd _389_/X sky130_fd_sc_hd__and3b_4
XFILLER_31_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output753_A wire1185/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1384_A _342_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output920_A wire1349/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] _261_/X vssd vssd vccd vccd wire1122/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_29_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1551_A wire1552/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1649_A wire1650/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__600__B _600_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1816_A wire1817/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__063__A _063_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4075 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput650 _021_/Y vssd vssd vccd vccd la_data_in_mprj[38] sky130_fd_sc_hd__buf_8
XFILLER_25_3341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput661 _031_/Y vssd vssd vccd vccd la_data_in_mprj[48] sky130_fd_sc_hd__buf_8
XFILLER_27_2949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput672 _041_/Y vssd vssd vccd vccd la_data_in_mprj[58] sky130_fd_sc_hd__buf_8
XFILLER_5_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput683 _051_/Y vssd vssd vccd vccd la_data_in_mprj[68] sky130_fd_sc_hd__buf_8
XFILLER_44_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2104 wire2104/A vssd vssd vccd vccd wire2104/X sky130_fd_sc_hd__buf_6
Xoutput694 _061_/Y vssd vssd vccd vccd la_data_in_mprj[78] sky130_fd_sc_hd__buf_8
Xwire2115 wire2116/X vssd vssd vccd vccd _572_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__510__B _510_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2126 wire2126/A vssd vssd vccd vccd _565_/B sky130_fd_sc_hd__buf_6
XFILLER_5_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2137 wire2137/A vssd vssd vccd vccd _521_/B sky130_fd_sc_hd__buf_6
Xwire2148 wire2148/A vssd vssd vccd vccd wire2148/X sky130_fd_sc_hd__buf_6
Xwire1403 _323_/X vssd vssd vccd vccd wire1403/X sky130_fd_sc_hd__buf_6
XFILLER_5_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1414 wire1415/X vssd vssd vccd vccd wire1414/X sky130_fd_sc_hd__buf_6
XFILLER_5_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2159 wire2159/A vssd vssd vccd vccd wire2159/X sky130_fd_sc_hd__buf_6
Xwire1425 _311_/X vssd vssd vccd vccd wire1425/X sky130_fd_sc_hd__buf_6
XFILLER_25_2695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1436 wire1437/X vssd vssd vccd vccd wire1436/X sky130_fd_sc_hd__buf_8
Xwire1447 wire1448/X vssd vssd vccd vccd wire1447/X sky130_fd_sc_hd__buf_6
Xwire1469 _253_/X vssd vssd vccd vccd wire1469/X sky130_fd_sc_hd__buf_8
XFILLER_28_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2032_A wire2033/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input115_A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__438__A_N _566_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__238__A _238_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_124 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2455 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _312_/A _312_/B vssd vssd vccd vccd _312_/X sky130_fd_sc_hd__and2_2
XFILLER_51_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_243_ _243_/A _243_/B vssd vssd vccd vccd _243_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1910 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput18 la_data_out_mprj[112] vssd vssd vccd vccd input18/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_input80_A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput29 la_data_out_mprj[122] vssd vssd vccd vccd _491_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_10_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_174_ _174_/A _174_/B vssd vssd vccd vccd _174_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3654 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__404__C _404_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2288 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1970 wire1971/X vssd vssd vccd vccd _175_/A sky130_fd_sc_hd__buf_6
XANTENNA_output501_A wire1275/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1981 wire1981/A vssd vssd vccd vccd wire1981/X sky130_fd_sc_hd__buf_6
XFILLER_19_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1992 wire1993/X vssd vssd vccd vccd _624_/B sky130_fd_sc_hd__buf_6
XFILLER_19_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1132_A wire1132/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_270 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_281 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output870_A _307_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1718 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] _176_/X vssd vssd vccd vccd _160_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] split5/A vssd vssd vccd vccd _140_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_20_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1599_A wire1600/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1766_A wire1767/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__611__A _611_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__330__B _330_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] _287_/X vssd vssd vccd vccd _107_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_42_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2686 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__058__A _058_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[10\]_B max_cap1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_477 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_rebuffer3_A split5/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__505__B _505_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3447 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__521__A _521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput480 _484_/X vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__buf_8
Xoutput491 wire1203/X vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__buf_8
XFILLER_40_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1200 _497_/X vssd vssd vccd vccd wire1200/X sky130_fd_sc_hd__buf_6
Xwire1211 _473_/X vssd vssd vccd vccd wire1211/X sky130_fd_sc_hd__buf_6
XFILLER_43_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1222 _460_/X vssd vssd vccd vccd wire1222/X sky130_fd_sc_hd__buf_6
XANTENNA_input232_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1233 _425_/X vssd vssd vccd vccd wire1233/X sky130_fd_sc_hd__buf_6
XFILLER_5_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1244 _418_/X vssd vssd vccd vccd wire1244/X sky130_fd_sc_hd__buf_6
XFILLER_21_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1255 _407_/X vssd vssd vccd vccd wire1255/X sky130_fd_sc_hd__buf_6
XFILLER_21_2367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1266 _396_/X vssd vssd vccd vccd wire1266/X sky130_fd_sc_hd__buf_6
Xwire1277 _386_/X vssd vssd vccd vccd wire1277/X sky130_fd_sc_hd__buf_6
XFILLER_19_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1288 _375_/X vssd vssd vccd vccd wire1288/X sky130_fd_sc_hd__buf_6
Xwire1299 wire1300/X vssd vssd vccd vccd wire1299/X sky130_fd_sc_hd__buf_8
XFILLER_38_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4152 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_226_ _226_/A _226_/B vssd vssd vccd vccd _226_/X sky130_fd_sc_hd__and2_2
XANTENNA__415__B _415_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_4196 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_157_ _157_/A vssd vssd vccd vccd _157_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_088_ _088_/A vssd vssd vccd vccd _088_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output549_A wire1225/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3981 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1082_A wire1083/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output716_A _081_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1347_A wire1348/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1514_A wire1514/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4085 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__606__A _606_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1883_A wire1883/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__325__B _325_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire967_A wire968/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1802 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3806 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__341__A _341_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4023 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput208 la_iena_mprj[53] vssd vssd vccd vccd _216_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput219 la_iena_mprj[63] vssd vssd vccd vccd _226_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3126 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__516__A _516_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__235__B _235_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_011_ _011_/A vssd vssd vccd vccd _011_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input182_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2197_A wire2198/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__251__A _251_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input447_A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input43_A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1030 _132_/Y vssd vssd vccd vccd wire1030/X sky130_fd_sc_hd__buf_6
XFILLER_40_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1041 wire1042/X vssd vssd vccd vccd wire1041/X sky130_fd_sc_hd__buf_6
XFILLER_2_3961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1052 wire1053/X vssd vssd vccd vccd wire1052/X sky130_fd_sc_hd__buf_6
XFILLER_38_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1063 wire1064/X vssd vssd vccd vccd wire1063/X sky130_fd_sc_hd__buf_6
XFILLER_53_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1074 wire1075/X vssd vssd vccd vccd wire1074/X sky130_fd_sc_hd__buf_6
XFILLER_48_889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1085 _121_/Y vssd vssd vccd vccd wire1085/X sky130_fd_sc_hd__buf_6
Xwire1096 wire1097/X vssd vssd vccd vccd wire1096/X sky130_fd_sc_hd__buf_6
XFILLER_1_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_528 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output499_A wire1277/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_209_ _209_/A _209_/B vssd vssd vccd vccd _209_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1297_A wire1298/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output833_A _585_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3907 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__161__A _161_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] wire1479/X vssd vssd vccd vccd wire1135/A
+ sky130_fd_sc_hd__nand2_4
XTAP_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1631_A wire1632/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__336__A _336_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__071__A _071_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3636 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_560_ _560_/A _560_/B vssd vssd vccd vccd _560_/X sky130_fd_sc_hd__and2_4
XTAP_3858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_491_ _619_/A _491_/B _491_/C vssd vssd vccd vccd _491_/X sky130_fd_sc_hd__and3b_1
XFILLER_35_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2112_A wire2112/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3980 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__246__A _246_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input397_A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__C _412_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4470 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3848 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1045_A _129_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3722 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3635 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_4011 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4180 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1212_A _472_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output783_A wire1166/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__156__A _156_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3332 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output950_A wire1445/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1581_A wire1581/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__603__B _603_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2126 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1846_A wire1846/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3759 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[2\]_B max_cap1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2832 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2854 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__471__A_N _599_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__066__A _066_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__513__B _513_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3400 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3444 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3466 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2062_A wire2063/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input145_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_612_ _612_/A _612_/B vssd vssd vccd vccd _612_/X sky130_fd_sc_hd__and2_4
XTAP_4378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input312_A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_543_ _543_/A _543_/B vssd vssd vccd vccd _543_/X sky130_fd_sc_hd__and2_4
XTAP_2932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_474_ _602_/A _474_/B _474_/C vssd vssd vccd vccd _474_/X sky130_fd_sc_hd__and3b_2
XFILLER_18_2339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__407__C _407_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3696 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__423__B _423_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output531_A wire1247/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output629_A _002_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3612 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1162_A wire1163/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput380 la_oenb_mprj[93] vssd vssd vccd vccd _590_/A sky130_fd_sc_hd__buf_6
XFILLER_42_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput391 mprj_adr_o_core[12] vssd vssd vccd vccd wire1670/A sky130_fd_sc_hd__buf_6
XFILLER_18_4220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1427_A wire1428/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__494__A_N _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] _206_/X vssd vssd vccd vccd _026_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_24_829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4128 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_166 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1796_A wire1797/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3162 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__A _614_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1963_A wire1964/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__333__B _333_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3720 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput810 _564_/X vssd vssd vccd vccd la_oenb_core[67] sky130_fd_sc_hd__buf_8
Xoutput821 _574_/X vssd vssd vccd vccd la_oenb_core[77] sky130_fd_sc_hd__buf_8
Xoutput832 _584_/X vssd vssd vccd vccd la_oenb_core[87] sky130_fd_sc_hd__buf_8
XFILLER_47_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput843 _594_/X vssd vssd vccd vccd la_oenb_core[97] sky130_fd_sc_hd__buf_8
XFILLER_9_3764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xoutput854 wire1407/X vssd vssd vccd vccd mprj_adr_o_user[15] sky130_fd_sc_hd__buf_8
XFILLER_5_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput865 _330_/X vssd vssd vccd vccd mprj_adr_o_user[25] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] _168_/X vssd vssd vccd vccd _152_/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_3786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput876 wire1424/X vssd vssd vccd vccd mprj_adr_o_user[6] sky130_fd_sc_hd__buf_8
XFILLER_8_2039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_4020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput887 wire1041/X vssd vssd vccd vccd mprj_dat_i_core[15] sky130_fd_sc_hd__buf_8
XFILLER_28_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2991 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput898 wire992/X vssd vssd vccd vccd mprj_dat_i_core[25] sky130_fd_sc_hd__buf_8
XFILLER_25_2844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1607 wire1608/X vssd vssd vccd vccd _332_/B sky130_fd_sc_hd__buf_8
XTAP_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1618 wire1619/X vssd vssd vccd vccd wire1618/X sky130_fd_sc_hd__buf_6
Xwire1629 wire1629/A vssd vssd vccd vccd wire1629/X sky130_fd_sc_hd__buf_6
XTAP_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__508__B _508_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_190_ _190_/A _190_/B vssd vssd vccd vccd _190_/X sky130_fd_sc_hd__and2_2
XFILLER_10_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__524__A _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__243__B _243_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input262_A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2277_A wire2277/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__418__B _418_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_526_ _526_/A _526_/B vssd vssd vccd vccd _526_/X sky130_fd_sc_hd__and2_4
XFILLER_50_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_457_ _585_/A _457_/B _457_/C vssd vssd vccd vccd _457_/X sky130_fd_sc_hd__and3b_4
XFILLER_53_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_388_ _516_/A _388_/B _388_/C vssd vssd vccd vccd _388_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output481_A _485_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1008_A wire1009/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output579_A wire1286/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output746_A _621_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1377_A wire1378/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output913_A wire1395/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1544_A wire1545/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1809_A wire1809/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__609__A _609_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_4050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__328__B _328_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire997_A wire998/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2692 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__344__A _344_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_30_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput640 _012_/Y vssd vssd vccd vccd la_data_in_mprj[29] sky130_fd_sc_hd__buf_8
XFILLER_5_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput651 _022_/Y vssd vssd vccd vccd la_data_in_mprj[39] sky130_fd_sc_hd__buf_8
XFILLER_25_4087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput662 _032_/Y vssd vssd vccd vccd la_data_in_mprj[49] sky130_fd_sc_hd__buf_8
Xoutput673 _042_/Y vssd vssd vccd vccd la_data_in_mprj[59] sky130_fd_sc_hd__buf_8
Xoutput684 _052_/Y vssd vssd vccd vccd la_data_in_mprj[69] sky130_fd_sc_hd__buf_8
Xwire2105 wire2106/X vssd vssd vccd vccd _577_/B sky130_fd_sc_hd__buf_6
XFILLER_40_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput695 _062_/Y vssd vssd vccd vccd la_data_in_mprj[79] sky130_fd_sc_hd__buf_8
Xwire2116 wire2116/A vssd vssd vccd vccd wire2116/X sky130_fd_sc_hd__buf_6
XFILLER_43_1517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2127 wire2127/A vssd vssd vccd vccd _564_/B sky130_fd_sc_hd__buf_6
Xwire2138 wire2138/A vssd vssd vccd vccd _520_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1404 wire1405/X vssd vssd vccd vccd wire1404/X sky130_fd_sc_hd__buf_6
Xwire2149 wire2150/X vssd vssd vccd vccd _510_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1415 wire1416/X vssd vssd vccd vccd wire1415/X sky130_fd_sc_hd__buf_6
Xwire1426 wire1427/X vssd vssd vccd vccd wire1426/X sky130_fd_sc_hd__buf_8
XFILLER_8_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1437 wire1438/X vssd vssd vccd vccd wire1437/X sky130_fd_sc_hd__buf_6
XFILLER_3_3171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1448 _300_/X vssd vssd vccd vccd wire1448/X sky130_fd_sc_hd__buf_6
XFILLER_28_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__519__A _519_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__238__B _238_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2025_A wire2025/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input108_A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _311_/A _311_/B vssd vssd vccd vccd _311_/X sky130_fd_sc_hd__and2_4
XTAP_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_242_ _242_/A _242_/B vssd vssd vccd vccd _242_/X sky130_fd_sc_hd__and2_2
XFILLER_52_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__254__A _254_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput19 la_data_out_mprj[113] vssd vssd vccd vccd input19/X sky130_fd_sc_hd__buf_6
XFILLER_7_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_173_ _173_/A _173_/B vssd vssd vccd vccd _173_/X sky130_fd_sc_hd__and2_1
XFILLER_32_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1977 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input73_A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1960 wire1960/A vssd vssd vccd vccd wire1960/X sky130_fd_sc_hd__buf_6
Xwire1971 wire1971/A vssd vssd vccd vccd wire1971/X sky130_fd_sc_hd__buf_6
XFILLER_20_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1982 wire1983/X vssd vssd vccd vccd _167_/A sky130_fd_sc_hd__buf_6
XFILLER_4_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1993 wire1994/X vssd vssd vccd vccd wire1993/X sky130_fd_sc_hd__buf_6
XTAP_3260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_4392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output696_A _154_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_271 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_509_ _509_/A _509_/B vssd vssd vccd vccd _509_/X sky130_fd_sc_hd__and2_1
XANTENNA_282 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output863_A wire1397/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__164__A _164_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] load_slew1458/X vssd vssd vccd vccd _133_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1494_A wire1495/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1661_A wire1662/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1759_A wire1759/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__611__B _611_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2073 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] _280_/X vssd vssd vccd vccd _100_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_0_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__074__A _074_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__521__B _521_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput470 wire1209/X vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__buf_8
XFILLER_44_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2769 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput481 _485_/X vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__buf_8
Xoutput492 wire1202/X vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__buf_8
XFILLER_40_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__405__A_N _405_/A_N vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1201 _496_/X vssd vssd vccd vccd wire1201/X sky130_fd_sc_hd__buf_6
XFILLER_25_2471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1212 _472_/X vssd vssd vccd vccd wire1212/X sky130_fd_sc_hd__buf_6
Xwire1223 _459_/X vssd vssd vccd vccd wire1223/X sky130_fd_sc_hd__buf_6
XFILLER_43_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1234 wire1235/X vssd vssd vccd vccd wire1234/X sky130_fd_sc_hd__buf_6
Xwire1245 _417_/X vssd vssd vccd vccd wire1245/X sky130_fd_sc_hd__buf_6
XFILLER_5_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1256 _406_/X vssd vssd vccd vccd wire1256/X sky130_fd_sc_hd__buf_6
Xwire1267 wire1268/X vssd vssd vccd vccd wire1267/X sky130_fd_sc_hd__buf_6
XANTENNA_input225_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1278 _385_/X vssd vssd vccd vccd wire1278/X sky130_fd_sc_hd__buf_6
Xwire1289 _374_/X vssd vssd vccd vccd wire1289/X sky130_fd_sc_hd__buf_6
XFILLER_34_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__249__A _249_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_4164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_225_ _225_/A _225_/B vssd vssd vccd vccd _225_/X sky130_fd_sc_hd__and2_2
XFILLER_11_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__415__C _415_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_156_ _156_/A vssd vssd vccd vccd _156_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1195 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_087_ _087_/A vssd vssd vccd vccd _087_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_49_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__B _431_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1075_A _123_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output709_A _074_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1242_A _420_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1790 wire1791/X vssd vssd vccd vccd _376_/B sky130_fd_sc_hd__buf_6
XFILLER_0_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_732 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1507_A wire1508/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2829 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__606__B _606_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1876_A wire1876/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__622__A _622_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_3818 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__341__B _341_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__428__A_N _556_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4254 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4035 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput209 la_iena_mprj[54] vssd vssd vccd vccd _217_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1022 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2885 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__069__A _069_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__516__B _516_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_010_ _010_/A vssd vssd vccd vccd _010_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__532__A _532_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3223 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2092_A wire2093/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input175_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input342_A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input36_A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1020 _134_/Y vssd vssd vccd vccd wire1020/X sky130_fd_sc_hd__buf_6
XFILLER_0_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1031 wire1032/X vssd vssd vccd vccd wire1031/X sky130_fd_sc_hd__buf_6
XFILLER_22_3890 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1042 wire1043/X vssd vssd vccd vccd wire1042/X sky130_fd_sc_hd__buf_6
Xwire1053 wire1054/X vssd vssd vccd vccd wire1053/X sky130_fd_sc_hd__buf_6
Xwire1064 wire1065/X vssd vssd vccd vccd wire1064/X sky130_fd_sc_hd__buf_6
XFILLER_38_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1075 _123_/Y vssd vssd vccd vccd wire1075/X sky130_fd_sc_hd__buf_6
Xwire1086 wire1087/X vssd vssd vccd vccd wire1086/X sky130_fd_sc_hd__buf_6
Xwire1097 wire1098/X vssd vssd vccd vccd wire1097/X sky130_fd_sc_hd__buf_6
XFILLER_53_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_4204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1235 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_208_ _208_/A _208_/B vssd vssd vccd vccd _208_/X sky130_fd_sc_hd__and2_2
XFILLER_45_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output561_A _442_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output659_A _029_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_139_ _139_/A vssd vssd vccd vccd _139_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2570 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output826_A _578_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] _236_/X vssd vssd vccd vccd _056_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1624_A wire1625/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_337 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__617__A _617_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1993_A wire1994/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__336__B _336_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_B wire1467/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__352__A _352_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3648 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3164 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_490_ _618_/A _490_/B _490_/C vssd vssd vccd vccd _490_/X sky130_fd_sc_hd__and3b_4
XANTENNA__527__A _527_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2105_A wire2106/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1435 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input292_A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_B wire1476/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__262__A _262_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1290 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4482 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1778 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1038_A wire1039/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4001 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3669 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2935 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output776_A _533_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_B _237_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output943_A wire1373/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__172__A _172_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1574_A wire1575/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3727 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1839_A wire1840/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2844 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__347__A _347_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__082__A _082_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3412 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3478 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input138_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2055_A wire2055/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_611_ _611_/A _611_/B vssd vssd vccd vccd _611_/X sky130_fd_sc_hd__and2_4
XFILLER_22_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_542_ _542_/A _542_/B vssd vssd vccd vccd _542_/X sky130_fd_sc_hd__and2_4
XTAP_3678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2222_A wire2223/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input305_A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__257__A _257_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_473_ _601_/A _473_/B _473_/C vssd vssd vccd vccd _473_/X sky130_fd_sc_hd__and3b_2
XFILLER_44_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_3691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3653 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[56\]_B _219_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__423__C _423_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3771 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output524_A wire1291/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3646 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1155_A _552_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput370 la_oenb_mprj[84] vssd vssd vccd vccd wire1688/A sky130_fd_sc_hd__buf_6
Xinput381 la_oenb_mprj[94] vssd vssd vccd vccd _591_/A sky130_fd_sc_hd__buf_6
XFILLER_7_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput392 mprj_adr_o_core[13] vssd vssd vccd vccd wire1667/A sky130_fd_sc_hd__buf_6
XFILLER_23_1367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4232 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output893_A wire1016/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_4167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__167__A _167_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] _199_/X vssd vssd vccd vccd _019_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2798 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[47\]_B _210_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1789_A wire1789/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__614__B _614_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1956_A wire1957/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput800 wire1150/X vssd vssd vccd vccd la_oenb_core[58] sky130_fd_sc_hd__buf_8
Xoutput811 _565_/X vssd vssd vccd vccd la_oenb_core[68] sky130_fd_sc_hd__buf_8
XFILLER_9_3732 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput822 _575_/X vssd vssd vccd vccd la_oenb_core[78] sky130_fd_sc_hd__buf_8
Xoutput833 _585_/X vssd vssd vccd vccd la_oenb_core[88] sky130_fd_sc_hd__buf_8
Xoutput844 _595_/X vssd vssd vccd vccd la_oenb_core[98] sky130_fd_sc_hd__buf_8
Xoutput855 wire1406/X vssd vssd vccd vccd mprj_adr_o_user[16] sky130_fd_sc_hd__buf_8
XFILLER_47_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput866 _331_/X vssd vssd vccd vccd mprj_adr_o_user[26] sky130_fd_sc_hd__buf_8
XFILLER_25_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput877 wire1423/X vssd vssd vccd vccd mprj_adr_o_user[7] sky130_fd_sc_hd__buf_8
Xoutput888 wire1036/X vssd vssd vccd vccd mprj_dat_i_core[16] sky130_fd_sc_hd__buf_8
XFILLER_28_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput899 wire987/X vssd vssd vccd vccd mprj_dat_i_core[26] sky130_fd_sc_hd__buf_8
XFILLER_25_3579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1608 wire1609/X vssd vssd vccd vccd wire1608/X sky130_fd_sc_hd__buf_6
XFILLER_28_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1619 wire1620/X vssd vssd vccd vccd wire1619/X sky130_fd_sc_hd__buf_6
XTAP_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2652 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__077__A _077_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3984 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_3848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[122\]_B _285_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__524__B _524_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_712 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__540__A _540_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3181 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2172_A wire2173/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input255_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_3056 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input422_A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[31\]_A mprj_dat_i_user[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_525_ _525_/A _525_/B vssd vssd vccd vccd _525_/X sky130_fd_sc_hd__and2_4
XTAP_2752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__418__C _418_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_456_ _584_/A _456_/B _456_/C vssd vssd vccd vccd _456_/X sky130_fd_sc_hd__and3b_4
XFILLER_18_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_387_ _515_/A _387_/B _387_/C vssd vssd vccd vccd _387_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__434__B _434_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[113\]_B _276_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1171 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output474_A wire1284/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3811 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output739_A _615_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3855 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1272_A _391_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__461__A_N _589_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4291 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3899 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output906_A wire1101/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__609__B _609_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1704_A wire1704/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[22\]_A mprj_dat_i_user[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__625__A _625_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1861 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__344__B _344_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_B _267_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput630 _148_/Y vssd vssd vccd vccd la_data_in_mprj[1] sky130_fd_sc_hd__buf_8
XANTENNA__360__A _360_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput641 _149_/Y vssd vssd vccd vccd la_data_in_mprj[2] sky130_fd_sc_hd__buf_8
Xoutput652 _150_/Y vssd vssd vccd vccd la_data_in_mprj[3] sky130_fd_sc_hd__buf_8
XFILLER_47_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput663 _151_/Y vssd vssd vccd vccd la_data_in_mprj[4] sky130_fd_sc_hd__buf_8
XFILLER_9_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput674 _152_/Y vssd vssd vccd vccd la_data_in_mprj[5] sky130_fd_sc_hd__buf_8
XFILLER_25_3354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput685 _153_/Y vssd vssd vccd vccd la_data_in_mprj[6] sky130_fd_sc_hd__buf_8
Xwire2106 wire2106/A vssd vssd vccd vccd wire2106/X sky130_fd_sc_hd__buf_6
XFILLER_47_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput696 _154_/Y vssd vssd vccd vccd la_data_in_mprj[7] sky130_fd_sc_hd__buf_8
Xwire2117 wire2117/A vssd vssd vccd vccd _571_/B sky130_fd_sc_hd__buf_6
Xwire2128 wire2128/A vssd vssd vccd vccd _563_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2139 wire2139/A vssd vssd vccd vccd _519_/B sky130_fd_sc_hd__buf_6
Xwire1405 _322_/X vssd vssd vccd vccd wire1405/X sky130_fd_sc_hd__buf_6
Xwire1416 _316_/X vssd vssd vccd vccd wire1416/X sky130_fd_sc_hd__buf_6
XFILLER_21_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1427 wire1428/X vssd vssd vccd vccd wire1427/X sky130_fd_sc_hd__buf_8
Xwire1438 wire1439/X vssd vssd vccd vccd wire1438/X sky130_fd_sc_hd__buf_6
XFILLER_41_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1449 wire1450/X vssd vssd vccd vccd wire1449/X sky130_fd_sc_hd__buf_6
XFILLER_3_3183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__519__B _519_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3136 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[13\]_A mprj_dat_i_user[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _310_/A _310_/B vssd vssd vccd vccd _310_/X sky130_fd_sc_hd__and2_4
XFILLER_42_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_660 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2018_A wire2019/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__535__A _535_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_241_ _241_/A _241_/B vssd vssd vccd vccd _241_/X sky130_fd_sc_hd__and2_4
XFILLER_51_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3612 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_172_ _172_/A _172_/B vssd vssd vccd vccd _172_/X sky130_fd_sc_hd__and2_4
XFILLER_49_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input372_A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__484__A_N _612_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input66_A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__270__A _270_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1950 wire1950/A vssd vssd vccd vccd _188_/A sky130_fd_sc_hd__buf_6
Xwire1961 wire1961/A vssd vssd vccd vccd _181_/A sky130_fd_sc_hd__buf_6
Xwire1972 wire1973/X vssd vssd vccd vccd _174_/A sky130_fd_sc_hd__buf_6
XFILLER_18_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1983 wire1983/A vssd vssd vccd vccd wire1983/X sky130_fd_sc_hd__buf_6
Xwire1994 wire1994/A vssd vssd vccd vccd wire1994/X sky130_fd_sc_hd__buf_6
XTAP_3250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__429__B _429_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_250 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1812 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_261 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_508_ _508_/A _508_/B vssd vssd vccd vccd _508_/X sky130_fd_sc_hd__and2_2
XFILLER_19_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_272 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1020_A _134_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_283 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1118_A wire1119/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output689_A _056_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ _567_/A _439_/B _439_/C vssd vssd vccd vccd _439_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output856_A wire1404/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_174 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__180__A _180_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_4228 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1654_A wire1654/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2179 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__339__B _339_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_446 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__355__A _355_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2381 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_3976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__090__A _090_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput471 wire1208/X vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__buf_8
Xoutput482 _486_/X vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__buf_8
Xoutput493 wire1201/X vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__buf_8
XFILLER_40_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1202 _495_/X vssd vssd vccd vccd wire1202/X sky130_fd_sc_hd__buf_6
XFILLER_5_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1213 _471_/X vssd vssd vccd vccd wire1213/X sky130_fd_sc_hd__buf_6
XFILLER_47_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1224 _458_/X vssd vssd vccd vccd wire1224/X sky130_fd_sc_hd__buf_6
Xwire1235 _424_/X vssd vssd vccd vccd wire1235/X sky130_fd_sc_hd__buf_6
Xwire1246 _416_/X vssd vssd vccd vccd wire1246/X sky130_fd_sc_hd__buf_6
XFILLER_5_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1257 _405_/X vssd vssd vccd vccd wire1257/X sky130_fd_sc_hd__buf_6
XFILLER_38_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1268 _395_/X vssd vssd vccd vccd wire1268/X sky130_fd_sc_hd__buf_6
Xwire1279 _384_/X vssd vssd vccd vccd wire1279/X sky130_fd_sc_hd__buf_6
XFILLER_1_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input120_A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input218_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4544 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2302_A wire2303/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__265__A _265_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_630 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_224_ _224_/A _224_/B vssd vssd vccd vccd _224_/X sky130_fd_sc_hd__and2_1
XFILLER_7_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_155_ _155_/A vssd vssd vccd vccd _155_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_6_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] max_cap1456/X vssd vssd vccd vccd _115_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_13_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3497 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_086_ _086_/A vssd vssd vccd vccd _086_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_23_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__C _431_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3983 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_2190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1068_A wire1069/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1780 wire1781/X vssd vssd vccd vccd _381_/B sky130_fd_sc_hd__buf_6
Xwire1791 wire1792/X vssd vssd vccd vccd wire1791/X sky130_fd_sc_hd__buf_6
XFILLER_19_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1402_A _324_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__175__A _175_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] rebuffer6/X vssd vssd vccd vccd _145_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_37_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3375 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1771_A wire1771/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__622__B _622_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4047 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1034 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1762 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__085__A _085_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3235 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input168_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2252_A wire2253/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input335_A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1010 _136_/Y vssd vssd vccd vccd wire1010/X sky130_fd_sc_hd__buf_6
XFILLER_25_2280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1021 wire1022/X vssd vssd vccd vccd wire1021/X sky130_fd_sc_hd__buf_6
Xwire1032 wire1033/X vssd vssd vccd vccd wire1032/X sky130_fd_sc_hd__buf_6
Xwire1043 wire1044/X vssd vssd vccd vccd wire1043/X sky130_fd_sc_hd__buf_6
XFILLER_47_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input29_A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_869 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1054 wire1055/X vssd vssd vccd vccd wire1054/X sky130_fd_sc_hd__buf_6
XFILLER_21_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1065 _125_/Y vssd vssd vccd vccd wire1065/X sky130_fd_sc_hd__buf_6
Xwire1076 wire1077/X vssd vssd vccd vccd wire1076/X sky130_fd_sc_hd__buf_6
XFILLER_1_2238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1087 wire1088/X vssd vssd vccd vccd wire1087/X sky130_fd_sc_hd__buf_6
XFILLER_38_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1098 wire1099/X vssd vssd vccd vccd wire1098/X sky130_fd_sc_hd__buf_6
XFILLER_38_2641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4396 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4238 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__426__C _426_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1203 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_207_ _207_/A _207_/B vssd vssd vccd vccd _207_/X sky130_fd_sc_hd__and2_4
XFILLER_50_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_138_ _138_/A vssd vssd vccd vccd _138_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__442__B _442_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output554_A _436_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2582 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_069_ _069_/A vssd vssd vccd vccd _069_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output721_A _598_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output819_A _572_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1352_A wire1353/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] _229_/X vssd vssd vccd vccd _049_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1617_A wire1618/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__617__B _617_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1986_A wire1987/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_1926 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire972_A wire973/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__352__B _352_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[5\]_A mprj_dat_i_user[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3132 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3176 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2683 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2000_A wire2000/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3868 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__543__A _543_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1870 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input285_A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__262__B _262_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1111 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1155 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input452_A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4494 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_1262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3724 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__437__B _437_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__418__A_N _546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1000 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output769_A wire1198/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output936_A wire1299/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4429 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1567_A wire1568/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_3739 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4186 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1901_A wire1902/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_390 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__347__B _347_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_894 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1567 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_2544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__A _363_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1516 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3227 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_610_ _610_/A _610_/B vssd vssd vccd vccd _610_/X sky130_fd_sc_hd__and2_4
XTAP_4358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2048_A wire2049/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__A _538_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_541_ _541_/A _541_/B vssd vssd vccd vccd _541_/X sky130_fd_sc_hd__and2_2
XTAP_2912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input200_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_472_ _600_/A _472_/B _472_/C vssd vssd vccd vccd _472_/X sky130_fd_sc_hd__and3b_4
XANTENNA__257__B _257_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1022 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2215_A wire2216/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_4480 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input96_A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__273__A _273_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2200 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output517_A wire1260/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput360 la_oenb_mprj[75] vssd vssd vccd vccd wire1697/A sky130_fd_sc_hd__buf_6
XFILLER_42_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput371 la_oenb_mprj[85] vssd vssd vccd vccd wire1687/A sky130_fd_sc_hd__buf_6
XFILLER_7_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput382 la_oenb_mprj[95] vssd vssd vccd vccd _592_/A sky130_fd_sc_hd__buf_6
XANTENNA_wire1050_A _128_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput393 mprj_adr_o_core[14] vssd vssd vccd vccd wire1665/A sky130_fd_sc_hd__buf_6
XFILLER_23_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4244 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1315_A wire1316/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output886_A wire1046/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] _192_/X vssd vssd vccd vccd _012_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA__390__A_N _518_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__183__A _183_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_3175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1684_A wire1684/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput801 _556_/X vssd vssd vccd vccd la_oenb_core[59] sky130_fd_sc_hd__buf_8
Xoutput812 _566_/X vssd vssd vccd vccd la_oenb_core[69] sky130_fd_sc_hd__buf_8
XANTENNA_wire1851_A wire1852/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput823 _576_/X vssd vssd vccd vccd la_oenb_core[79] sky130_fd_sc_hd__buf_8
XFILLER_9_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3503 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1949_A wire1949/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput834 wire1147/X vssd vssd vccd vccd la_oenb_core[89] sky130_fd_sc_hd__buf_8
Xoutput845 _596_/X vssd vssd vccd vccd la_oenb_core[99] sky130_fd_sc_hd__buf_8
Xoutput856 wire1404/X vssd vssd vccd vccd mprj_adr_o_user[17] sky130_fd_sc_hd__buf_8
XFILLER_3_4000 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput867 _332_/X vssd vssd vccd vccd mprj_adr_o_user[27] sky130_fd_sc_hd__buf_8
XFILLER_25_3547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput878 wire1422/X vssd vssd vccd vccd mprj_adr_o_user[8] sky130_fd_sc_hd__buf_8
XFILLER_47_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput889 wire1031/X vssd vssd vccd vccd mprj_dat_i_core[17] sky130_fd_sc_hd__buf_8
XFILLER_3_4033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1609 wire1610/X vssd vssd vccd vccd wire1609/X sky130_fd_sc_hd__buf_6
XFILLER_6_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4008 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2664 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__358__A _358_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_658 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2287 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__093__A _093_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3193 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_768 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input150_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2165_A wire2166/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input248_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input415_A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__268__A _268_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_524_ _524_/A _524_/B vssd vssd vccd vccd _524_/X sky130_fd_sc_hd__and2_4
XTAP_2742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_2029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_3727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_455_ _583_/A _455_/B _455_/C vssd vssd vccd vccd _455_/X sky130_fd_sc_hd__and3b_4
XTAP_2797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_386_ _514_/A _386_/B _386_/C vssd vssd vccd vccd _386_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__434__C _434_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1183 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1096 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4513 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output467_A wire1212/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3823 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1098_A wire1099/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__450__B _450_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output634_A _006_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3867 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1265_A _397_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4156 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output801_A _556_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1432_A wire1433/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_934 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput190 la_iena_mprj[37] vssd vssd vccd vccd _200_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__178__A _178_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_B split5/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1899_A wire1900/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput620 _109_/Y vssd vssd vccd vccd la_data_in_mprj[126] sky130_fd_sc_hd__buf_8
XFILLER_47_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput631 _003_/Y vssd vssd vccd vccd la_data_in_mprj[20] sky130_fd_sc_hd__buf_8
XFILLER_9_3552 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__360__B _360_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3311 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput642 _013_/Y vssd vssd vccd vccd la_data_in_mprj[30] sky130_fd_sc_hd__buf_8
XFILLER_43_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput653 _023_/Y vssd vssd vccd vccd la_data_in_mprj[40] sky130_fd_sc_hd__buf_8
XFILLER_47_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput664 _033_/Y vssd vssd vccd vccd la_data_in_mprj[50] sky130_fd_sc_hd__buf_8
XFILLER_28_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput675 _043_/Y vssd vssd vccd vccd la_data_in_mprj[60] sky130_fd_sc_hd__buf_8
XFILLER_5_3438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput686 _053_/Y vssd vssd vccd vccd la_data_in_mprj[70] sky130_fd_sc_hd__buf_8
Xwire2107 wire2108/X vssd vssd vccd vccd _576_/B sky130_fd_sc_hd__buf_6
XFILLER_29_2790 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput697 _063_/Y vssd vssd vccd vccd la_data_in_mprj[80] sky130_fd_sc_hd__buf_8
XFILLER_8_1115 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3208 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2118 wire2118/A vssd vssd vccd vccd _570_/B sky130_fd_sc_hd__buf_6
XFILLER_25_2643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2129 wire2129/A vssd vssd vccd vccd _562_/B sky130_fd_sc_hd__buf_6
XANTENNA_input3_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1406 _321_/X vssd vssd vccd vccd wire1406/X sky130_fd_sc_hd__buf_6
Xwire1417 wire1418/X vssd vssd vccd vccd wire1417/X sky130_fd_sc_hd__buf_6
XFILLER_47_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1428 wire1429/X vssd vssd vccd vccd wire1428/X sky130_fd_sc_hd__buf_6
XFILLER_23_3090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1439 _302_/X vssd vssd vccd vccd wire1439/X sky130_fd_sc_hd__buf_6
XFILLER_38_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__088__A _088_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3749 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_3148 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[13\]_B split4/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_240_ _240_/A _240_/B vssd vssd vccd vccd _240_/X sky130_fd_sc_hd__and2_2
XFILLER_32_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__535__B _535_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_171_ _171_/A _171_/B vssd vssd vccd vccd _171_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3624 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input198_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__551__A _551_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input365_A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2282_A wire2282/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__270__B _270_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[0\] user_irq_core[0] _291_/X vssd vssd vccd vccd _111_/A sky130_fd_sc_hd__nand2_2
XANTENNA_input59_A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3764 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1940 wire1940/A vssd vssd vccd vccd _196_/A sky130_fd_sc_hd__buf_6
XFILLER_4_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1951 wire1951/A vssd vssd vccd vccd _187_/A sky130_fd_sc_hd__buf_6
XFILLER_1_3869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1962 wire1962/A vssd vssd vccd vccd _180_/A sky130_fd_sc_hd__buf_6
Xwire1973 wire1973/A vssd vssd vccd vccd wire1973/X sky130_fd_sc_hd__buf_6
Xwire1984 wire1985/X vssd vssd vccd vccd _166_/A sky130_fd_sc_hd__buf_6
XFILLER_18_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1995 wire1996/X vssd vssd vccd vccd _623_/B sky130_fd_sc_hd__buf_6
XTAP_3251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_240 _256_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_251 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ _507_/A _507_/B vssd vssd vccd vccd _507_/X sky130_fd_sc_hd__and2_2
XANTENNA_262 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_273 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_284 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__445__B _445_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1013_A wire1014/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ _566_/A _438_/B _438_/C vssd vssd vccd vccd _438_/X sky130_fd_sc_hd__and3b_4
XANTENNA_output584_A wire1219/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_369_ _497_/A _369_/B _369_/C vssd vssd vccd vccd _369_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output751_A wire1187/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xrebuffer1 split4/A vssd vssd vccd vccd rebuffer1/X sky130_fd_sc_hd__bufbuf_8
XANTENNA_output849_A wire1417/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1382_A wire1383/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_893 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__180__B _180_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1931 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] wire1464/X vssd vssd vccd vccd _079_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3675 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1647_A wire1647/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1814_A wire1815/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_3285 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_2551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_753 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_701 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_789 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__355__B _355_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3988 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput472 wire1207/X vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__buf_8
XFILLER_47_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput483 _487_/X vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__buf_8
Xoutput494 wire1282/X vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__buf_8
XFILLER_9_2681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1203 _494_/X vssd vssd vccd vccd wire1203/X sky130_fd_sc_hd__buf_6
XFILLER_5_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1214 _470_/X vssd vssd vccd vccd wire1214/X sky130_fd_sc_hd__buf_6
XFILLER_25_2484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1225 _431_/X vssd vssd vccd vccd wire1225/X sky130_fd_sc_hd__buf_6
XFILLER_47_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1236 wire1237/X vssd vssd vccd vccd wire1236/X sky130_fd_sc_hd__buf_6
XFILLER_19_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1247 _415_/X vssd vssd vccd vccd wire1247/X sky130_fd_sc_hd__buf_6
XFILLER_5_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1258 _404_/X vssd vssd vccd vccd wire1258/X sky130_fd_sc_hd__buf_6
Xwire1269 _394_/X vssd vssd vccd vccd wire1269/X sky130_fd_sc_hd__buf_6
XFILLER_38_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2030_A wire2031/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input113_A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2128_A wire2128/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__A _546_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__265__B _265_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__451__A_N _579_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_223_ _223_/A _223_/B vssd vssd vccd vccd _223_/X sky130_fd_sc_hd__and2_2
XFILLER_23_491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_154_ _154_/A vssd vssd vccd vccd _154_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__281__A _281_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_085_ _085_/A vssd vssd vccd vccd _085_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_49_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3951 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3995 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_395 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1770 wire1771/X vssd vssd vccd vccd _385_/B sky130_fd_sc_hd__buf_6
XFILLER_4_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1781 wire1781/A vssd vssd vccd vccd wire1781/X sky130_fd_sc_hd__buf_6
XFILLER_53_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1792 wire1792/A vssd vssd vccd vccd wire1792/X sky130_fd_sc_hd__buf_6
XFILLER_20_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1130_A wire1130/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1228_A _428_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output799_A wire1152/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__175__B _175_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1031 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] _174_/X vssd vssd vccd vccd _158_/A
+ sky130_fd_sc_hd__nand2_2
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] rebuffer3/X vssd vssd vccd vccd _138_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_50_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1597_A wire1598/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__191__A _191_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1764_A wire1765/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2760 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_3419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] _285_/X vssd vssd vccd vccd wire1140/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_1046 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__A_N _602_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__366__A _366_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_586 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_737 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_rebuffer1_A split4/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3752 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2078_A wire2079/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1000 wire1001/X vssd vssd vccd vccd wire999/A sky130_fd_sc_hd__buf_6
XFILLER_40_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1011 wire1012/X vssd vssd vccd vccd wire1011/X sky130_fd_sc_hd__buf_6
XFILLER_25_2270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1022 wire1023/X vssd vssd vccd vccd wire1022/X sky130_fd_sc_hd__buf_6
XANTENNA_input230_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1033 wire1034/X vssd vssd vccd vccd wire1033/X sky130_fd_sc_hd__buf_6
XANTENNA_input328_A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1044 wire1045/X vssd vssd vccd vccd wire1044/X sky130_fd_sc_hd__buf_6
XANTENNA_wire2245_A wire2245/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3892 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1055 _127_/Y vssd vssd vccd vccd wire1055/X sky130_fd_sc_hd__buf_6
XFILLER_2_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1066 wire1067/X vssd vssd vccd vccd wire1066/X sky130_fd_sc_hd__buf_6
Xwire1077 wire1078/X vssd vssd vccd vccd wire1077/X sky130_fd_sc_hd__buf_8
Xwire1088 wire1089/X vssd vssd vccd vccd wire1088/X sky130_fd_sc_hd__buf_6
Xwire1099 wire1100/X vssd vssd vccd vccd wire1099/X sky130_fd_sc_hd__buf_6
XFILLER_28_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__276__A _276_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4364 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_973 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_206_ _206_/A _206_/B vssd vssd vccd vccd _206_/X sky130_fd_sc_hd__and2_4
XFILLER_10_3273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_137_ _137_/A vssd vssd vccd vccd _137_/Y sky130_fd_sc_hd__inv_12
XFILLER_8_999 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__442__C _442_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_068_ _068_/A vssd vssd vccd vccd _068_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_2594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output547_A wire1227/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1080_A _122_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1178_A _519_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output714_A _079_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1345_A _355_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2290 wire2290/A vssd vssd vccd vccd wire2290/X sky130_fd_sc_hd__buf_6
XFILLER_39_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] _222_/X vssd vssd vccd vccd _042_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_306 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1090 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3496 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__186__A _186_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_3140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1881_A wire1882/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1979_A wire1979/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire965_A _146_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[5\]_B split4/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2695 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__096__A _096_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_4504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1882 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_914 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input180_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2195_A wire2196/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input278_A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1167 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3077 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input445_A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input41_A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2150 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_851 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__437__C _437_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output497_A wire1279/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_4058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__453__B _453_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output664_A _033_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1295_A wire1296/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output831_A _583_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output929_A wire1323/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3202 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__363__B _363_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_939 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__B _538_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_540_ _540_/A _540_/B vssd vssd vccd vccd _540_/X sky130_fd_sc_hd__and2_4
XTAP_2913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_4069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_471_ _599_/A _471_/B _471_/C vssd vssd vccd vccd _471_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2110_A wire2110/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2208_A wire2208/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__554__A _554_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input395_A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input89_A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput350 la_oenb_mprj[66] vssd vssd vccd vccd wire1706/A sky130_fd_sc_hd__buf_6
XFILLER_23_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xinput361 la_oenb_mprj[76] vssd vssd vccd vccd wire1696/A sky130_fd_sc_hd__buf_6
Xinput372 la_oenb_mprj[86] vssd vssd vccd vccd wire1686/A sky130_fd_sc_hd__buf_6
XFILLER_40_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput383 la_oenb_mprj[96] vssd vssd vccd vccd wire1683/A sky130_fd_sc_hd__buf_6
XFILLER_48_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput394 mprj_adr_o_core[15] vssd vssd vccd vccd wire1662/A sky130_fd_sc_hd__buf_6
XFILLER_53_4103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4114 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__448__B _448_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1043_A wire1044/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output781_A _537_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1308_A wire1309/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output879_A wire1420/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_3132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__183__B _183_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1677_A wire1678/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput802 wire1195/X vssd vssd vccd vccd la_oenb_core[5] sky130_fd_sc_hd__buf_8
Xoutput813 wire1194/X vssd vssd vccd vccd la_oenb_core[6] sky130_fd_sc_hd__buf_8
Xoutput824 wire1193/X vssd vssd vccd vccd la_oenb_core[7] sky130_fd_sc_hd__buf_8
Xoutput835 wire1192/X vssd vssd vccd vccd la_oenb_core[8] sky130_fd_sc_hd__buf_8
XFILLER_6_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput846 wire1191/X vssd vssd vccd vccd la_oenb_core[9] sky130_fd_sc_hd__buf_8
XFILLER_29_3695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput857 wire1403/X vssd vssd vccd vccd mprj_adr_o_user[18] sky130_fd_sc_hd__buf_8
XANTENNA_wire1844_A wire1845/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput868 _333_/X vssd vssd vccd vccd mprj_adr_o_user[28] sky130_fd_sc_hd__buf_8
XFILLER_42_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_4012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput879 wire1420/X vssd vssd vccd vccd mprj_adr_o_user[9] sky130_fd_sc_hd__buf_8
XTAP_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_604 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2593 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2676 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__358__B _358_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2965 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_2244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_559 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2554 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2060_A wire2061/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input143_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2158_A wire2159/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__549__A _549_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__268__B _268_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input310_A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1992 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input408_A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_523_ _523_/A _523_/B vssd vssd vccd vccd _523_/X sky130_fd_sc_hd__and2_4
XTAP_3488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3864 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3886 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_454_ _582_/A _454_/B _454_/C vssd vssd vccd vccd _454_/X sky130_fd_sc_hd__and3b_4
XFILLER_32_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__284__A _284_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_191 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_385_ _513_/A _385_/B _385_/C vssd vssd vccd vccd _385_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_4197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1140 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1042 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1649 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__450__C _450_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3879 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output627_A _000_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1160_A wire1161/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1258_A _404_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput180 la_iena_mprj[28] vssd vssd vccd vccd wire1743/A sky130_fd_sc_hd__buf_6
XFILLER_42_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput191 la_iena_mprj[38] vssd vssd vccd vccd _201_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__178__B _178_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1425_A _311_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] _204_/X vssd vssd vccd vccd _024_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_33_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3221 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__194__A _194_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1794_A wire1795/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1874 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1104 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1961_A wire1961/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput610 _100_/Y vssd vssd vccd vccd la_data_in_mprj[117] sky130_fd_sc_hd__buf_8
Xoutput621 _110_/Y vssd vssd vccd vccd la_data_in_mprj[127] sky130_fd_sc_hd__buf_8
Xoutput632 _004_/Y vssd vssd vccd vccd la_data_in_mprj[21] sky130_fd_sc_hd__buf_8
XFILLER_47_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput643 _014_/Y vssd vssd vccd vccd la_data_in_mprj[31] sky130_fd_sc_hd__buf_8
XFILLER_9_3564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3323 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput654 _024_/Y vssd vssd vccd vccd la_data_in_mprj[41] sky130_fd_sc_hd__buf_8
XFILLER_5_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput665 _034_/Y vssd vssd vccd vccd la_data_in_mprj[51] sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] _166_/X vssd vssd vccd vccd _150_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput676 _044_/Y vssd vssd vccd vccd la_data_in_mprj[61] sky130_fd_sc_hd__buf_8
XFILLER_28_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput687 _054_/Y vssd vssd vccd vccd la_data_in_mprj[71] sky130_fd_sc_hd__buf_8
Xwire2108 wire2108/A vssd vssd vccd vccd wire2108/X sky130_fd_sc_hd__buf_6
XFILLER_25_2633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput698 _064_/Y vssd vssd vccd vccd la_data_in_mprj[81] sky130_fd_sc_hd__buf_8
Xwire2119 wire2120/X vssd vssd vccd vccd _569_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1127 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1407 _320_/X vssd vssd vccd vccd wire1407/X sky130_fd_sc_hd__buf_6
Xwire1418 wire1419/X vssd vssd vccd vccd wire1418/X sky130_fd_sc_hd__buf_6
Xwire1429 _304_/X vssd vssd vccd vccd wire1429/X sky130_fd_sc_hd__buf_6
XTAP_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3990 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2495 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_4153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_170_ _170_/A _170_/B vssd vssd vccd vccd _170_/X sky130_fd_sc_hd__and2_4
XFILLER_32_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_389 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__551__B _551_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input260_A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2275_A wire2276/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input358_A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_566 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__380__A_N _508_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__279__A _279_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1930 wire1930/A vssd vssd vccd vccd _334_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3776 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1941 wire1941/A vssd vssd vccd vccd _195_/A sky130_fd_sc_hd__buf_6
Xwire1952 wire1952/A vssd vssd vccd vccd _186_/A sky130_fd_sc_hd__buf_6
XFILLER_19_935 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1963 wire1964/X vssd vssd vccd vccd _179_/A sky130_fd_sc_hd__buf_6
Xwire1974 wire1974/A vssd vssd vccd vccd _173_/A sky130_fd_sc_hd__buf_6
XFILLER_20_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1985 wire1985/A vssd vssd vccd vccd wire1985/X sky130_fd_sc_hd__buf_6
XFILLER_19_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1996 wire1997/X vssd vssd vccd vccd wire1996/X sky130_fd_sc_hd__buf_6
XFILLER_19_979 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_230 wire2235/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_241 wire1989/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_506_ _506_/A _506_/B vssd vssd vccd vccd _506_/X sky130_fd_sc_hd__and2_2
XANTENNA_252 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1847 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_437_ _565_/A _437_/B _437_/C vssd vssd vccd vccd _437_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__445__C _445_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_368_ _368_/A _368_/B vssd vssd vccd vccd _368_/X sky130_fd_sc_hd__and2_2
XANTENNA_wire1006_A wire1007/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output577_A _457_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_299_ _299_/A _299_/B vssd vssd vccd vccd _299_/X sky130_fd_sc_hd__and2_4
Xrebuffer2 split4/A vssd vssd vccd vccd rebuffer2/X sky130_fd_sc_hd__bufbuf_8
XFILLER_31_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__461__B _461_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output744_A _619_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2021 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1375_A _345_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] wire1470/X vssd vssd vccd vccd _072_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_output911_A wire1076/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3687 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1542_A wire1543/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__189__A _189_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1002 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_2602 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1013 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1807_A wire1807/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire995_A wire996/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_459 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_4119 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__B _371_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput473 _478_/X vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__buf_8
Xoutput484 _488_/X vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__buf_8
XFILLER_43_2029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput495 wire1281/X vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__buf_8
XFILLER_25_2441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1204 _493_/X vssd vssd vccd vccd wire1204/X sky130_fd_sc_hd__buf_6
XFILLER_40_2939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__099__A _099_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1215 _469_/X vssd vssd vccd vccd wire1215/X sky130_fd_sc_hd__buf_6
Xwire1226 _430_/X vssd vssd vccd vccd wire1226/X sky130_fd_sc_hd__buf_6
XFILLER_9_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1237 _423_/X vssd vssd vccd vccd wire1237/X sky130_fd_sc_hd__buf_6
XFILLER_47_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1248 _414_/X vssd vssd vccd vccd wire1248/X sky130_fd_sc_hd__buf_6
XFILLER_47_57 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1259 _403_/X vssd vssd vccd vccd wire1259/X sky130_fd_sc_hd__buf_6
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_754 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__546__B _546_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2023_A wire2024/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3878 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_222_ _222_/A _222_/B vssd vssd vccd vccd _222_/X sky130_fd_sc_hd__and2_2
XFILLER_8_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__562__A _562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3444 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_153_ _153_/A vssd vssd vccd vccd _153_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__281__B _281_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input71_A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_084_ _084_/A vssd vssd vccd vccd _084_/Y sky130_fd_sc_hd__inv_4
XFILLER_45_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3963 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_4313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4493 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1491 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1760 wire1760/A vssd vssd vccd vccd _391_/B sky130_fd_sc_hd__buf_6
Xwire1771 wire1771/A vssd vssd vccd vccd wire1771/X sky130_fd_sc_hd__buf_6
Xwire1782 wire1783/X vssd vssd vccd vccd _380_/B sky130_fd_sc_hd__buf_6
XFILLER_18_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1793 wire1794/X vssd vssd vccd vccd _375_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_735 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__456__B _456_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1043 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output861_A _326_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1087 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] load_slew1458/X vssd vssd vccd vccd _131_/A
+ sky130_fd_sc_hd__nand2_8
XANTENNA_wire1492_A wire1493/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__191__B _191_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1924_A wire1924/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] _278_/X vssd vssd vccd vccd _098_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_39_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__366__B _366_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_B wire1465/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1001 _138_/Y vssd vssd vccd vccd wire1001/X sky130_fd_sc_hd__buf_6
Xwire1012 wire1013/X vssd vssd vccd vccd wire1012/X sky130_fd_sc_hd__buf_6
XFILLER_22_3860 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1023 wire1024/X vssd vssd vccd vccd wire1023/X sky130_fd_sc_hd__buf_6
Xwire1034 wire1035/X vssd vssd vccd vccd wire1034/X sky130_fd_sc_hd__buf_6
XFILLER_43_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3965 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1045 _129_/Y vssd vssd vccd vccd wire1045/X sky130_fd_sc_hd__buf_6
XFILLER_21_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1056 wire1057/X vssd vssd vccd vccd wire1056/X sky130_fd_sc_hd__buf_6
XFILLER_5_2398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1067 wire1068/X vssd vssd vccd vccd wire1067/X sky130_fd_sc_hd__buf_6
XFILLER_2_3987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2140_A wire2140/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input223_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1078 wire1079/X vssd vssd vccd vccd wire1078/X sky130_fd_sc_hd__buf_8
XANTENNA_wire2238_A wire2238/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1089 wire1090/X vssd vssd vccd vccd wire1089/X sky130_fd_sc_hd__buf_6
XANTENNA__557__A _557_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__276__B _276_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3631 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[86\]_B wire1473/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__292__A _292_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_205_ _205_/A _205_/B vssd vssd vccd vccd _205_/X sky130_fd_sc_hd__and2_4
XFILLER_12_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_136_ _136_/A vssd vssd vccd vccd _136_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_7_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4450 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_067_ _067_/A vssd vssd vccd vccd _067_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_45_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1073_A wire1074/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2280 wire2280/A vssd vssd vccd vccd _445_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1240_A wire1241/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2291 wire2291/A vssd vssd vccd vccd _436_/B sky130_fd_sc_hd__buf_6
XANTENNA_wire1338_A wire1339/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2407 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1590 wire1591/X vssd vssd vccd vccd wire1590/X sky130_fd_sc_hd__buf_6
XFILLER_4_1185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__186__B _186_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1505_A wire1506/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_B wire1482/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1874_A wire1874/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1062 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1647 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__441__A_N _569_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_2591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2549 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1594 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3826 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4240 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2090_A wire2091/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input173_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2188_A wire2189/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1179 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3911 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3955 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input340_A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input438_A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1737 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input34_A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__287__A _287_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3704 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2938 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__453__C _453_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1057 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_2679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output657_A _027_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_119_ _119_/A vssd vssd vccd vccd _119_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1190_A _507_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4100 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1288_A _375_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__464__A_N _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output824_A wire1193/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1455_A _296_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1203 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] _234_/X vssd vssd vccd vccd _054_/A
+ sky130_fd_sc_hd__nand2_4
XTAP_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1175 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1028 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_4505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1622_A wire1623/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__197__A _197_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3214 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1525 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_351 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_2579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1466 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_470_ _598_/A _470_/B _470_/C vssd vssd vccd vccd _470_/X sky130_fd_sc_hd__and3b_2
XTAP_2958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_535 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4368 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2103_A wire2104/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input290_A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input388_A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__487__A_N _615_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__570__A _570_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2428 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4431 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput340 la_oenb_mprj[57] vssd vssd vccd vccd _554_/A sky130_fd_sc_hd__buf_6
XFILLER_2_4282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput351 la_oenb_mprj[67] vssd vssd vccd vccd wire1705/A sky130_fd_sc_hd__buf_6
Xinput362 la_oenb_mprj[77] vssd vssd vccd vccd wire1695/A sky130_fd_sc_hd__buf_6
XFILLER_49_977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput373 la_oenb_mprj[87] vssd vssd vccd vccd wire1685/A sky130_fd_sc_hd__buf_6
Xinput384 la_oenb_mprj[97] vssd vssd vccd vccd wire1682/A sky130_fd_sc_hd__buf_6
Xinput395 mprj_adr_o_core[16] vssd vssd vccd vccd wire1658/A sky130_fd_sc_hd__buf_6
XFILLER_40_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__448__C _448_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1036_A wire1037/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_599_ _599_/A _599_/B vssd vssd vccd vccd _599_/X sky130_fd_sc_hd__and2_4
XFILLER_43_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__B _464_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_B _279_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output774_A wire1171/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output941_A wire1379/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput803 wire1149/X vssd vssd vccd vccd la_oenb_core[60] sky130_fd_sc_hd__buf_8
XANTENNA_wire1572_A wire1573/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput814 _567_/X vssd vssd vccd vccd la_oenb_core[70] sky130_fd_sc_hd__buf_8
Xoutput825 _577_/X vssd vssd vccd vccd la_oenb_core[80] sky130_fd_sc_hd__buf_8
XFILLER_47_1805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput836 wire1146/X vssd vssd vccd vccd la_oenb_core[90] sky130_fd_sc_hd__buf_8
Xoutput847 wire961/X vssd vssd vccd vccd mprj_ack_i_core sky130_fd_sc_hd__buf_8
XFILLER_25_3527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput858 wire1402/X vssd vssd vccd vccd mprj_adr_o_user[19] sky130_fd_sc_hd__buf_8
XFILLER_25_2804 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_2973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput869 _334_/X vssd vssd vccd vccd mprj_adr_o_user[29] sky130_fd_sc_hd__buf_8
XFILLER_47_1849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[25\]_A mprj_dat_i_user[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4508 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__374__B _374_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[107\]_B _270_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1399 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2376 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3987 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1566 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2511 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2566 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1821 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_2347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1865 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_4124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__549__B _549_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2053_A wire2053/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input136_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_605 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_wb_dat_gates\[16\]_A mprj_dat_i_user[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_522_ _522_/A _522_/B vssd vssd vccd vccd _522_/X sky130_fd_sc_hd__and2_2
XTAP_2722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2220_A wire2221/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input303_A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__565__A _565_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_453_ _581_/A _453_/B _453_/C vssd vssd vccd vccd _453_/X sky130_fd_sc_hd__and3b_4
XTAP_2777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__284__B _284_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_384_ _512_/A _384_/B _384_/C vssd vssd vccd vccd _384_/X sky130_fd_sc_hd__and3b_4
XFILLER_35_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4515 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output522_A wire1255/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1101 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_741 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__459__B _459_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1153_A wire1154/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_3529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3468 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput170 la_iena_mprj[19] vssd vssd vccd vccd _182_/B sky130_fd_sc_hd__buf_4
XFILLER_23_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput181 la_iena_mprj[29] vssd vssd vccd vccd _192_/B sky130_fd_sc_hd__buf_4
XFILLER_4_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput192 la_iena_mprj[39] vssd vssd vccd vccd _202_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1320_A wire1321/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1418_A wire1419/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output891_A wire1021/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] _197_/X vssd vssd vccd vccd _017_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_14_3206 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_2641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3277 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__194__B _194_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1787_A wire1787/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3597 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1954_A wire1955/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput600 _091_/Y vssd vssd vccd vccd la_data_in_mprj[108] sky130_fd_sc_hd__buf_8
Xoutput611 _101_/Y vssd vssd vccd vccd la_data_in_mprj[118] sky130_fd_sc_hd__buf_8
Xoutput622 _159_/Y vssd vssd vccd vccd la_data_in_mprj[12] sky130_fd_sc_hd__buf_8
XFILLER_29_3471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput633 _005_/Y vssd vssd vccd vccd la_data_in_mprj[22] sky130_fd_sc_hd__buf_8
XFILLER_44_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput644 _015_/Y vssd vssd vccd vccd la_data_in_mprj[32] sky130_fd_sc_hd__buf_8
XFILLER_25_3335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput655 _025_/Y vssd vssd vccd vccd la_data_in_mprj[42] sky130_fd_sc_hd__buf_8
XFILLER_9_3576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput666 _035_/Y vssd vssd vccd vccd la_data_in_mprj[52] sky130_fd_sc_hd__buf_8
XFILLER_47_1646 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput677 _045_/Y vssd vssd vccd vccd la_data_in_mprj[62] sky130_fd_sc_hd__buf_8
XFILLER_29_2781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput688 _055_/Y vssd vssd vccd vccd la_data_in_mprj[72] sky130_fd_sc_hd__buf_8
Xwire2109 wire2110/X vssd vssd vccd vccd _575_/B sky130_fd_sc_hd__buf_6
XFILLER_45_2071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput699 _065_/Y vssd vssd vccd vccd la_data_in_mprj[82] sky130_fd_sc_hd__buf_8
XFILLER_3_3120 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1408 wire1409/X vssd vssd vccd vccd wire1408/X sky130_fd_sc_hd__buf_6
XFILLER_42_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1419 _315_/X vssd vssd vccd vccd wire1419/X sky130_fd_sc_hd__buf_6
XFILLER_45_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__369__B _369_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1773 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4029 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4452 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2785 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4338 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3762 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_2373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1650 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1071 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input253_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2170_A wire2170/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2268_A wire2269/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input420_A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1920 wire1920/A vssd vssd vccd vccd _250_/A sky130_fd_sc_hd__buf_6
Xwire1931 wire1931/A vssd vssd vccd vccd _232_/A sky130_fd_sc_hd__buf_6
XFILLER_1_3849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1942 wire1942/A vssd vssd vccd vccd _194_/A sky130_fd_sc_hd__buf_6
XFILLER_19_925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1953 wire1953/A vssd vssd vccd vccd _185_/A sky130_fd_sc_hd__buf_6
XFILLER_21_3788 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1964 wire1964/A vssd vssd vccd vccd wire1964/X sky130_fd_sc_hd__buf_6
XTAP_3220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1975 wire1975/A vssd vssd vccd vccd _172_/A sky130_fd_sc_hd__buf_6
XFILLER_19_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1986 wire1987/X vssd vssd vccd vccd _165_/A sky130_fd_sc_hd__buf_6
XFILLER_20_1329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_755 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1997 wire1997/A vssd vssd vccd vccd wire1997/X sky130_fd_sc_hd__buf_6
XFILLER_19_4352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_4363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_220 wire2085/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 wire2243/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_4396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_505_ _505_/A _505_/B vssd vssd vccd vccd _505_/X sky130_fd_sc_hd__and2_2
XTAP_2552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_242 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_275 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_436_ _564_/A _436_/B _436_/C vssd vssd vccd vccd _436_/X sky130_fd_sc_hd__and3b_4
XTAP_1862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2104 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_367_ _367_/A _367_/B vssd vssd vccd vccd _367_/X sky130_fd_sc_hd__and2_2
XFILLER_32_3873 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_2159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_298_ _298_/A _298_/B vssd vssd vccd vccd _298_/X sky130_fd_sc_hd__and2_1
XANTENNA_output472_A wire1207/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xrebuffer3 split5/A vssd vssd vccd vccd rebuffer3/X sky130_fd_sc_hd__bufbuf_8
XFILLER_9_199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3705 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output737_A _613_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1270_A _393_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1368_A wire1369/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4005 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output904_A wire970/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__189__B _189_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1902 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1058 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_950 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire988_A wire989/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2925 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3394 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__371__C _371_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1391 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3143 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput463 wire1294/X vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__buf_8
Xoutput474 wire1284/X vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__buf_8
Xoutput485 wire1283/X vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__buf_8
Xoutput496 wire1280/X vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__buf_8
XFILLER_9_2683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1205 _492_/X vssd vssd vccd vccd wire1205/X sky130_fd_sc_hd__buf_6
Xwire1216 _468_/X vssd vssd vccd vccd wire1216/X sky130_fd_sc_hd__buf_6
XFILLER_5_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1227 _429_/X vssd vssd vccd vccd wire1227/X sky130_fd_sc_hd__buf_6
XFILLER_5_2569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1238 wire1239/X vssd vssd vccd vccd wire1238/X sky130_fd_sc_hd__buf_6
XFILLER_38_4227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1249 _413_/X vssd vssd vccd vccd wire1249/X sky130_fd_sc_hd__buf_6
XFILLER_5_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_4561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_69 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2260 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_703 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2279 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2016_A wire2017/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_994 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_221_ _221_/A _221_/B vssd vssd vccd vccd _221_/X sky130_fd_sc_hd__and2_2
XFILLER_14_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_152_ _152_/A vssd vssd vccd vccd _152_/Y sky130_fd_sc_hd__inv_2
XANTENNA__562__B _562_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3456 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_083_ _083_/A vssd vssd vccd vccd _083_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input370_A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_input64_A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_821 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_320 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_3975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4231 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_load_slew1458_A split5/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2002 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1750 wire1750/A vssd vssd vccd vccd _452_/C sky130_fd_sc_hd__buf_6
XFILLER_18_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1761 wire1761/A vssd vssd vccd vccd _390_/B sky130_fd_sc_hd__buf_6
XFILLER_19_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1772 wire1773/X vssd vssd vccd vccd _303_/A sky130_fd_sc_hd__buf_6
Xwire1783 wire1783/A vssd vssd vccd vccd wire1783/X sky130_fd_sc_hd__buf_6
XFILLER_37_3025 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1794 wire1795/X vssd vssd vccd vccd wire1794/X sky130_fd_sc_hd__buf_6
XTAP_3050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__456__C _456_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1116_A wire1117/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output687_A _054_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_419_ _547_/A _419_/B _419_/C vssd vssd vccd vccd _419_/X sky130_fd_sc_hd__and3b_4
XTAP_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1689 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__472__B _472_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1099 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output854_A wire1407/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1485_A input96/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1652_A wire1653/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_3474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3316 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3134 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] _271_/X vssd vssd vccd vccd _091_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_17_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__370__A_N _498_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__382__B _382_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2799 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3191 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[8\]_A mprj_dat_i_user[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmax_length1714 _416_/A_N vssd vssd vccd vccd wire1713/A sky130_fd_sc_hd__buf_6
XFILLER_49_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1002 wire1003/X vssd vssd vccd vccd wire1002/X sky130_fd_sc_hd__buf_6
XFILLER_5_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1013 wire1014/X vssd vssd vccd vccd wire1013/X sky130_fd_sc_hd__buf_6
XFILLER_22_3872 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1024 wire1025/X vssd vssd vccd vccd wire1024/X sky130_fd_sc_hd__buf_6
XFILLER_5_2366 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1035 _131_/Y vssd vssd vccd vccd wire1035/X sky130_fd_sc_hd__buf_6
Xwire1046 wire1047/X vssd vssd vccd vccd wire1046/X sky130_fd_sc_hd__buf_6
XFILLER_38_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1057 wire1058/X vssd vssd vccd vccd wire1057/X sky130_fd_sc_hd__buf_6
XFILLER_5_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1068 wire1069/X vssd vssd vccd vccd wire1068/X sky130_fd_sc_hd__buf_6
XFILLER_1_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3999 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1079 wire1080/X vssd vssd vccd vccd wire1079/X sky130_fd_sc_hd__buf_6
XANTENNA__557__B _557_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input216_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3643 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2300_A wire2300/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__573__A _573_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3698 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4090 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_204_ _204_/A _204_/B vssd vssd vccd vccd _204_/X sky130_fd_sc_hd__and2_4
XFILLER_12_975 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3220 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_3231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_135_ _135_/A vssd vssd vccd vccd _135_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_49_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_066_ _066_/A vssd vssd vccd vccd _066_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4462 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3603 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1066_A wire1067/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2270 wire2270/A vssd vssd vccd vccd wire2270/X sky130_fd_sc_hd__buf_6
Xwire2281 wire2281/A vssd vssd vccd vccd _309_/A sky130_fd_sc_hd__buf_6
XFILLER_1_3454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire2292 wire2292/A vssd vssd vccd vccd _435_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1580 wire1581/X vssd vssd vccd vccd wire1580/X sky130_fd_sc_hd__buf_6
XANTENNA__467__B _467_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1591 wire1591/A vssd vssd vccd vccd wire1591/X sky130_fd_sc_hd__buf_6
XFILLER_0_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__393__A_N _521_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1400_A wire1401/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1306 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1867_A wire1868/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1930 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__B _377_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3529 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_3838 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3540 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_4296 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3584 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3035 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2301 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input166_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2083_A wire2083/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3967 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input333_A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_698 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3680 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__568__A _568_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input27_A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1833 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__287__B _287_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_1276 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_4130 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3738 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4038 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_3397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4535 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_118_ _118_/A vssd vssd vccd vccd _118_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_29_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output552_A _434_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4112 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_049_ _049_/A vssd vssd vccd vccd _049_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3889 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1183_A _514_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_3641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3591 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output817_A _570_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1350_A wire1351/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1448_A _300_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1259 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] _227_/X vssd vssd vccd vccd _047_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_1187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1615_A wire1616/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3805 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3106 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3226 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2514 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_897 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1984_A wire1985/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire970_A wire971/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1158 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1423 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1920 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2518 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1986 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_4306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2325 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_3638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4336 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_547 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input283_A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_3392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2298_A wire2298/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__B _570_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1091 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_4443 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1007 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3972 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xsplit4 split4/A vssd vssd vccd vccd split4/X sky130_fd_sc_hd__buf_8
XFILLER_40_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput330 la_oenb_mprj[48] vssd vssd vccd vccd _545_/A sky130_fd_sc_hd__buf_8
XFILLER_2_4261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__298__A _298_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput341 la_oenb_mprj[58] vssd vssd vccd vccd wire1711/A sky130_fd_sc_hd__buf_6
XFILLER_48_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput352 la_oenb_mprj[68] vssd vssd vccd vccd wire1704/A sky130_fd_sc_hd__buf_6
Xinput363 la_oenb_mprj[78] vssd vssd vccd vccd _447_/A_N sky130_fd_sc_hd__buf_6
Xinput374 la_oenb_mprj[88] vssd vssd vccd vccd wire1684/A sky130_fd_sc_hd__buf_6
XFILLER_29_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput385 la_oenb_mprj[98] vssd vssd vccd vccd wire1681/A sky130_fd_sc_hd__buf_6
XFILLER_48_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput396 mprj_adr_o_core[17] vssd vssd vccd vccd wire1654/A sky130_fd_sc_hd__buf_6
XFILLER_35_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3524 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2714 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_374 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1029_A wire1030/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_598_ _598_/A _598_/B vssd vssd vccd vccd _598_/X sky130_fd_sc_hd__and2_4
XFILLER_32_834 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__C _464_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__431__A_N _559_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output767_A wire1173/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1398_A wire1399/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__480__B _480_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4207 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1 la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput804 wire1148/X vssd vssd vccd vccd la_oenb_core[61] sky130_fd_sc_hd__buf_8
XANTENNA_output934_A wire1303/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput815 _568_/X vssd vssd vccd vccd la_oenb_core[71] sky130_fd_sc_hd__buf_8
Xoutput826 _578_/X vssd vssd vccd vccd la_oenb_core[81] sky130_fd_sc_hd__buf_8
XFILLER_42_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput837 wire1145/X vssd vssd vccd vccd la_oenb_core[91] sky130_fd_sc_hd__buf_8
XFILLER_6_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1565_A wire1566/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput848 _305_/X vssd vssd vccd vccd mprj_adr_o_user[0] sky130_fd_sc_hd__buf_8
XFILLER_28_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput859 _306_/X vssd vssd vccd vccd mprj_adr_o_user[1] sky130_fd_sc_hd__buf_8
XFILLER_42_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3302 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[25\]_B split5/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__001__A _001_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_2300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__374__C _374_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2388 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__390__B _390_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_3185 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2523 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_wb_dat_gates\[16\]_B load_slew1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2046_A wire2046/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input129_A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_521_ _521_/A _521_/B vssd vssd vccd vccd _521_/X sky130_fd_sc_hd__and2_4
XTAP_2723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_4100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__565__B _565_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_452_ _580_/A _452_/B _452_/C vssd vssd vccd vccd _452_/X sky130_fd_sc_hd__and3b_4
XFILLER_17_4280 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2213_A wire2214/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__454__A_N _582_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4144 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_383_ _511_/A _383_/B _383_/C vssd vssd vccd vccd _383_/X sky130_fd_sc_hd__and3b_4
XFILLER_50_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input94_A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4480 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__A _581_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1271 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output515_A wire1262/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput160 la_iena_mprj[125] vssd vssd vccd vccd _288_/B sky130_fd_sc_hd__buf_4
XFILLER_4_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput171 la_iena_mprj[1] vssd vssd vccd vccd _164_/B sky130_fd_sc_hd__clkbuf_4
Xinput182 la_iena_mprj[2] vssd vssd vccd vccd _165_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput193 la_iena_mprj[3] vssd vssd vccd vccd _166_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1146_A _587_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_4044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3343 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__475__B _475_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1313_A wire1314/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output884_A wire1056/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] _190_/X vssd vssd vccd vccd _010_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_18_2664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2577 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4212 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3500 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput601 _092_/Y vssd vssd vccd vccd la_data_in_mprj[109] sky130_fd_sc_hd__buf_8
Xoutput612 _102_/Y vssd vssd vccd vccd la_data_in_mprj[119] sky130_fd_sc_hd__buf_8
XFILLER_25_3303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput623 _160_/Y vssd vssd vccd vccd la_data_in_mprj[13] sky130_fd_sc_hd__buf_8
Xoutput634 _006_/Y vssd vssd vccd vccd la_data_in_mprj[23] sky130_fd_sc_hd__buf_8
Xoutput645 _016_/Y vssd vssd vccd vccd la_data_in_mprj[33] sky130_fd_sc_hd__buf_8
XFILLER_47_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput656 _026_/Y vssd vssd vccd vccd la_data_in_mprj[43] sky130_fd_sc_hd__buf_8
Xoutput667 _036_/Y vssd vssd vccd vccd la_data_in_mprj[53] sky130_fd_sc_hd__buf_8
XFILLER_9_3588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2613 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput678 _046_/Y vssd vssd vccd vccd la_data_in_mprj[63] sky130_fd_sc_hd__buf_8
Xoutput689 _056_/Y vssd vssd vccd vccd la_data_in_mprj[73] sky130_fd_sc_hd__buf_8
XFILLER_42_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1409 _319_/X vssd vssd vccd vccd wire1409/X sky130_fd_sc_hd__buf_6
XFILLER_3_3143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__369__C _369_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__477__A_N _605_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__385__B _385_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_4420 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4464 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2797 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_513 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2375 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input246_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2163_A wire2164/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_split4_A split4/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3975 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1910 wire1910/A vssd vssd vccd vccd wire1910/X sky130_fd_sc_hd__buf_6
Xwire1921 wire1921/A vssd vssd vccd vccd _249_/A sky130_fd_sc_hd__buf_6
XFILLER_41_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1932 wire1932/A vssd vssd vccd vccd _231_/A sky130_fd_sc_hd__buf_6
XFILLER_46_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1943 wire1943/A vssd vssd vccd vccd _193_/A sky130_fd_sc_hd__buf_6
Xwire1954 wire1955/X vssd vssd vccd vccd _184_/A sky130_fd_sc_hd__buf_6
XTAP_3210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1965 wire1966/X vssd vssd vccd vccd _178_/A sky130_fd_sc_hd__buf_6
XTAP_3221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input413_A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1976 wire1976/A vssd vssd vccd vccd _171_/A sky130_fd_sc_hd__buf_6
XTAP_3232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1987 wire1987/A vssd vssd vccd vccd wire1987/X sky130_fd_sc_hd__buf_6
XANTENNA__576__A _576_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1998 wire1999/X vssd vssd vccd vccd _622_/B sky130_fd_sc_hd__buf_6
XFILLER_41_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _574_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 wire2093/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__295__B _295_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_504_ _504_/A _504_/B vssd vssd vccd vccd _504_/X sky130_fd_sc_hd__and2_2
XANTENNA_232 _440_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 _351_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3696 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_435_ _563_/A _435_/B _435_/C vssd vssd vccd vccd _435_/X sky130_fd_sc_hd__and3b_4
XANTENNA_287 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_366_ _366_/A _366_/B vssd vssd vccd vccd _366_/X sky130_fd_sc_hd__and2_2
XFILLER_31_2127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_297_ _297_/A _297_/B vssd vssd vccd vccd _297_/X sky130_fd_sc_hd__and2_4
XFILLER_48_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_189 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output465_A wire1214/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1096_A wire1097/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output632_A _004_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_3667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1427 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2966 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_2690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1430_A wire1431/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1528_A wire1528/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1037 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_406 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1897_A wire1898/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2937 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4064 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_3352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput464 wire1215/X vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput475 _479_/X vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__buf_8
XFILLER_9_2651 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput486 _489_/X vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__buf_8
XFILLER_25_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput497 wire1279/X vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__buf_8
XFILLER_5_3249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_3199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input1_A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1206 _491_/X vssd vssd vccd vccd wire1206/X sky130_fd_sc_hd__buf_6
XFILLER_47_15 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1217 _465_/X vssd vssd vccd vccd wire1217/X sky130_fd_sc_hd__buf_6
Xwire1228 _428_/X vssd vssd vccd vccd wire1228/X sky130_fd_sc_hd__buf_6
XFILLER_41_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1239 _422_/X vssd vssd vccd vccd wire1239/X sky130_fd_sc_hd__buf_6
XFILLER_28_701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2272 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_715 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_3749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_220_ _220_/A _220_/B vssd vssd vccd vccd _220_/X sky130_fd_sc_hd__and2_2
XFILLER_49_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2009_A wire2009/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_151_ _151_/A vssd vssd vccd vccd _151_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input196_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_082_ _082_/A vssd vssd vccd vccd _082_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2280_A wire2280/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input363_A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_332 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input57_A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4243 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2014 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1460 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3553 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1740 input21/X vssd vssd vccd vccd _484_/C sky130_fd_sc_hd__buf_6
XFILLER_1_2913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_2069 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1751 wire1751/A vssd vssd vccd vccd _451_/C sky130_fd_sc_hd__buf_6
XFILLER_1_2924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1762 wire1763/X vssd vssd vccd vccd _389_/B sky130_fd_sc_hd__buf_6
XFILLER_46_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1773 wire1773/A vssd vssd vccd vccd wire1773/X sky130_fd_sc_hd__buf_6
XFILLER_1_2946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1784 wire1785/X vssd vssd vccd vccd _379_/B sky130_fd_sc_hd__buf_6
XTAP_3040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1795 wire1795/A vssd vssd vccd vccd wire1795/X sky130_fd_sc_hd__buf_6
XTAP_3051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_4014 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_4047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2060 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_418_ _546_/A _418_/B _418_/C vssd vssd vccd vccd _418_/X sky130_fd_sc_hd__and3b_4
XANTENNA_wire1011_A wire1012/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output582_A wire1221/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1109_A wire1110/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_349_ _349_/A _349_/B vssd vssd vccd vccd _349_/X sky130_fd_sc_hd__and2_4
XFILLER_35_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1245 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output847_A wire961/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_4121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1380_A wire1381/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1478_A _244_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3431 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] _257_/X vssd vssd vccd vccd _077_/A
+ sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1645_A wire1646/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1812_A wire1813/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_4125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2701 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_2881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2745 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_475 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3777 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_wb_dat_gates\[8\]_B max_cap1456/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2527 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2262 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_3079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1003 wire1004/X vssd vssd vccd vccd wire1003/X sky130_fd_sc_hd__buf_6
XFILLER_2_3923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1014 wire1015/X vssd vssd vccd vccd wire1014/X sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[8\]_B _171_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1025 _133_/Y vssd vssd vccd vccd wire1025/X sky130_fd_sc_hd__buf_6
XFILLER_25_2284 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1036 wire1037/X vssd vssd vccd vccd wire1036/X sky130_fd_sc_hd__buf_6
Xwire1047 wire1048/X vssd vssd vccd vccd wire1047/X sky130_fd_sc_hd__buf_6
XFILLER_5_2378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1058 wire1059/X vssd vssd vccd vccd wire1058/X sky130_fd_sc_hd__buf_6
Xwire1069 wire1070/X vssd vssd vccd vccd wire1069/X sky130_fd_sc_hd__buf_6
XFILLER_38_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1436 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input111_A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input209_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2126_A wire2126/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3655 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__573__B _573_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_203_ _203_/A _203_/B vssd vssd vccd vccd _203_/X sky130_fd_sc_hd__and2_4
XFILLER_19_1398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_134_ _134_/A vssd vssd vccd vccd _134_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3276 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_065_ _065_/A vssd vssd vccd vccd _065_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_49_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4474 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_151 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3795 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1314 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_4281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_3411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2260 wire2260/A vssd vssd vccd vccd wire2260/X sky130_fd_sc_hd__buf_6
XFILLER_43_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2271 wire2272/X vssd vssd vccd vccd _451_/B sky130_fd_sc_hd__buf_6
Xwire2282 wire2282/A vssd vssd vccd vccd _444_/B sky130_fd_sc_hd__buf_6
Xwire2293 wire2293/A vssd vssd vccd vccd _308_/A sky130_fd_sc_hd__buf_6
XANTENNA_wire1059_A wire1060/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1570 wire1571/X vssd vssd vccd vccd wire1570/X sky130_fd_sc_hd__buf_6
XFILLER_39_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1581 wire1581/A vssd vssd vccd vccd wire1581/X sky130_fd_sc_hd__buf_6
XANTENNA__467__C _467_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1592 wire1593/X vssd vssd vccd vccd _307_/B sky130_fd_sc_hd__buf_6
XFILLER_21_2693 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_4445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1226_A _430_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output797_A wire1155/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_4309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__B _483_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] split5/A vssd vssd vccd vccd _136_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_33_1318 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_773 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1595_A wire1596/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_2486 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1616 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1762_A wire1763/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3333 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__004__A _004_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_2435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] _283_/X vssd vssd vccd vccd wire1142/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_29_317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__C _377_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_810 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3920 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3806 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__393__B _393_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_283 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_3596 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire2076_A wire2077/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_4421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input159_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__568__B _568_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2243_A wire2243/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_3692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input326_A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1845 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4142 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__584__A _584_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_3430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4066 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1763 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_3474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2620 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2615 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2063 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2648 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_1985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_117_ _117_/A vssd vssd vccd vccd _117_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_2372 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_3857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_048_ _048_/A vssd vssd vccd vccd _048_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_4_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4124 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output545_A wire1228/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_4207 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_4168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1176_A _521_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2952 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_3697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output712_A _077_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__478__B _478_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1343_A wire1344/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2090 wire2091/X vssd vssd vccd vccd _584_/B sky130_fd_sc_hd__buf_6
XFILLER_26_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] _220_/X vssd vssd vccd vccd _040_/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_3817 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1510_A wire1510/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1608_A wire1609/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_17_2504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_504 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4117 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2715 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1977_A wire1978/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire963_A wire964/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1435 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1479 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2633 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2855 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__388__B _388_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3305 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_876 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4348 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_3073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2962 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3360 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1693 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2193_A wire2193/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input276_A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1980 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__383__A_N _511_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input443_A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3984 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3743 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4499 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__579__A _579_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3787 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xsplit5 split5/A vssd vssd vccd vccd split5/X sky130_fd_sc_hd__buf_8
XFILLER_48_401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput320 la_oenb_mprj[39] vssd vssd vccd vccd _536_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xinput331 la_oenb_mprj[49] vssd vssd vccd vccd _546_/A sky130_fd_sc_hd__buf_4
XFILLER_0_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput342 la_oenb_mprj[59] vssd vssd vccd vccd _556_/A sky130_fd_sc_hd__buf_6
XANTENNA__298__B _298_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput353 la_oenb_mprj[69] vssd vssd vccd vccd wire1703/A sky130_fd_sc_hd__buf_6
XFILLER_48_445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput364 la_oenb_mprj[79] vssd vssd vccd vccd wire1693/A sky130_fd_sc_hd__buf_6
Xinput375 la_oenb_mprj[89] vssd vssd vccd vccd _586_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput386 la_oenb_mprj[99] vssd vssd vccd vccd wire1680/A sky130_fd_sc_hd__buf_6
Xinput397 mprj_adr_o_core[18] vssd vssd vccd vccd wire1651/A sky130_fd_sc_hd__buf_6
XFILLER_48_489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_4139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_597_ _597_/A _597_/B vssd vssd vccd vccd _597_/X sky130_fd_sc_hd__and2_4
XFILLER_43_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_386 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_846 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output495_A wire1281/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2169 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4311 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output662_A _032_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__480__C _480_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2 la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1293_A _370_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4219 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput805 _559_/X vssd vssd vccd vccd la_oenb_core[62] sky130_fd_sc_hd__buf_8
XFILLER_47_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput816 _569_/X vssd vssd vccd vccd la_oenb_core[72] sky130_fd_sc_hd__buf_8
Xoutput827 _579_/X vssd vssd vccd vccd la_oenb_core[82] sky130_fd_sc_hd__buf_8
Xoutput838 _589_/X vssd vssd vccd vccd la_oenb_core[92] sky130_fd_sc_hd__buf_8
XFILLER_42_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output927_A wire1331/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput849 wire1417/X vssd vssd vccd vccd mprj_adr_o_user[10] sky130_fd_sc_hd__buf_8
XFILLER_6_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1460_A wire1461/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1558_A wire1559/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3297 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_3060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_2025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3625 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4061 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_194 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_2356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__390__C _390_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_520_ _520_/A _520_/B vssd vssd vccd vccd _520_/X sky130_fd_sc_hd__and2_4
XTAP_2702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3834 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2039_A wire2039/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_451_ _579_/A _451_/B _451_/C vssd vssd vccd vccd _451_/X sky130_fd_sc_hd__and3b_4
XFILLER_26_662 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_150 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_4292 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_382_ _510_/A _382_/B _382_/C vssd vssd vccd vccd _382_/X sky130_fd_sc_hd__and3b_4
XFILLER_15_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2206_A wire2207/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2489 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2770 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_input393_A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_349 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__B _581_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input87_A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1007 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3190 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4263 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__102__A _102_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3667 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput150 la_iena_mprj[116] vssd vssd vccd vccd _279_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput161 la_iena_mprj[126] vssd vssd vccd vccd _289_/B sky130_fd_sc_hd__buf_4
XFILLER_48_253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput172 la_iena_mprj[20] vssd vssd vccd vccd _183_/B sky130_fd_sc_hd__buf_4
XTAP_4660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput183 la_iena_mprj[30] vssd vssd vccd vccd _193_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_output508_A wire1269/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_3901 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput194 la_iena_mprj[40] vssd vssd vccd vccd _203_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3300 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_4693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1041_A wire1042/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1483 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3945 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__475__C _475_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_3355 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4201 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_3989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_3388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_643 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1306_A _366_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output877_A wire1423/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1877 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__491__B _491_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_4224 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1675_A wire1676/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_3512 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput602 _157_/Y vssd vssd vccd vccd la_data_in_mprj[10] sky130_fd_sc_hd__buf_8
XFILLER_9_4268 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput613 _158_/Y vssd vssd vccd vccd la_data_in_mprj[11] sky130_fd_sc_hd__buf_8
Xoutput624 _161_/Y vssd vssd vccd vccd la_data_in_mprj[14] sky130_fd_sc_hd__buf_8
XFILLER_29_3473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput635 _007_/Y vssd vssd vccd vccd la_data_in_mprj[24] sky130_fd_sc_hd__buf_8
Xoutput646 _017_/Y vssd vssd vccd vccd la_data_in_mprj[34] sky130_fd_sc_hd__buf_8
XFILLER_5_3409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput657 _027_/Y vssd vssd vccd vccd la_data_in_mprj[44] sky130_fd_sc_hd__buf_8
XFILLER_29_2761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1842_A wire1843/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput668 _037_/Y vssd vssd vccd vccd la_data_in_mprj[54] sky130_fd_sc_hd__buf_8
Xoutput679 _047_/Y vssd vssd vccd vccd la_data_in_mprj[64] sky130_fd_sc_hd__buf_8
XFILLER_29_2794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_905 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3108 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__385__C _385_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_4481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_4432 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3499 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3731 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4476 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_153 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3702 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3871 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2354 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2387 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1900 wire1900/A vssd vssd vccd vccd wire1900/X sky130_fd_sc_hd__buf_6
XANTENNA_input141_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1911 wire1911/A vssd vssd vccd vccd _259_/A sky130_fd_sc_hd__buf_6
XANTENNA_wire2156_A wire2156/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1922 wire1922/A vssd vssd vccd vccd _248_/A sky130_fd_sc_hd__buf_4
XANTENNA_input239_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1933 wire1933/A vssd vssd vccd vccd _230_/A sky130_fd_sc_hd__buf_4
XANTENNA__421__A_N _549_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1944 wire1944/A vssd vssd vccd vccd _330_/A sky130_fd_sc_hd__buf_6
XTAP_3200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1539 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1955 wire1955/A vssd vssd vccd vccd wire1955/X sky130_fd_sc_hd__buf_6
XTAP_3211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1966 wire1966/A vssd vssd vccd vccd wire1966/X sky130_fd_sc_hd__buf_6
XTAP_3222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1977 wire1978/X vssd vssd vccd vccd _170_/A sky130_fd_sc_hd__buf_6
XTAP_3233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1988 wire1989/X vssd vssd vccd vccd _164_/A sky130_fd_sc_hd__buf_6
XFILLER_45_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1999 wire2000/X vssd vssd vccd vccd wire1999/X sky130_fd_sc_hd__buf_6
XANTENNA__576__B _576_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input406_A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_200 _340_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _526_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_503_ _503_/A _503_/B vssd vssd vccd vccd _503_/X sky130_fd_sc_hd__and2_4
XTAP_2532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _438_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_993 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_244 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_429 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_266 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_434_ _562_/A _434_/B _434_/C vssd vssd vccd vccd _434_/X sky130_fd_sc_hd__and3b_4
XTAP_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1118 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2253 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__592__A _592_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _365_/A _365_/B vssd vssd vccd vccd _365_/X sky130_fd_sc_hd__and2_2
XFILLER_9_113 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2297 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_296_ _296_/A _296_/B vssd vssd vccd vccd _296_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_831 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_4347 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1089_A wire1090/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[40\]_B _203_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1345 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_2945 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1256_A _406_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__486__B _486_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1423_A _312_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3753 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_4031 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3948 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4032 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_3134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] _164_/X vssd vssd vccd vccd _148_/A
+ sky130_fd_sc_hd__nand2_1
Xoutput465 wire1214/X vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__buf_8
XFILLER_5_3217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[31\]_B _194_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput476 _480_/X vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__buf_8
XFILLER_44_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__444__A_N _572_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput487 _490_/X vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__buf_8
XFILLER_9_2663 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput498 wire1278/X vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__buf_8
XFILLER_25_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1207 _477_/X vssd vssd vccd vccd wire1207/X sky130_fd_sc_hd__buf_6
Xwire1218 _464_/X vssd vssd vccd vccd wire1218/X sky130_fd_sc_hd__buf_6
XFILLER_47_27 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1229 wire1230/X vssd vssd vccd vccd wire1229/X sky130_fd_sc_hd__buf_6
XFILLER_5_1837 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_223 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__396__B _396_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_2827 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[98\]_B _261_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_4104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2573 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2437 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_150_ _150_/A vssd vssd vccd vccd _150_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_657 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_081_ _081_/A vssd vssd vccd vccd _081_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input189_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire2273_A wire2274/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input356_A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3808 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3751 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2026 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__587__A _587_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3565 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1730 wire1730/A vssd vssd vccd vccd _614_/A sky130_fd_sc_hd__buf_6
XFILLER_1_2903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1741 input20/X vssd vssd vccd vccd _483_/C sky130_fd_sc_hd__buf_6
XFILLER_1_3659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1752 wire1752/A vssd vssd vccd vccd _450_/C sky130_fd_sc_hd__buf_6
Xwire1763 wire1763/A vssd vssd vccd vccd wire1763/X sky130_fd_sc_hd__buf_6
XFILLER_1_2936 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_3005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1774 wire1775/X vssd vssd vccd vccd _384_/B sky130_fd_sc_hd__buf_6
XTAP_3030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_757 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1785 wire1785/A vssd vssd vccd vccd wire1785/X sky130_fd_sc_hd__buf_6
XTAP_3041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_768 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xwire1796 wire1797/X vssd vssd vccd vccd _302_/A sky130_fd_sc_hd__buf_6
XTAP_3052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2969 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4184 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[89\]_B wire1470/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_3472 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3358 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_417_ _545_/A _417_/B _417_/C vssd vssd vccd vccd _417_/X sky130_fd_sc_hd__and3b_4
XTAP_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4395 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_3661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_348_ _348_/A _348_/B vssd vssd vccd vccd _348_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1004_A wire1005/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3082 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output575_A _455_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_279_ _279_/A _279_/B vssd vssd vccd vccd _279_/X sky130_fd_sc_hd__and2_4
XFILLER_48_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__467__A_N _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A _617_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1373_A wire1374/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] wire1472/X vssd vssd vccd vccd wire1128/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_29_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2043 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1540_A wire1541/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3250 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1638_A wire1639/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__497__A _497_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1805_A wire1805/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2385 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1734 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_4137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire993_A wire994/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4560 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2713 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4424 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2757 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3756 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1482 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_3193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2539 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2471 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2717 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1004 wire1005/X vssd vssd vccd vccd wire1004/X sky130_fd_sc_hd__buf_6
Xwire1015 _135_/Y vssd vssd vccd vccd wire1015/X sky130_fd_sc_hd__buf_6
Xwire1026 wire1027/X vssd vssd vccd vccd wire1026/X sky130_fd_sc_hd__buf_6
XFILLER_2_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1037 wire1038/X vssd vssd vccd vccd wire1037/X sky130_fd_sc_hd__buf_6
XFILLER_5_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1048 wire1049/X vssd vssd vccd vccd wire1048/X sky130_fd_sc_hd__buf_6
Xwire1059 wire1060/X vssd vssd vccd vccd wire1059/X sky130_fd_sc_hd__buf_6
XANTENNA__200__A _200_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_4059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1667 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2021_A wire2022/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input104_A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2119_A wire2120/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_782 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1989 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_202_ _202_/A _202_/B vssd vssd vccd vccd _202_/X sky130_fd_sc_hd__and2_4
XFILLER_23_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_133_ _133_/A vssd vssd vccd vccd _133_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_10_3255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2543 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3288 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_4431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_064_ _064_/A vssd vssd vccd vccd _064_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_3581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire2250 wire2250/A vssd vssd vccd vccd _459_/B sky130_fd_sc_hd__buf_6
Xwire2261 wire2261/A vssd vssd vccd vccd _310_/A sky130_fd_sc_hd__buf_6
XFILLER_40_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2272 wire2272/A vssd vssd vccd vccd wire2272/X sky130_fd_sc_hd__buf_6
XFILLER_43_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2283 wire2283/A vssd vssd vccd vccd _443_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2294 wire2294/A vssd vssd vccd vccd _434_/B sky130_fd_sc_hd__buf_6
XFILLER_47_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1560 wire1561/X vssd vssd vccd vccd _312_/B sky130_fd_sc_hd__buf_6
Xwire1571 wire1571/A vssd vssd vccd vccd wire1571/X sky130_fd_sc_hd__buf_6
Xwire1582 wire1583/X vssd vssd vccd vccd _336_/B sky130_fd_sc_hd__buf_6
Xwire1593 wire1594/X vssd vssd vccd vccd wire1593/X sky130_fd_sc_hd__buf_6
XFILLER_17_3409 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_3723 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_557 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output692_A _059_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1219_A _463_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_3133 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_2192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__C _483_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1021 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] load_slew1458/X vssd vssd vccd vccd _129_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_11_1606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1588_A wire1589/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1065 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3301 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1755_A wire1755/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1022 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3389 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1976 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] _276_/X vssd vssd vccd vccd _096_/A
+ sky130_fd_sc_hd__nand2_8
XFILLER_2_1818 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3932 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_365 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_3976 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__393__C _393_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2521 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_273 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1252 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_295 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2303 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2069_A wire2069/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_3660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4408 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input221_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2236_A wire2236/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input319_A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_3133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4012 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4154 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__584__B _584_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4029 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_2627 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_116_ _116_/A vssd vssd vccd vccd _116_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_51_1997 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__105__A _105_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_4261 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_047_ _047_/A vssd vssd vccd vccd _047_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_10_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3571 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_461 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output538_A wire1240/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1071_A wire1072/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_3529 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1169_A _536_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2817 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_2997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__478__C _478_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output705_A _071_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire2080 wire2081/X vssd vssd vccd vccd _591_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2091 wire2091/A vssd vssd vccd vccd wire2091/X sky130_fd_sc_hd__buf_6
XFILLER_21_3192 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_wire1336_A _358_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1390 _340_/X vssd vssd vccd vccd wire1390/X sky130_fd_sc_hd__buf_6
XFILLER_19_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__494__B _494_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_B _282_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_4265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1503_A wire1504/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_2527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_516 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4129 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1706 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2841 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1127 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2885 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2148 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__015__A _015_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2801 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_A mprj_dat_i_user[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_2906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_866 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_888 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_685 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_195 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_2941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1959 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3973 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input171_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1970 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input269_A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2186_A wire2187/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3996 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__579__B _579_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_3755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[19\]_A mprj_dat_i_user[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input436_A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3849 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput310 la_oenb_mprj[2] vssd vssd vccd vccd _499_/A sky130_fd_sc_hd__buf_4
Xinput321 la_oenb_mprj[3] vssd vssd vccd vccd _500_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3799 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input32_A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput332 la_oenb_mprj[4] vssd vssd vccd vccd _501_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput343 la_oenb_mprj[5] vssd vssd vccd vccd _502_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput354 la_oenb_mprj[6] vssd vssd vccd vccd _503_/A sky130_fd_sc_hd__buf_4
Xinput365 la_oenb_mprj[7] vssd vssd vccd vccd _504_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_48_457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1621 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput376 la_oenb_mprj[8] vssd vssd vccd vccd _505_/A sky130_fd_sc_hd__buf_6
XFILLER_36_608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput387 la_oenb_mprj[9] vssd vssd vccd vccd _506_/A sky130_fd_sc_hd__buf_4
Xinput398 mprj_adr_o_core[19] vssd vssd vccd vccd wire1647/A sky130_fd_sc_hd__buf_6
XANTENNA__595__A _595_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1665 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_596_ _596_/A _596_/B vssd vssd vccd vccd _596_/X sky130_fd_sc_hd__and2_4
XFILLER_16_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_93 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_398 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output488_A wire1206/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_4367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_3633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output655_A _025_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_3 la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_3081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput806 _560_/X vssd vssd vccd vccd la_oenb_core[63] sky130_fd_sc_hd__buf_8
XFILLER_42_4501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput817 _570_/X vssd vssd vccd vccd la_oenb_core[73] sky130_fd_sc_hd__buf_8
XFILLER_6_65 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput828 _580_/X vssd vssd vccd vccd la_oenb_core[83] sky130_fd_sc_hd__buf_8
XFILLER_29_2932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1286_A _377_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput839 _590_/X vssd vssd vccd vccd la_oenb_core[93] sky130_fd_sc_hd__buf_8
XFILLER_42_4545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output822_A _575_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4185 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2807 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_2277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3473 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__B _489_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1453_A wire1454/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3254 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1620_A wire1621/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3637 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_162 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3946 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_52_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4423 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1211 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3204 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1255 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4033 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2328 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_3917 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1020 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4536 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_3448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1373 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ _578_/A _450_/B _450_/C vssd vssd vccd vccd _450_/X sky130_fd_sc_hd__and3b_4
XTAP_2747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_674 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4173 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_381_ _509_/A _381_/B _381_/C vssd vssd vccd vccd _381_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_324 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3581 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3434 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2101_A wire2102/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_4209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input386_A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_3781 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1199 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2829 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_4231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3107 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1527 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4275 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3613 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_2417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3563 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2057 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_250 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2934 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput140 la_iena_mprj[107] vssd vssd vccd vccd _270_/B sky130_fd_sc_hd__clkbuf_4
Xinput151 la_iena_mprj[117] vssd vssd vccd vccd _280_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xinput162 la_iena_mprj[127] vssd vssd vccd vccd _290_/B sky130_fd_sc_hd__buf_4
XFILLER_37_928 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput173 la_iena_mprj[21] vssd vssd vccd vccd _184_/B sky130_fd_sc_hd__buf_4
XTAP_4650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput184 la_iena_mprj[31] vssd vssd vccd vccd _194_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_4661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 la_iena_mprj[41] vssd vssd vccd vccd _204_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_4683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3312 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2691 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_641 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1034_A wire1035/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2611 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_3247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3367 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2081 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_579_ _579_/A _579_/B vssd vssd vccd vccd _579_/X sky130_fd_sc_hd__and2_4
XFILLER_53_2546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4257 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1201_A _496_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_output772_A _529_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__491__C _491_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_53_1889 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4236 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4006 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1570_A wire1571/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_3917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput603 _093_/Y vssd vssd vccd vccd la_data_in_mprj[110] sky130_fd_sc_hd__buf_8
XFILLER_9_3524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput614 _103_/Y vssd vssd vccd vccd la_data_in_mprj[120] sky130_fd_sc_hd__buf_8
XANTENNA_wire1668_A wire1669/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_4039 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput625 _162_/Y vssd vssd vccd vccd la_data_in_mprj[15] sky130_fd_sc_hd__buf_8
XFILLER_47_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput636 _008_/Y vssd vssd vccd vccd la_data_in_mprj[25] sky130_fd_sc_hd__buf_8
XFILLER_29_3485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput647 _018_/Y vssd vssd vccd vccd la_data_in_mprj[35] sky130_fd_sc_hd__buf_8
XFILLER_42_4353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xoutput658 _028_/Y vssd vssd vccd vccd la_data_in_mprj[45] sky130_fd_sc_hd__buf_8
XFILLER_45_2041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput669 _038_/Y vssd vssd vccd vccd la_data_in_mprj[55] sky130_fd_sc_hd__buf_8
XFILLER_28_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_2995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_3445 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4580 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4308 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4488 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2045 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2067 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_165 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1339 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4404 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__203__A _203_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3933 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4448 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3883 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3977 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1901 wire1902/X vssd vssd vccd vccd _264_/A sky130_fd_sc_hd__buf_6
XFILLER_41_3173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2399 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1912 wire1912/A vssd vssd vccd vccd _258_/A sky130_fd_sc_hd__buf_6
Xwire1923 wire1923/A vssd vssd vccd vccd _243_/A sky130_fd_sc_hd__buf_4
Xwire1934 wire1934/A vssd vssd vccd vccd _333_/A sky130_fd_sc_hd__buf_6
Xwire1945 wire1945/A vssd vssd vccd vccd _192_/A sky130_fd_sc_hd__buf_6
XTAP_3201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input134_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2051_A wire2051/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1956 wire1957/X vssd vssd vccd vccd _183_/A sky130_fd_sc_hd__buf_6
XTAP_3212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire2149_A wire2150/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xwire1967 wire1967/A vssd vssd vccd vccd _177_/A sky130_fd_sc_hd__buf_6
XFILLER_46_725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_3223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1978 wire1978/A vssd vssd vccd vccd wire1978/X sky130_fd_sc_hd__buf_6
XTAP_3234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1989 wire1989/A vssd vssd vccd vccd wire1989/X sky130_fd_sc_hd__buf_6
XTAP_3245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _340_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _284_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_502_ _502_/A _502_/B vssd vssd vccd vccd _502_/X sky130_fd_sc_hd__and2_4
XFILLER_27_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2519 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input301_A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_223 _563_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_3289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 _342_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_433_ _561_/A _433_/B _433_/C vssd vssd vccd vccd _433_/X sky130_fd_sc_hd__and3b_4
XTAP_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2221 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_289 wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_2599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_1865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__592__B _592_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_1876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_1887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_364_ _364_/A _364_/B vssd vssd vccd vccd _364_/X sky130_fd_sc_hd__and2_2
XFILLER_35_2265 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_2107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_125 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_187 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_295_ _295_/A_N _295_/B vssd vssd vccd vccd _295_/X sky130_fd_sc_hd__and2b_4
XFILLER_9_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xrebuffer6 wire1460/X vssd vssd vccd vccd rebuffer6/X sky130_fd_sc_hd__bufbuf_8
XFILLER_6_843 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_4359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3051 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2659 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1407 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2361 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1969 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4133 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_4019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_output520_A wire1257/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_3224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_2269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2742 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1151_A _555_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1249_A _413_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_2545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__486__C _486_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__396__A_N _524_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_4491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3721 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_961 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3120 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] _195_/X vssd vssd vccd vccd _015_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_18_3164 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_51_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2441 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3186 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1317 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_474 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_4087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_3353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2630 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_669 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1785_A wire1785/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2641 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_670 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_4022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4044 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1952_A wire1952/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4088 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1413 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__023__A _023_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput466 wire1213/X vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__buf_8
Xoutput477 _481_/X vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__buf_8
XFILLER_47_1457 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xoutput488 wire1206/X vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__buf_8
Xoutput499 wire1277/X vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__buf_8
XFILLER_9_2675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xwire1208 _476_/X vssd vssd vccd vccd wire1208/X sky130_fd_sc_hd__buf_6
XFILLER_41_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1219 _463_/X vssd vssd vccd vccd wire1219/X sky130_fd_sc_hd__buf_6
XFILLER_9_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4492 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1849 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_2241 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3780 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__396__C _396_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_4506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_791 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_3275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_953 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2405 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4116 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2585 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_2449 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4337 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_629 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2703 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_080_ _080_/A vssd vssd vccd vccd _080_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_2913 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2099_A wire2100/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2501 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4212 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input251_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_3730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input349_A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2266_A wire2267/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2545 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4256 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2589 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1720 _400_/A_N vssd vssd vccd vccd _528_/A sky130_fd_sc_hd__buf_6
Xwire1731 wire1731/A vssd vssd vccd vccd _613_/A sky130_fd_sc_hd__buf_6
XANTENNA__587__B _587_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_3577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1742 input19/X vssd vssd vccd vccd _482_/C sky130_fd_sc_hd__buf_6
XFILLER_21_3588 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1753 wire1753/A vssd vssd vccd vccd _449_/C sky130_fd_sc_hd__buf_6
XFILLER_24_1265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1107 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1764 wire1765/X vssd vssd vccd vccd _388_/B sky130_fd_sc_hd__buf_6
XFILLER_46_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1775 wire1775/A vssd vssd vccd vccd wire1775/X sky130_fd_sc_hd__buf_6
XTAP_3031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire1786 wire1787/X vssd vssd vccd vccd _378_/B sky130_fd_sc_hd__buf_6
XFILLER_37_3017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1797 wire1797/A vssd vssd vccd vccd wire1797/X sky130_fd_sc_hd__buf_6
XTAP_3053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3304 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_2374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3949 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_4341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_416_ _416_/A_N _416_/B _416_/C vssd vssd vccd vccd _416_/X sky130_fd_sc_hd__and3b_4
XTAP_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_2505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_2636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_2073 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__108__A _108_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_2549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_347_ _347_/A _347_/B vssd vssd vccd vccd _347_/X sky130_fd_sc_hd__and2_4
X_278_ _278_/A _278_/B vssd vssd vccd vccd _278_/X sky130_fd_sc_hd__and2_4
XFILLER_31_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output470_A wire1209/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_2371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3960 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output568_A wire1287/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_3709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4123 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1199_A _498_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output735_A _611_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1733 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1121 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1777 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1366_A _348_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_2607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_output902_A wire974/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_3262 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__497__B _497_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_3137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2331 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3415 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_4572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_901 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2725 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_783 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4436 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1147 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_3773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_2769 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3161 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__411__A_N _539_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_49_2209 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1309 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2507 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3151 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_3555 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4532 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_838 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_3820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2865 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1287 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_2483 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1005 _137_/Y vssd vssd vccd vccd wire1005/X sky130_fd_sc_hd__buf_6
XFILLER_40_2729 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1016 wire1017/X vssd vssd vccd vccd wire1016/X sky130_fd_sc_hd__buf_6
XFILLER_38_4005 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1027 wire1028/X vssd vssd vccd vccd wire1027/X sky130_fd_sc_hd__buf_6
Xwire1038 wire1039/X vssd vssd vccd vccd wire1038/X sky130_fd_sc_hd__buf_6
XFILLER_0_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire1049 wire1050/X vssd vssd vccd vccd wire1049/X sky130_fd_sc_hd__buf_6
XFILLER_0_4383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1679 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_2603 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_503 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1381 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_249 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_709 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1957 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3668 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4060 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1345 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2014_A wire2015/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_2825 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2213 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4101 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2393 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_201_ _201_/A _201_/B vssd vssd vccd vccd _201_/X sky130_fd_sc_hd__and2_2
XFILLER_11_433 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input299_A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_132_ _132_/A vssd vssd vccd vccd _132_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_32_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_477 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1545 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_2680 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_063_ _063_/A vssd vssd vccd vccd _063_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_2555 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_4537 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input62_A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2599 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4487 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1917 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3869 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__598__A _598_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_809 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2240 wire2241/X vssd vssd vccd vccd _467_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_4086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_4169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2251 wire2251/A vssd vssd vccd vccd _458_/B sky130_fd_sc_hd__buf_6
Xwire2262 wire2263/X vssd vssd vccd vccd _454_/B sky130_fd_sc_hd__buf_6
XFILLER_40_3997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xwire2273 wire2274/X vssd vssd vccd vccd _450_/B sky130_fd_sc_hd__buf_6
XFILLER_21_3374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire2284 wire2284/A vssd vssd vccd vccd _442_/B sky130_fd_sc_hd__buf_6
XFILLER_1_2712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1550 wire1551/X vssd vssd vccd vccd wire1550/X sky130_fd_sc_hd__buf_6
XFILLER_21_3385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2295 wire2295/A vssd vssd vccd vccd _433_/B sky130_fd_sc_hd__buf_6
XFILLER_5_2892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire1561 wire1562/X vssd vssd vccd vccd wire1561/X sky130_fd_sc_hd__buf_6
XFILLER_47_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2745 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xwire1572 wire1573/X vssd vssd vccd vccd _309_/B sky130_fd_sc_hd__buf_6
Xwire1583 wire1584/X vssd vssd vccd vccd wire1583/X sky130_fd_sc_hd__buf_6
XFILLER_1_2756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xwire1594 wire1595/X vssd vssd vccd vccd wire1594/X sky130_fd_sc_hd__buf_6
XFILLER_21_2695 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3893 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1401 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3123 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_569 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_3779 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire1114_A wire1115/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__434__A_N _562_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_4171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_2909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2319 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output852_A wire1410/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1689 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1077 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4003 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1541 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1650_A wire1651/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1748_A wire1748/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1034 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__301__A _301_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2595 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4325 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1173 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] wire1462/X vssd vssd vccd vccd
+ _089_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_2266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2967 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_3944 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_4200 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4380 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2533 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2577 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2017 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1286 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_4053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2315 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2409 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4340 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2359 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2673 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2291 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__211__A _211_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_3891 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2166 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_820 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1246 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_3145 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input214_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_85 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2131_A wire2131/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4122 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__457__A_N _585_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire2229_A wire2229/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_51_4024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3009 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3189 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_867 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_4166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_517 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3919 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1765 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3307 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3329 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_3498 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1921 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1039 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_4505 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2677 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_2639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2087 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1353 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4549 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_115_ _115_/A vssd vssd vccd vccd _115_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_45_3105 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2352 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1397 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3285 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_046_ _046_/A vssd vssd vccd vccd _046_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_3600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_3149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1662 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_49_1861 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_473 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_4451 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3761 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1229 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1064_A wire1065/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_3160 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2070 wire2071/X vssd vssd vccd vccd _297_/A sky130_fd_sc_hd__buf_6
Xwire2081 wire2081/A vssd vssd vccd vccd wire2081/X sky130_fd_sc_hd__buf_6
XFILLER_36_4509 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xwire2092 wire2093/X vssd vssd vccd vccd _583_/B sky130_fd_sc_hd__buf_6
XFILLER_43_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1380 wire1381/X vssd vssd vccd vccd wire1380/X sky130_fd_sc_hd__buf_6
XFILLER_35_812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xwire1391 wire1392/X vssd vssd vccd vccd wire1391/X sky130_fd_sc_hd__buf_6
XANTENNA_wire1231_A _426_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_2492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2575 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1329_A wire1330/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_52_3109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_867 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__494__C _494_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_377 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_837 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4520 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2853 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4564 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_2897 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1865_A wire1866/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_50_1497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1448 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_4237 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2813 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3165 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_3176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2993 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_B split5/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__031__A _031_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2857 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_3608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1605 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_149 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_2907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_4199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_3465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_2918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_4333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3329 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_193 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3610 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_52_3621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_1290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3752 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1905 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3638 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1326 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3985 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__206__A _206_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_727 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_3425 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_49_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3469 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_53 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1157 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2081_A wire2081/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input164_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2217 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2179_A wire2180/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1909 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[19\]_B load_slew1458/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput300 la_oenb_mprj[20] vssd vssd vccd vccd _517_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput311 la_oenb_mprj[30] vssd vssd vccd vccd wire1721/A sky130_fd_sc_hd__buf_6
Xinput322 la_oenb_mprj[40] vssd vssd vccd vccd _409_/A_N sky130_fd_sc_hd__buf_6
XFILLER_40_2323 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput333 la_oenb_mprj[50] vssd vssd vccd vccd _547_/A sky130_fd_sc_hd__buf_4
XANTENNA_input331_A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput344 la_oenb_mprj[60] vssd vssd vccd vccd _557_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input429_A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput355 la_oenb_mprj[70] vssd vssd vccd vccd wire1702/A sky130_fd_sc_hd__buf_6
XFILLER_2_4297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput366 la_oenb_mprj[80] vssd vssd vccd vccd wire1692/A sky130_fd_sc_hd__buf_6
XANTENNA_input25_A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput377 la_oenb_mprj[90] vssd vssd vccd vccd _587_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1633 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput388 mprj_adr_o_core[0] vssd vssd vccd vccd wire1679/A sky130_fd_sc_hd__buf_6
Xinput399 mprj_adr_o_core[1] vssd vssd vccd vccd wire1644/A sky130_fd_sc_hd__buf_6
XFILLER_21_1032 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_4228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__595__B _595_/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1677 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1065 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_595_ _595_/A _595_/B vssd vssd vccd vccd _595_/X sky130_fd_sc_hd__and2_4
XFILLER_31_4417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_3863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_2739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_2149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1426 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_2463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_2583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_881 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4313 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA__116__A _116_/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_2458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1172 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_4 la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput807 _561_/X vssd vssd vccd vccd la_oenb_core[64] sky130_fd_sc_hd__buf_8
XFILLER_10_2171 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput818 _571_/X vssd vssd vccd vccd la_oenb_core[74] sky130_fd_sc_hd__buf_8
XFILLER_49_3093 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output550_A _432_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput829 _581_/X vssd vssd vccd vccd la_oenb_core[84] sky130_fd_sc_hd__buf_8
XFILLER_6_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_029_ _029_/A vssd vssd vccd vccd _029_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_2955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1181_A _516_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_wire1279_A _384_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__489__C _489_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2109 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output815_A _568_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XTAP_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1446_A wire1447/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1037 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] _225_/X vssd vssd vccd vccd _045_/A
+ sky130_fd_sc_hd__nand2_4
XFILLER_23_2587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_wire1613_A wire1614/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_3605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2350 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4041 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3649 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2303 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_2314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4085 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_174 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_50_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1982_A wire1983/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2661 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_369 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_50_1261 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1835 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_4479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_3745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4001 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3609 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1267 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_3789 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4181 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2421 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3177 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4045 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2465 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__399__C _399_/C vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_4089 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_4106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2687 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_3405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1341 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_4548 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1385 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3836 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_2726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3273 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_2737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3137 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_461 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_686 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_380_ _508_/A _380_/B _380_/C vssd vssd vccd vccd _380_/X sky130_fd_sc_hd__and3b_4
XFILLER_13_3413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_4158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4450 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1735 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_3446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_177 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_892 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_391 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_3793 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input281_A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1481 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3192 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2296_A wire2296/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_input379_A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_3277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_3761 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_3531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_4287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3575 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1875 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_3417 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4061 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_23_1105 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput130 la_data_out_mprj[99] vssd vssd vccd vccd _468_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2863 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput141 la_iena_mprj[108] vssd vssd vccd vccd _271_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1357 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_233 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput152 la_iena_mprj[118] vssd vssd vccd vccd _281_/B sky130_fd_sc_hd__clkbuf_4
Xinput163 la_iena_mprj[12] vssd vssd vccd vccd _175_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 la_iena_mprj[22] vssd vssd vccd vccd _185_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1441 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xinput185 la_iena_mprj[32] vssd vssd vccd vccd _195_/B sky130_fd_sc_hd__clkbuf_4
XTAP_4662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_277 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xinput196 la_iena_mprj[42] vssd vssd vccd vccd _205_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_36_417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_4673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1485 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_951 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_3324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_3972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XTAP_3983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_3969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_141 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_601 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4225 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
X_578_ _578_/A _578_/B vssd vssd vccd vccd _578_/X sky130_fd_sc_hd__and2_4
XANTENNA_wire1027_A wire1028/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_53_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output598_A _089_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_2667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4269 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_2801 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_53_1846 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_2981 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XPHY_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output765_A wire1174/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_4143 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_51_1581 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1396_A _337_/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_4248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4018 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output932_A wire1311/X vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput604 _094_/Y vssd vssd vccd vccd la_data_in_mprj[111] sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3453 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput615 _104_/Y vssd vssd vccd vccd la_data_in_mprj[121] sky130_fd_sc_hd__buf_8
XFILLER_44_3929 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4321 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput626 _163_/Y vssd vssd vccd vccd la_data_in_mprj[16] sky130_fd_sc_hd__buf_8
XFILLER_47_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xoutput637 _009_/Y vssd vssd vccd vccd la_data_in_mprj[26] sky130_fd_sc_hd__buf_8
Xoutput648 _019_/Y vssd vssd vccd vccd la_data_in_mprj[36] sky130_fd_sc_hd__buf_8
XANTENNA_wire1563_A wire1563/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_3497 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
Xoutput659 _029_/Y vssd vssd vccd vccd la_data_in_mprj[46] sky130_fd_sc_hd__buf_8
XFILLER_42_4365 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2053 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1049 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2941 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2097 vssd vssd vccd vccd sky130_ef_sc_hd__decap_12
.ends

