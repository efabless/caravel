VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravan_core
  CLASS BLOCK ;
  FOREIGN caravan_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 3165.000 BY 4767.000 ;
END caravan_core
END LIBRARY