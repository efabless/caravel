magic
tech sky130A
magscale 1 2
timestamp 1686151263
<< checkpaint >>
rect 674245 108867 676990 111443
rect 674143 103403 677009 105940
rect 674244 103347 676989 103403
<< metal1 >>
rect 675778 117266 675830 117272
rect 675778 117208 675830 117214
rect 675682 113371 675734 115709
rect 675586 112665 675638 112671
rect 675586 112487 675638 112493
rect 675490 109630 675542 109636
rect 675490 109452 675542 109458
rect 675492 101631 675540 109452
rect 675588 108347 675636 112487
rect 675682 109050 675734 113199
rect 675586 108341 675638 108347
rect 675586 108163 675638 108169
rect 675490 101625 675542 101631
rect 675490 101567 675542 101573
rect 675492 100265 675540 101567
rect 675588 100462 675636 108163
rect 675586 100456 675638 100462
rect 675586 100278 675638 100284
rect 675588 100265 675636 100278
rect 675682 99896 675734 108866
rect 675780 102183 675828 117208
rect 675778 102177 675830 102183
rect 675778 102119 675830 102125
rect 675780 102106 675828 102119
<< via1 >>
rect 675778 117214 675830 117266
rect 675682 113199 675734 113371
rect 675586 112493 675638 112665
rect 675490 109458 675542 109630
rect 675682 108866 675734 109050
rect 675586 108169 675638 108341
rect 675490 101573 675542 101625
rect 675586 100284 675638 100456
rect 675778 102125 675830 102177
<< metal2 >>
rect 675772 117214 675778 117266
rect 675830 117264 675836 117266
rect 676699 117264 676708 117270
rect 675830 117216 676708 117264
rect 675830 117214 675836 117216
rect 676699 117210 676708 117216
rect 676768 117210 676777 117270
rect 675495 115647 675505 115703
rect 675730 115647 675740 115703
rect 675495 115095 675505 115151
rect 675730 115095 675740 115151
rect 675490 114451 675506 114507
rect 675731 114451 675747 114507
rect 675496 113807 675506 113863
rect 675731 113807 675741 113863
rect 675676 113311 675682 113371
rect 675407 113255 675682 113311
rect 675676 113199 675682 113255
rect 675734 113311 675740 113371
rect 675734 113255 675887 113311
rect 675734 113199 675740 113255
rect 675407 112665 675887 112667
rect 675407 112611 675586 112665
rect 675580 112493 675586 112611
rect 675638 112611 675887 112665
rect 675638 112493 675644 112611
rect 675496 111967 675506 112023
rect 675731 111967 675741 112023
rect 675495 111415 675505 111471
rect 675730 111415 675740 111471
rect 675495 110771 675505 110827
rect 675730 110771 675740 110827
rect 675407 109630 675887 109631
rect 675407 109575 675490 109630
rect 675484 109458 675490 109575
rect 675542 109575 675887 109630
rect 675542 109458 675548 109575
rect 675676 108866 675682 109050
rect 675734 108866 675740 109050
rect 675407 108341 675887 108343
rect 675407 108287 675586 108341
rect 675580 108169 675586 108287
rect 675638 108287 675887 108341
rect 675638 108169 675644 108287
rect 675496 107643 675505 107699
rect 675730 107643 675739 107699
rect 675496 107091 675506 107147
rect 675731 107091 675741 107147
rect 675496 106447 675506 106503
rect 675731 106447 675741 106503
rect 675495 105803 675505 105859
rect 675730 105803 675740 105859
rect 675494 105251 675504 105307
rect 675729 105251 675739 105307
rect 675496 103411 675506 103467
rect 675731 103411 675741 103467
rect 675495 102767 675505 102823
rect 675730 102767 675740 102823
rect 675762 102177 675840 102179
rect 675762 102125 675778 102177
rect 675830 102125 675840 102177
rect 675762 102123 675840 102125
rect 675407 101625 675887 101627
rect 675407 101573 675490 101625
rect 675542 101573 675887 101625
rect 675407 101571 675887 101573
rect 675495 100927 675505 100983
rect 675730 100927 675740 100983
rect 675580 100339 675586 100456
rect 675407 100284 675586 100339
rect 675638 100339 675644 100456
rect 675638 100284 675887 100339
rect 675407 100283 675887 100284
<< via2 >>
rect 676708 117210 676768 117270
rect 675505 115647 675730 115703
rect 675505 115095 675730 115151
rect 675506 114451 675731 114507
rect 675506 113807 675731 113863
rect 675506 111967 675731 112023
rect 675505 111415 675730 111471
rect 675505 110771 675730 110827
rect 675505 110127 675730 110183
rect 675505 107643 675730 107699
rect 675506 107091 675731 107147
rect 675506 106447 675731 106503
rect 675505 105803 675730 105859
rect 675504 105251 675729 105307
rect 675504 104607 675729 104663
rect 675506 103411 675731 103467
rect 675505 102767 675730 102823
rect 675505 100927 675730 100983
<< metal3 >>
rect 676708 117275 676768 117452
rect 676703 117270 676773 117275
rect 676703 117210 676708 117270
rect 676768 117210 676773 117270
rect 676703 117205 676773 117210
rect 675407 115703 675887 115710
rect 675407 115647 675505 115703
rect 675730 115647 675887 115703
rect 675407 115640 675887 115647
rect 675407 115151 675887 115158
rect 675407 115095 675505 115151
rect 675730 115095 675887 115151
rect 675407 115088 675887 115095
rect 675407 114507 675887 114514
rect 675407 114451 675506 114507
rect 675731 114451 675887 114507
rect 675407 114444 675887 114451
rect 675407 113863 675887 113870
rect 675407 113807 675506 113863
rect 675731 113807 675887 113863
rect 675407 113800 675887 113807
rect 675407 112023 675887 112030
rect 675407 111967 675506 112023
rect 675731 111967 675887 112023
rect 675407 111960 675887 111967
rect 675407 111471 675887 111478
rect 675407 111415 675505 111471
rect 675730 111415 675887 111471
rect 675407 111408 675887 111415
rect 675407 110827 675887 110834
rect 675407 110771 675505 110827
rect 675730 110771 675887 110827
rect 675407 110764 675887 110771
rect 675407 110183 675887 110190
rect 675407 110127 675505 110183
rect 675730 110127 675887 110183
rect 675407 110120 675887 110127
rect 675407 107699 675887 107706
rect 675407 107643 675505 107699
rect 675730 107643 675887 107699
rect 675407 107636 675887 107643
rect 675407 107147 675887 107154
rect 675407 107091 675506 107147
rect 675731 107091 675887 107147
rect 675407 107084 675887 107091
rect 675407 106503 675887 106510
rect 675407 106447 675506 106503
rect 675731 106447 675887 106503
rect 675407 106440 675887 106447
rect 675407 105859 675887 105866
rect 675407 105803 675505 105859
rect 675730 105803 675887 105859
rect 675407 105796 675887 105803
rect 675406 105307 675886 105314
rect 675406 105251 675504 105307
rect 675729 105251 675886 105307
rect 675406 105244 675886 105251
rect 675407 104663 675887 104670
rect 675407 104607 675504 104663
rect 675729 104607 675887 104663
rect 675407 104600 675887 104607
rect 675407 103467 675887 103474
rect 675407 103411 675506 103467
rect 675731 103411 675887 103467
rect 675407 103404 675887 103411
rect 675407 102823 675887 102830
rect 675407 102767 675505 102823
rect 675730 102767 675887 102823
rect 675407 102760 675887 102767
rect 675407 100983 675887 100990
rect 675407 100927 675505 100983
rect 675730 100927 675887 100983
rect 675407 100920 675887 100927
<< properties >>
string flatten true
<< end >>
