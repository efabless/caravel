* NGSPICE file created from housekeeping_alt.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_2 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_4 abstract view
.subckt sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt housekeeping_alt VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0]
+ irq[1] irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XANTENNA__3691__A2 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5968__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6914_ _6926_/CLK _6914_/D fanout566/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_hold2978_A _7183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6845_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6845_/X sky130_fd_sc_hd__and2_1
XFILLER_0_193_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6776_ _6751_/S _6776_/A2 _6774_/Y _6775_/X VGND VGND VPWR VPWR _6776_/X sky130_fd_sc_hd__a22o_1
X_3988_ _3988_/A _3988_/B _3988_/C _3988_/D VGND VGND VPWR VPWR _3995_/C sky130_fd_sc_hd__nor4_1
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5727_ _5727_/A0 hold84/X _5730_/S VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3746__A3 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6145__A1 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5658_ _5955_/A1 _5658_/A1 _5658_/S VGND VGND VPWR VPWR _5658_/X sky130_fd_sc_hd__mux2_1
X_4609_ _4887_/D _4747_/B _4887_/B _4879_/C _4805_/B VGND VGND VPWR VPWR _4909_/A
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__6696__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5589_ _5589_/A0 _5805_/A1 _5589_/S VGND VGND VPWR VPWR _5589_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold340 hold340/A VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7328_ _7359_/CLK _7328_/D fanout576/X VGND VGND VPWR VPWR _7328_/Q sky130_fd_sc_hd__dfstp_4
Xhold351 _5933_/X VGND VGND VPWR VPWR _7522_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold362 hold362/A VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold373 hold373/A VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4829__B _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold384 hold384/A VGND VGND VPWR VPWR hold384/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__A2 _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7259_ _7510_/CLK _7259_/D fanout603/X VGND VGND VPWR VPWR _7259_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4459__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5656__A0 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5120__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4845__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 hold2891/X VGND VGND VPWR VPWR _7260_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1051 hold2748/X VGND VGND VPWR VPWR hold2749/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1062 hold2798/X VGND VGND VPWR VPWR hold2799/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input127_A wb_adr_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1073 _4492_/X VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5959__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1084 hold2917/X VGND VGND VPWR VPWR hold2918/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _4377_/X VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6620__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A3 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4580__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_38_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5187__A2 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input92_A spimemio_flash_io3_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4395__A0 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6687__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5895__A0 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6439__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5647__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4905__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6611__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4960_ _4960_/A _4960_/B VGND VGND VPWR VPWR _5252_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_188_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3911_ _6912_/Q _5612_/B _5947_/A _3657_/X _6958_/Q VGND VGND VPWR VPWR _3911_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4891_ _5222_/B _5222_/C _4937_/C _4891_/D VGND VGND VPWR VPWR _4891_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3976__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6630_ _7574_/Q _6424_/X _6628_/X _6629_/X VGND VGND VPWR VPWR _6630_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5178__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3842_ _7505_/Q _5983_/A _5938_/C _3841_/X VGND VGND VPWR VPWR _3842_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5032__D1 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4921__C _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4386__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6561_ _7371_/Q _6459_/B _6429_/X _6468_/X _7411_/Q VGND VGND VPWR VPWR _6561_/X
+ sky130_fd_sc_hd__a32o_1
X_3773_ _7490_/Q _3569_/X _3765_/X _3772_/X VGND VGND VPWR VPWR _3773_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3728__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5512_ _5512_/A _5575_/A _5548_/A _5512_/D VGND VGND VPWR VPWR _5512_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3537__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6492_ _7312_/Q _6419_/D _6452_/X _7344_/Q VGND VGND VPWR VPWR _6492_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6127__B2 _7336_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6678__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5443_ _4601_/Y _4956_/B _4659_/Y VGND VGND VPWR VPWR _5541_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5350__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5374_ _4703_/Y _4846_/Y _4428_/B _5373_/X VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__o211a_1
X_7113_ _7196_/CLK _7113_/D fanout589/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3553__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4325_ _5950_/A1 _4325_/A1 _4327_/S VGND VGND VPWR VPWR _4325_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5638__A0 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7044_ _7201_/CLK _7044_/D _6839_/A VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_4
X_4256_ _4256_/A0 _4256_/A1 _4258_/S VGND VGND VPWR VPWR _4256_/X sky130_fd_sc_hd__mux2_1
X_4187_ _4187_/A0 _7640_/Q _4429_/B VGND VGND VPWR VPWR _4187_/X sky130_fd_sc_hd__mux2_8
XANTENNA_fanout377_A _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6063__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6602__A2 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3967__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6828_ hold45/A _7107_/Q _6798_/C VGND VGND VPWR VPWR _6828_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6366__A1 _6965_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4831__C _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3719__A3 _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6759_ _7015_/Q _4105_/B _6459_/B _6467_/X _7156_/Q VGND VGND VPWR VPWR _6759_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6669__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6120__A _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold170 hold170/A VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold181 hold181/A VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold192 hold192/A VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4301__A0 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4575__A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4852__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A3 _3496_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3591__A1 input59/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3654__A _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3894__A2 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4110_ _7110_/Q _4084_/X _4425_/B VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__a21o_1
X_5090_ _4774_/Y _4960_/A _5089_/Y _5088_/Y VGND VGND VPWR VPWR _5090_/Y sky130_fd_sc_hd__o211ai_1
Xhold1809 _7525_/Q VGND VGND VPWR VPWR hold116/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6293__B1 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4041_ _4041_/A1 _4040_/D _4040_/A _4044_/A1 VGND VGND VPWR VPWR _4042_/B sky130_fd_sc_hd__a22oi_1
XANTENNA__4485__A _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5992_ hold36/X hold22/X _5992_/C _5992_/D VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__and4_4
XFILLER_0_189_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4943_ _5248_/B _4943_/B VGND VGND VPWR VPWR _4944_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3949__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4932__B _4932_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7662_ _7662_/A VGND VGND VPWR VPWR _7662_/X sky130_fd_sc_hd__clkbuf_2
X_4874_ _4984_/B _4984_/A _4668_/C _5100_/A VGND VGND VPWR VPWR _5203_/B sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_145_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6613_ _7317_/Q _6419_/D _6424_/X _7573_/Q _6612_/X VGND VGND VPWR VPWR _6613_/X
+ sky130_fd_sc_hd__a221o_1
X_3825_ _7174_/Q _4509_/A _5623_/B _5581_/A _7211_/Q VGND VGND VPWR VPWR _3825_/X
+ sky130_fd_sc_hd__a32o_1
X_7593_ _7593_/CLK _7593_/D fanout567/X VGND VGND VPWR VPWR _7593_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_15_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6544_ _6544_/A _6544_/B _6544_/C _6544_/D VGND VGND VPWR VPWR _6545_/C sky130_fd_sc_hd__nor4_2
X_3756_ _7554_/Q _3508_/X _4422_/S input46/X _3755_/X VGND VGND VPWR VPWR _3759_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_172_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_6475_ _7448_/Q _6467_/A _6574_/C _6408_/B _7376_/Q VGND VGND VPWR VPWR _6475_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5859__A0 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3687_ _7176_/Q _5875_/A _5623_/B _3537_/X _7427_/Q VGND VGND VPWR VPWR _3687_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3564__A _3564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5426_ _5158_/A _5342_/B _5038_/B _5183_/A VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__o211a_1
Xoutput220 _7658_/X VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
XANTENNA__5323__A2 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput231 _7668_/X VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput242 _7652_/X VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
Xoutput253 _4132_/A VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
Xoutput264 _7228_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
X_5357_ _4947_/C _5213_/C _5346_/X _5102_/B _5357_/B2 VGND VGND VPWR VPWR _5357_/X
+ sky130_fd_sc_hd__a32o_1
Xoutput275 _6918_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
Xoutput286 _6928_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
XANTENNA__3885__A2 _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput297 _7246_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4308_ _4308_/A0 _5754_/A1 _4308_/S VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__mux2_1
X_5288_ _4847_/X _5061_/X _5286_/X _5123_/X VGND VGND VPWR VPWR _5288_/Y sky130_fd_sc_hd__o31ai_2
X_7027_ _7196_/CLK _7027_/D fanout589/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfrtp_4
X_4239_ _4239_/A0 _4238_/X _4249_/S VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_179_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5938__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1943_A _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire347 _6647_/Y VGND VGND VPWR VPWR wire347/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3157_A _7243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input55_A mgmt_gpio_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3876__A2 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5078__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6275__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3628__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout480 _5735_/A1 VGND VGND VPWR VPWR _5951_/A1 sky130_fd_sc_hd__buf_12
XANTENNA__4736__C _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout491 _5940_/A1 VGND VGND VPWR VPWR _5583_/A0 sky130_fd_sc_hd__clkbuf_16
XANTENNA__6290__A3 _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6009__B _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6027__B1 _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4455__D hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5848__B hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5250__A1 _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3649__A _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4244__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_732 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3800__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3610_ _7356_/Q _5803_/A _4212_/A _3494_/X _7476_/Q VGND VGND VPWR VPWR _3610_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_71_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4590_ _5071_/A _4825_/A VGND VGND VPWR VPWR _4591_/B sky130_fd_sc_hd__and2b_4
XANTENNA_max_cap557_A _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6750__B2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3541_ _5938_/B _4491_/A VGND VGND VPWR VPWR _3541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold906 _4379_/X VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold917 hold917/A VGND VGND VPWR VPWR hold917/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold928 _4507_/X VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6260_ _6649_/S _6260_/A2 _6258_/X _6259_/X _6777_/S VGND VGND VPWR VPWR _6260_/X
+ sky130_fd_sc_hd__a221o_1
Xhold939 hold939/A VGND VGND VPWR VPWR hold939/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4108__A3 _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3472_ _4551_/A _3507_/A _3576_/C VGND VGND VPWR VPWR _3472_/X sky130_fd_sc_hd__and3_2
X_5211_ _4716_/Y _4886_/Y _4906_/B VGND VGND VPWR VPWR _5224_/A sky130_fd_sc_hd__o21ai_1
Xhold3008 _6915_/Q VGND VGND VPWR VPWR hold730/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_110_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6191_ _6649_/S _7604_/Q _6777_/S _6190_/X VGND VGND VPWR VPWR _6191_/X sky130_fd_sc_hd__a211o_1
Xhold3019 _7032_/Q VGND VGND VPWR VPWR hold3019/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_1_1__f_user_clock clkbuf_0_user_clock/X VGND VGND VPWR VPWR _4161_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3867__A2 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2307 hold584/X VGND VGND VPWR VPWR _5964_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5142_ _4956_/A _4690_/Y _4713_/X _4720_/Y _4706_/Y VGND VGND VPWR VPWR _5143_/C
+ sky130_fd_sc_hd__o32a_1
Xhold2318 _6956_/Q VGND VGND VPWR VPWR hold612/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2329 _7388_/Q VGND VGND VPWR VPWR hold965/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1606 _7497_/Q VGND VGND VPWR VPWR hold275/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1617 hold259/X VGND VGND VPWR VPWR _4444_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4419__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1628 hold247/X VGND VGND VPWR VPWR _5915_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5073_ _5073_/A _5073_/B VGND VGND VPWR VPWR _5081_/A sky130_fd_sc_hd__nand2_8
Xhold1639 _4435_/X VGND VGND VPWR VPWR hold254/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4024_ _4024_/A1 _4040_/A _4023_/X VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__o21a_1
XANTENNA__3550__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4292__A2 _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4943__A _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5758__B hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5975_ _5993_/A1 _5975_/A1 _5982_/S VGND VGND VPWR VPWR _5975_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2960_A _7504_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4154__S _6898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4926_ _4932_/B _4954_/C _4929_/A _5260_/D VGND VGND VPWR VPWR _4927_/B sky130_fd_sc_hd__and4_1
XFILLER_0_176_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4857_ _4856_/A _5072_/B _5058_/D VGND VGND VPWR VPWR _4859_/C sky130_fd_sc_hd__and3b_4
X_7645_ _4164_/A1 _7645_/D _4309_/B VGND VGND VPWR VPWR _7645_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3808_ _7305_/Q _5686_/A _5704_/A _7321_/Q _3807_/X VGND VGND VPWR VPWR _3808_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_172_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7576_ _7581_/CLK hold68/X fanout585/X VGND VGND VPWR VPWR _7576_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_117_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5544__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4788_ _4790_/C _5089_/B _4823_/C VGND VGND VPWR VPWR _5096_/A sky130_fd_sc_hd__and3_4
XANTENNA__6741__B2 _7185_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6527_ _7370_/Q _6459_/B _6651_/C _6455_/X _7458_/Q VGND VGND VPWR VPWR _6527_/X
+ sky130_fd_sc_hd__a32o_1
X_3739_ _7290_/Q _4212_/A _3669_/C _4322_/A _7004_/Q VGND VGND VPWR VPWR _3739_/X
+ sky130_fd_sc_hd__a32o_1
X_6458_ _7431_/Q _6747_/B _6645_/C _6457_/X _7471_/Q VGND VGND VPWR VPWR _6458_/X
+ sky130_fd_sc_hd__a32o_1
X_5409_ _4687_/Y _5406_/Y _4761_/Y _5140_/X _5303_/D VGND VGND VPWR VPWR _5569_/A
+ sky130_fd_sc_hd__o311a_1
X_6389_ _7030_/Q _6099_/X _6111_/X _7040_/Q _6388_/X VGND VGND VPWR VPWR _6389_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2830 hold2830/A VGND VGND VPWR VPWR _5840_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2841 _6874_/Q VGND VGND VPWR VPWR hold2841/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2852 _6972_/Q VGND VGND VPWR VPWR _4278_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2863 hold2863/A VGND VGND VPWR VPWR hold2863/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2874 _7127_/Q VGND VGND VPWR VPWR hold2874/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2885 hold2885/A VGND VGND VPWR VPWR _5868_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2896 hold2896/A VGND VGND VPWR VPWR hold2896/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5480__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5480__B2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3491__B1 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5668__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4572__B _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5387__C _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3546__A1 _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3546__B2 _7350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5299__A1 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6496__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__A2 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4747__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6248__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3651__B _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4239__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6799__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6799__B2 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6263__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4663__B1_N _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5471__A1 _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5760_ hold43/X _5760_/A1 _5766_/S VGND VGND VPWR VPWR _5760_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_174_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4711_ _4753_/C _4767_/B VGND VGND VPWR VPWR _5404_/B sky130_fd_sc_hd__and2_2
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5691_ hold84/X _5691_/A1 _5694_/S VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__mux2_1
XFILLER_0_126_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7430_ _7555_/CLK _7430_/D fanout594/X VGND VGND VPWR VPWR _7430_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2374_A _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4642_ _4675_/A _4675_/B _4643_/C _4645_/D VGND VGND VPWR VPWR _4648_/A sky130_fd_sc_hd__nand4_4
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7361_ _7537_/CLK _7361_/D fanout575/X VGND VGND VPWR VPWR _7361_/Q sky130_fd_sc_hd__dfrtp_4
X_4573_ _5058_/D _4888_/B _5282_/A VGND VGND VPWR VPWR _4667_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_141_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap400 _4758_/B VGND VGND VPWR VPWR _5328_/A sky130_fd_sc_hd__buf_6
XFILLER_0_188_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold703 hold703/A VGND VGND VPWR VPWR _7264_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold714 hold714/A VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6312_ _7042_/Q _6089_/X _6308_/X _6309_/X _6311_/X VGND VGND VPWR VPWR _6312_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3545__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3524_ _3524_/A _3524_/B _3524_/C _3524_/D VGND VGND VPWR VPWR _3570_/B sky130_fd_sc_hd__nor4_2
Xhold725 _5796_/X VGND VGND VPWR VPWR _7400_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7292_ _7366_/CLK _7292_/D fanout579/X VGND VGND VPWR VPWR _7292_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold736 hold736/A VGND VGND VPWR VPWR hold736/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold747 hold747/A VGND VGND VPWR VPWR hold747/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap455 _4815_/B VGND VGND VPWR VPWR _4790_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__6487__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold758 hold758/A VGND VGND VPWR VPWR _7435_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold769 hold769/A VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6243_ _7381_/Q _6089_/X _6239_/X _6240_/X _6242_/X VGND VGND VPWR VPWR _6243_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ _6904_/Q hold396/X _4025_/A VGND VGND VPWR VPWR _3455_/X sky130_fd_sc_hd__mux2_1
Xhold2104 _5844_/X VGND VGND VPWR VPWR hold148/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6174_ _7378_/Q _6089_/X _6144_/C _6173_/X VGND VGND VPWR VPWR _6174_/X sky130_fd_sc_hd__a31o_1
Xhold2115 _6935_/Q VGND VGND VPWR VPWR hold799/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2126 _7126_/Q VGND VGND VPWR VPWR hold149/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3561__B _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6239__B1 _6093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2137 hold2137/A VGND VGND VPWR VPWR _4460_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5125_ _4851_/Y _5294_/A _5064_/Y _4968_/X _5124_/X VGND VGND VPWR VPWR _5125_/Y
+ sky130_fd_sc_hd__a221oi_2
Xhold1403 hold5/X VGND VGND VPWR VPWR _5735_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4149__S _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2148 _4472_/X VGND VGND VPWR VPWR hold168/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2159 hold169/X VGND VGND VPWR VPWR _4445_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1414 _5968_/X VGND VGND VPWR VPWR hold1414/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1425 hold194/X VGND VGND VPWR VPWR _7329_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4376__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1436 _5725_/X VGND VGND VPWR VPWR hold202/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1447 _3569_/X VGND VGND VPWR VPWR _5893_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6254__A3 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5056_ _5056_/A _5056_/B _5056_/C VGND VGND VPWR VPWR _5060_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_137_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1458 hold178/X VGND VGND VPWR VPWR _7270_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1469 _3543_/X VGND VGND VPWR VPWR _5668_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4007_ _4062_/A _4025_/A VGND VGND VPWR VPWR _4040_/D sky130_fd_sc_hd__nand2_4
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout457_A _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7219__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7556__RESET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6411__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4823__D _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5958_ _5958_/A0 _5985_/A1 _5964_/S VGND VGND VPWR VPWR _5958_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3776__A1 _6965_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4909_ _4909_/A _4929_/A _4909_/C _4909_/D VGND VGND VPWR VPWR _4915_/C sky130_fd_sc_hd__and4_2
X_5889_ _5889_/A0 _5997_/A1 _5892_/S VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__mux2_1
X_7628_ _7644_/CLK _7628_/D _4309_/B VGND VGND VPWR VPWR _7628_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3528__A1 _7510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3528__B2 _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6190__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6112__B _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7559_ _7563_/CLK _7559_/D fanout602/X VGND VGND VPWR VPWR _7559_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_132_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1739_A _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input157_A wb_dat_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4567__B _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3700__B2 _7201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2660 _5850_/X VGND VGND VPWR VPWR _7448_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2671 _7475_/Q VGND VGND VPWR VPWR hold742/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2682 _5817_/X VGND VGND VPWR VPWR hold768/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2693 hold761/X VGND VGND VPWR VPWR _5826_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1970 _4368_/X VGND VGND VPWR VPWR hold423/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input18_A mask_rev_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1981 _4477_/X VGND VGND VPWR VPWR hold453/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1992 _5815_/X VGND VGND VPWR VPWR hold550/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_97_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3767__A1 _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3767__B2 _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6705__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6705__B2 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3646__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6181__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4192__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_5 _3725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6469__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4758__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3662__A _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5141__B1 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6641__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6930_ _7601_/CLK _6930_/D fanout565/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfrtp_4
X_6861_ _6873_/A _6869_/B VGND VGND VPWR VPWR _6861_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_6_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7211_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4643__D _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5812_ _5866_/B _5884_/B hold48/A VGND VGND VPWR VPWR _5820_/S sky130_fd_sc_hd__and3_4
X_6792_ _3570_/Y _6792_/A1 _6792_/S VGND VGND VPWR VPWR _7636_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3758__A1 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5743_ _5743_/A0 _5896_/A0 _5748_/S VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5674_ _5953_/A1 _5674_/A1 _5676_/S VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3556__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7413_ _7478_/CLK _7413_/D fanout581/X VGND VGND VPWR VPWR _7413_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4625_ _5058_/D _4856_/A _5399_/A VGND VGND VPWR VPWR _4956_/A sky130_fd_sc_hd__nand3_4
XANTENNA__6172__A2 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7344_ _7539_/CLK _7344_/D fanout578/X VGND VGND VPWR VPWR _7344_/Q sky130_fd_sc_hd__dfstp_2
Xhold500 hold500/A VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4556_ _5586_/A0 _4556_/A1 _4556_/S VGND VGND VPWR VPWR _4556_/X sky130_fd_sc_hd__mux2_1
Xhold511 hold511/A VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold522 hold522/A VGND VGND VPWR VPWR hold522/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold533 _5715_/X VGND VGND VPWR VPWR _7328_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3507_ _3507_/A hold20/A _4491_/C VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__and3_4
Xhold544 hold544/A VGND VGND VPWR VPWR _7470_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7275_ _7429_/CLK _7275_/D fanout583/X VGND VGND VPWR VPWR _7275_/Q sky130_fd_sc_hd__dfrtp_1
Xhold555 hold555/A VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4487_ _5805_/A1 _4487_/A1 _4490_/S VGND VGND VPWR VPWR _4487_/X sky130_fd_sc_hd__mux2_1
Xhold566 hold566/A VGND VGND VPWR VPWR _7322_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold577 _5706_/X VGND VGND VPWR VPWR _7320_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold588 hold588/A VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6226_ _7300_/Q _6074_/X _6379_/B1 _7396_/Q _6225_/X VGND VGND VPWR VPWR _6226_/X
+ sky130_fd_sc_hd__a221o_1
X_3438_ _7338_/Q VGND VGND VPWR VPWR _3438_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6475__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold599 hold599/A VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5683__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6152_/X _6157_/B _6157_/C VGND VGND VPWR VPWR _6157_/Y sky130_fd_sc_hd__nand3b_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout574_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1200 hold1200/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
Xhold1211 hold2840/X VGND VGND VPWR VPWR hold1211/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 hold3061/X VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5108_ _5107_/A _4743_/Y wire529/X _5107_/X VGND VGND VPWR VPWR _5111_/B sky130_fd_sc_hd__a31o_1
XANTENNA__6227__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1233 hold2964/X VGND VGND VPWR VPWR hold2965/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1244 _5622_/X VGND VGND VPWR VPWR _7249_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6088_ _7495_/Q _6085_/X _6087_/X _7463_/Q _6083_/X VGND VGND VPWR VPWR _6102_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1255 hold3066/X VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1266 hold3119/X VGND VGND VPWR VPWR hold3120/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6632__B1 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1277 hold3115/X VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5039_ _5039_/A _5039_/B _5039_/C VGND VGND VPWR VPWR _5041_/A sky130_fd_sc_hd__nor3_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 hold3144/X VGND VGND VPWR VPWR hold3145/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1299 _4365_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3749__B2 _7034_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1856_A _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6699__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6163__A2 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4578__A _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3482__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR _4089_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput131 wb_cyc_i VGND VGND VPWR VPWR _4093_/A sky130_fd_sc_hd__clkbuf_2
Xhold3180 _3797_/X VGND VGND VPWR VPWR _7217_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5901__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6809_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3191 _6701_/X VGND VGND VPWR VPWR _7624_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6814_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_4
XANTENNA__4857__A_N _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5426__A1 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2490 hold963/X VGND VGND VPWR VPWR _4186_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6623__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6387__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3657__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6154__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4410_ _4442_/A0 _5985_/A1 _4422_/S VGND VGND VPWR VPWR _4410_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4165__A1 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5390_ _5390_/A _5518_/C _5473_/C VGND VGND VPWR VPWR _5394_/A sky130_fd_sc_hd__and3_1
XFILLER_0_111_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4341_ _5714_/A0 _4341_/A1 _4345_/S VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7060_ _7170_/CLK _7060_/D fanout573/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4272_ _4272_/A0 _5840_/A1 _4276_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6011_ _7585_/Q _7584_/Q _6932_/Q _6751_/S VGND VGND VPWR VPWR _6011_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5665__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5811__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2504_A _7400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3691__A3 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3979__A1 _7439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6913_ _6926_/CLK _6913_/D fanout566/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_178_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6844_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6844_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6775_ _6961_/Q _6431_/Y _6775_/B1 VGND VGND VPWR VPWR _6775_/X sky130_fd_sc_hd__o21a_1
X_3987_ _7287_/Q _3543_/X _3983_/X _3985_/X _3986_/X VGND VGND VPWR VPWR _3988_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_190_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5726_ _5726_/A0 _5987_/A1 _5730_/S VGND VGND VPWR VPWR _5726_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3600__B1 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5657_ _5954_/A1 _5657_/A1 _5658_/S VGND VGND VPWR VPWR _5657_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4156__A1 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4608_ _4887_/D _4747_/B _4887_/B _4879_/C VGND VGND VPWR VPWR _4608_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_142_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5588_ _5588_/A0 _5948_/A1 _5589_/S VGND VGND VPWR VPWR _5588_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_102_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3903__A1 _7448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold330 hold330/A VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7327_ _7359_/CLK _7327_/D fanout575/X VGND VGND VPWR VPWR _7327_/Q sky130_fd_sc_hd__dfstp_2
X_4539_ hold36/X _5612_/C hold56/X _5902_/B VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__and4_1
Xhold341 hold341/A VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3903__B2 _7440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold352 hold352/A VGND VGND VPWR VPWR hold352/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold363 _5932_/X VGND VGND VPWR VPWR _7521_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold374 hold374/A VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_159_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6448__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold385 _4404_/X VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_159_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold396 _6903_/Q VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7258_ _7578_/CLK _7258_/D fanout604/X VGND VGND VPWR VPWR _7258_/Q sky130_fd_sc_hd__dfrtp_4
X_6209_ _7459_/Q _6080_/X _6092_/X _7531_/Q _6208_/X VGND VGND VPWR VPWR _6209_/X
+ sky130_fd_sc_hd__a221o_1
X_7189_ _7189_/CLK _7189_/D fanout574/X VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfstp_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 _5687_/X VGND VGND VPWR VPWR _7303_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5408__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1041 hold2878/X VGND VGND VPWR VPWR hold2879/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 hold2750/X VGND VGND VPWR VPWR _7271_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6605__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 _4450_/X VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1074 hold2803/X VGND VGND VPWR VPWR hold2804/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 _4273_/X VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5022__A _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 hold2892/X VGND VGND VPWR VPWR hold2893/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4580__B _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6384__A2 _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3187_A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input85_A spimemio_flash_io0_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6788__A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6727__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4855__C1 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_71_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7024_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4247__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4607__C1 _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6611__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3910_ _7496_/Q _5902_/A _3651_/X _7047_/Q _3909_/X VGND VGND VPWR VPWR _3913_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4890_ _5222_/B _5222_/C _5260_/D _4891_/D VGND VGND VPWR VPWR _5223_/D sky130_fd_sc_hd__nand4_2
X_3841_ _7393_/Q _5785_/A _3933_/A _3665_/X _7124_/Q VGND VGND VPWR VPWR _3841_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4921__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5583__A0 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3772_ _7049_/Q _3651_/X _3767_/X _3769_/X _3771_/X VGND VGND VPWR VPWR _3772_/X
+ sky130_fd_sc_hd__a2111o_1
X_6560_ _7379_/Q _6408_/B _6555_/X _6557_/X _6559_/X VGND VGND VPWR VPWR _6570_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_70_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5511_ _4843_/A _4659_/Y _5081_/A _5541_/D _5247_/C VGND VGND VPWR VPWR _5512_/D
+ sky130_fd_sc_hd__o311a_1
X_6491_ _7464_/Q _6434_/X _6460_/X _7384_/Q _6490_/X VGND VGND VPWR VPWR _6494_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5806__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4138__A1 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5442_ _5107_/A _5342_/A _5342_/B _5205_/X VGND VGND VPWR VPWR _5442_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_125_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6678__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5886__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5373_ _4744_/Y _4844_/Y _4880_/Y _4846_/Y VGND VGND VPWR VPWR _5373_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3897__B1 _3889_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7487_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5107__A _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4324_ _5805_/A1 _4324_/A1 _4327_/S VGND VGND VPWR VPWR _4324_/X sky130_fd_sc_hd__mux2_1
X_7112_ _7112_/CLK _7112_/D fanout589/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7043_ _7156_/CLK _7043_/D _6833_/A VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfstp_4
X_4255_ _4255_/A0 _5997_/A1 _4258_/S VGND VGND VPWR VPWR _4255_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4186_ _4186_/A0 _5914_/A1 _4190_/S VGND VGND VPWR VPWR _4186_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4665__B _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7551_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_3_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_1_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5810__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4681__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3821__B1 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6827_ _6827_/A _6827_/B VGND VGND VPWR VPWR _6827_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6366__A2 _6072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4377__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire507 wire508/X VGND VGND VPWR VPWR _4075_/S sky130_fd_sc_hd__buf_6
X_6758_ _7136_/Q _6409_/X _6753_/X _6757_/X _6430_/X VGND VGND VPWR VPWR _6758_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_45_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3719__A4 _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire529 _5072_/D VGND VGND VPWR VPWR wire529/X sky130_fd_sc_hd__buf_2
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5709_ hold84/X _5709_/A1 _5712_/S VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6689_ _7198_/Q _6463_/A _6771_/A3 _6408_/D _7168_/Q VGND VGND VPWR VPWR _6689_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5877__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6120__B _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold160 hold160/A VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold171 hold171/A VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold182 hold182/A VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5629__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold193 hold193/A VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5058__A_N _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4856__A _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4575__B _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__A2 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4368__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output289_A _6923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3591__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5868__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3654__B _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4540__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3894__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3670__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4040_ _4040_/A _6900_/Q _6901_/Q _4040_/D VGND VGND VPWR VPWR _4042_/A sky130_fd_sc_hd__and4_1
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4485__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6045__A1 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2202_A _7302_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6596__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5991_ _5991_/A0 _5991_/A1 _5991_/S VGND VGND VPWR VPWR _5991_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4942_ _4942_/A _5248_/B _4948_/C _5180_/B VGND VGND VPWR VPWR _4944_/B sky130_fd_sc_hd__nand4_1
XANTENNA__3803__B1 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7661_ _7661_/A VGND VGND VPWR VPWR _7661_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6348__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4873_ _4667_/A _4667_/B _4984_/B _4984_/A VGND VGND VPWR VPWR _4873_/X sky130_fd_sc_hd__o22a_4
XFILLER_0_129_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6612_ _7593_/Q _7581_/Q _6408_/C _6611_/X VGND VGND VPWR VPWR _6612_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4359__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3824_ _7252_/Q _5640_/C _5623_/B _3663_/X _7164_/Q VGND VGND VPWR VPWR _3824_/X
+ sky130_fd_sc_hd__a32o_1
X_7592_ _7593_/CLK _7592_/D fanout568/X VGND VGND VPWR VPWR _7592_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_27_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6543_ _7314_/Q _6419_/D _6454_/X _7490_/Q _6542_/X VGND VGND VPWR VPWR _6544_/D
+ sky130_fd_sc_hd__a221o_1
X_3755_ _4168_/D _4248_/S _3652_/X _7150_/Q VGND VGND VPWR VPWR _3755_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3582__A2 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3686_ _7233_/Q _3617_/X _3681_/X _3683_/X _3685_/X VGND VGND VPWR VPWR _3686_/X
+ sky130_fd_sc_hd__a2111o_2
X_6474_ _7593_/Q _7576_/Q _6408_/C _6058_/X _7528_/Q VGND VGND VPWR VPWR _6474_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3564__B _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput210 _3438_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
X_5425_ _5282_/A _5339_/A _5199_/C _4758_/X VGND VGND VPWR VPWR _5425_/X sky130_fd_sc_hd__a31o_2
Xoutput221 _7659_/X VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6520__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput232 _7669_/X VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput243 _4152_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XANTENNA__4531__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput254 _4132_/Y VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
X_5356_ _5094_/A _5183_/C _4877_/A VGND VGND VPWR VPWR _5450_/B sky130_fd_sc_hd__o21ai_1
Xoutput265 _7222_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
Xoutput276 _7235_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
XFILLER_0_11_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput287 _6921_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XANTENNA__3885__A3 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4307_ _4307_/A0 _5647_/A0 _4308_/S VGND VGND VPWR VPWR _4307_/X sky130_fd_sc_hd__mux2_1
Xoutput298 _7247_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
X_5287_ _5061_/B _5453_/C _4845_/X VGND VGND VPWR VPWR _5294_/B sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout487_A _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4238_ _5653_/A1 _5896_/A0 _4248_/S VGND VGND VPWR VPWR _4238_/X sky130_fd_sc_hd__mux2_1
X_7026_ _7196_/CLK _7026_/D fanout590/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfrtp_4
X_4169_ _7084_/Q _4169_/A2 _4168_/Y _4169_/B2 VGND VGND VPWR VPWR _4169_/X sky130_fd_sc_hd__a22o_2
XANTENNA__4047__A0 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6587__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5795__A0 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5938__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire348 _6440_/Y VGND VGND VPWR VPWR wire348/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6511__A2 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4522__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3876__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input48_A mgmt_gpio_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3490__A _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6275__A1 _7470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6275__B2 _7510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout470 hold1662/X VGND VGND VPWR VPWR hold1663/A sky130_fd_sc_hd__buf_6
Xfanout481 _5735_/A1 VGND VGND VPWR VPWR _5987_/A1 sky130_fd_sc_hd__clkbuf_16
XANTENNA__3628__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5483__C1 _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout492 _5940_/A1 VGND VGND VPWR VPWR _5985_/A1 sky130_fd_sc_hd__buf_12
XANTENNA__4598__A_N _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6290__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3649__B hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5250__A2 _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3800__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3665__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3540_ _7438_/Q _3525_/X _3528_/X _3534_/X _3539_/X VGND VGND VPWR VPWR _3568_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_51_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold907 hold907/A VGND VGND VPWR VPWR hold907/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold918 _4519_/X VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold929 hold929/A VGND VGND VPWR VPWR hold929/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3471_ _3507_/A hold20/X VGND VGND VPWR VPWR _3537_/A sky130_fd_sc_hd__and2_4
XANTENNA__6502__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5210_ _4601_/Y _4716_/Y _4726_/Y _4906_/B VGND VGND VPWR VPWR _5210_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5710__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4513__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6190_ _7282_/Q _6036_/Y _6178_/X _6189_/X _6775_/B1 VGND VGND VPWR VPWR _6190_/X
+ sky130_fd_sc_hd__o221a_1
Xhold3009 hold730/X VGND VGND VPWR VPWR _4196_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_20_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5141_ _4706_/Y _4741_/Y _4759_/Y _4761_/Y _5139_/X VGND VGND VPWR VPWR _5143_/B
+ sky130_fd_sc_hd__o221a_1
Xhold2308 _5964_/X VGND VGND VPWR VPWR hold585/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2319 hold612/X VGND VGND VPWR VPWR _4258_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5072_ _5399_/B _5072_/B _5072_/C _5072_/D VGND VGND VPWR VPWR _5072_/Y sky130_fd_sc_hd__nand4_1
Xhold1607 hold275/X VGND VGND VPWR VPWR _5905_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1618 _4444_/X VGND VGND VPWR VPWR hold260/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1629 _5915_/X VGND VGND VPWR VPWR hold248/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4023_ _4028_/A0 _4025_/A _4022_/X VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5777__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5974_ hold72/X _5992_/D VGND VGND VPWR VPWR _5982_/S sky130_fd_sc_hd__nand2_8
XANTENNA__3788__C1 _3787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4925_ _4925_/A _5444_/C _4925_/C VGND VGND VPWR VPWR _4927_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_136_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6650__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7644_ _7644_/CLK _7644_/D _6780_/B VGND VGND VPWR VPWR _7644_/Q sky130_fd_sc_hd__dfrtp_1
X_4856_ _4856_/A _4888_/B _5058_/D VGND VGND VPWR VPWR _4856_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_0_145_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3807_ _6990_/Q _5731_/B _5623_/B _3531_/X _7337_/Q VGND VGND VPWR VPWR _3807_/X
+ sky130_fd_sc_hd__a32o_1
X_7575_ _7575_/CLK _7575_/D fanout595/X VGND VGND VPWR VPWR _7575_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6741__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4787_ _4836_/C _4797_/B VGND VGND VPWR VPWR _4787_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6526_ _7562_/Q _6419_/C _6466_/X _7506_/Q _6525_/X VGND VGND VPWR VPWR _6526_/X
+ sky130_fd_sc_hd__a221o_1
X_3738_ _7261_/Q _5619_/B _5659_/B VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__and3_1
X_6457_ _7595_/Q _6574_/B _6600_/B _7596_/Q VGND VGND VPWR VPWR _6457_/X sky130_fd_sc_hd__and4b_4
X_3669_ _4491_/A _4491_/C _3669_/C VGND VGND VPWR VPWR _3669_/X sky130_fd_sc_hd__and3_4
XFILLER_0_30_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4504__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5408_ _5113_/A _5295_/C _5410_/A VGND VGND VPWR VPWR _5408_/Y sky130_fd_sc_hd__o21ai_2
X_6388_ _7060_/Q _6110_/A _6084_/X _6082_/X _7010_/Q VGND VGND VPWR VPWR _6388_/X
+ sky130_fd_sc_hd__a32o_1
X_5339_ _5339_/A _5339_/B _5339_/C _5339_/D VGND VGND VPWR VPWR _5340_/A sky130_fd_sc_hd__nand4_2
Xhold2820 hold2820/A VGND VGND VPWR VPWR hold2820/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2831 _5840_/X VGND VGND VPWR VPWR hold2831/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2842 hold2842/A VGND VGND VPWR VPWR _4182_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2853 hold2853/A VGND VGND VPWR VPWR hold2853/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2864 _7147_/Q VGND VGND VPWR VPWR hold2864/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5014__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2875 hold2875/A VGND VGND VPWR VPWR _4468_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7009_ _7190_/CLK _7009_/D fanout573/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2886 _5868_/X VGND VGND VPWR VPWR hold2886/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2897 _6950_/Q VGND VGND VPWR VPWR hold2897/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4853__B _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5030__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4572__C _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input102_A wb_adr_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4440__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5965__A _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6193__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6732__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3546__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5904__S _5910_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5299__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__C _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3651__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5471__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5759__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6036__A _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5875__A _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _5113_/A _5089_/B _5089_/C VGND VGND VPWR VPWR _4803_/A sky130_fd_sc_hd__and3_2
XANTENNA_clkbuf_leaf_29_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3785__A2 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5690_ _5951_/A1 _5690_/A1 _5694_/S VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4641_ _4694_/B _4641_/B _4730_/C _4768_/B VGND VGND VPWR VPWR _4811_/A sky130_fd_sc_hd__nor4_2
XFILLER_0_142_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6723__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2367_A _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5931__A0 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7360_ _7537_/CLK _7360_/D fanout577/X VGND VGND VPWR VPWR _7360_/Q sky130_fd_sc_hd__dfstp_2
X_4572_ _5058_/D _4888_/B _5282_/A VGND VGND VPWR VPWR _4668_/C sky130_fd_sc_hd__and3_4
XFILLER_0_188_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap401 _4647_/Y VGND VGND VPWR VPWR _5222_/B sky130_fd_sc_hd__buf_6
XFILLER_0_25_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold704 hold704/A VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6311_ _7113_/Q _6317_/C _6074_/X _6968_/Q _6310_/X VGND VGND VPWR VPWR _6311_/X
+ sky130_fd_sc_hd__a221o_1
Xhold715 hold715/A VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold56_A hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3523_ _7374_/Q _5758_/A _3519_/X _7550_/Q _3522_/X VGND VGND VPWR VPWR _3524_/D
+ sky130_fd_sc_hd__a221o_1
X_7291_ _7539_/CLK hold85/X fanout577/X VGND VGND VPWR VPWR _7291_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold726 hold726/A VGND VGND VPWR VPWR hold726/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold737 hold737/A VGND VGND VPWR VPWR _7250_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5814__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap456 _5059_/B VGND VGND VPWR VPWR _4815_/B sky130_fd_sc_hd__buf_4
Xhold748 _4363_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold759 hold759/A VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6242_ _7389_/Q _6317_/C _6379_/B1 _7397_/Q _6241_/X VGND VGND VPWR VPWR _6242_/X
+ sky130_fd_sc_hd__a221o_1
X_3454_ _4429_/B hold52/X hold529/X VGND VGND VPWR VPWR _3454_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4498__A0 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6173_ _7410_/Q _6144_/C _6097_/B _6144_/B VGND VGND VPWR VPWR _6173_/X sky130_fd_sc_hd__o211a_1
Xhold2105 _7156_/Q VGND VGND VPWR VPWR hold158/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2116 hold799/X VGND VGND VPWR VPWR _4222_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5115__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2127 hold149/X VGND VGND VPWR VPWR _4466_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2138 _4460_/X VGND VGND VPWR VPWR hold157/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3561__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5124_ _5122_/Y _5123_/X _5580_/A2 VGND VGND VPWR VPWR _5124_/X sky130_fd_sc_hd__a21o_1
Xhold2149 _7451_/Q VGND VGND VPWR VPWR hold141/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1404 _5735_/X VGND VGND VPWR VPWR hold1404/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1415 _7646_/Q VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1426 _7473_/Q VGND VGND VPWR VPWR hold221/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4376__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1437 hold202/X VGND VGND VPWR VPWR _7337_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5055_ _5295_/A _5113_/A _5118_/C _5295_/D VGND VGND VPWR VPWR _5056_/C sky130_fd_sc_hd__nand4_1
Xhold1448 _5893_/Y VGND VGND VPWR VPWR _5901_/S sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1459 _7516_/Q VGND VGND VPWR VPWR hold171/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_137_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4006_ _4006_/A _4006_/B VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__nor2_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4670__B1 _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5214__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6411__A1 _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5957_ _5957_/A0 _5993_/A1 _5964_/S VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5785__A _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3776__A2 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4973__A1 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4908_ wire533/X _4877_/A _4907_/X _4906_/Y VGND VGND VPWR VPWR _4913_/A sky130_fd_sc_hd__a211oi_1
XANTENNA_fanout617_A _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5888_ _5888_/A0 _5996_/A1 _5892_/S VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7627_ _7627_/CLK _7627_/D fanout566/X VGND VGND VPWR VPWR _7627_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6175__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4839_ _5011_/B _4839_/B VGND VGND VPWR VPWR _5496_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6714__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5922__A0 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3528__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7558_ _7582_/CLK hold32/X fanout585/X VGND VGND VPWR VPWR _7558_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_160_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6509_ _7313_/Q _6419_/D _6424_/X _7569_/Q _6508_/X VGND VGND VPWR VPWR _6509_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7489_ _7489_/CLK _7489_/D fanout586/X VGND VGND VPWR VPWR _7489_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5724__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6478__A1 _7400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4489__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3700__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__clkbuf_4
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2650 _5970_/X VGND VGND VPWR VPWR hold689/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2661 _7523_/Q VGND VGND VPWR VPWR hold734/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2672 hold742/X VGND VGND VPWR VPWR _5880_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2683 _6940_/Q VGND VGND VPWR VPWR hold893/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2694 _5826_/X VGND VGND VPWR VPWR hold762/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1960 _7361_/Q VGND VGND VPWR VPWR hold553/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1971 hold423/X VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4583__B _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1982 hold453/X VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4661__B1 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1993 _7155_/Q VGND VGND VPWR VPWR hold478/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_168_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5205__A2 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5695__A _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3767__A2 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3927__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6166__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6705__A2 _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4786__A_N _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3646__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_6 _3774_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6469__A1 _7367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6469__B2 _7407_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4758__B _4758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3662__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4774__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6641__B2 _7366_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4924__D _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6860_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6860_/X sky130_fd_sc_hd__and2_1
XFILLER_0_190_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_187_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5811_ _5811_/A0 _5955_/A1 _5811_/S VGND VGND VPWR VPWR _5811_/X sky130_fd_sc_hd__mux2_1
X_6791_ _3607_/Y _6791_/A1 _6792_/S VGND VGND VPWR VPWR _7635_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5809__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3758__A2 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5742_ _5742_/A0 _5985_/A1 _5748_/S VGND VGND VPWR VPWR _5742_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4955__B2 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4940__C _4940_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5673_ hold84/X _5673_/A1 _5676_/S VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__mux2_1
XFILLER_0_155_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7412_ _7412_/CLK _7412_/D fanout581/X VGND VGND VPWR VPWR _7412_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5904__A0 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3556__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4624_ _5058_/D _4856_/A _5399_/A VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__and3_4
XFILLER_0_114_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7343_ _7537_/CLK _7343_/D fanout577/X VGND VGND VPWR VPWR _7343_/Q sky130_fd_sc_hd__dfstp_2
Xhold501 hold501/A VGND VGND VPWR VPWR _7272_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4555_ _5852_/A0 _4555_/A1 _4556_/S VGND VGND VPWR VPWR _4555_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold512 hold512/A VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold523 hold523/A VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold534 hold534/A VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold545 hold545/A VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3506_ _4473_/A hold22/A _3931_/D VGND VGND VPWR VPWR _3506_/X sky130_fd_sc_hd__and3_4
X_7274_ _7278_/CLK _7274_/D fanout580/X VGND VGND VPWR VPWR _7274_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold556 _5892_/X VGND VGND VPWR VPWR _7486_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4486_ _5948_/A1 _4486_/A1 _4490_/S VGND VGND VPWR VPWR _4486_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4668__B _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold567 hold567/A VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold578 hold578/A VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5132__A1 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold589 _5688_/X VGND VGND VPWR VPWR _7304_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6225_ _7292_/Q _6144_/A _6136_/C _6332_/C _7364_/Q VGND VGND VPWR VPWR _6225_/X
+ sky130_fd_sc_hd__a32o_1
X_3437_ _7346_/Q VGND VGND VPWR VPWR _3437_/Y sky130_fd_sc_hd__inv_2
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _7369_/Q _6111_/X _6121_/X _7305_/Q _6155_/X VGND VGND VPWR VPWR _6157_/C
+ sky130_fd_sc_hd__a221oi_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 hold2861/X VGND VGND VPWR VPWR hold1201/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 hold1212/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 hold3033/X VGND VGND VPWR VPWR hold3034/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5107_ _5107_/A _5118_/A _5387_/C VGND VGND VPWR VPWR _5107_/X sky130_fd_sc_hd__and3_1
Xhold1234 hold3088/X VGND VGND VPWR VPWR hold3089/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6087_ _6110_/A _6121_/A _6120_/B VGND VGND VPWR VPWR _6087_/X sky130_fd_sc_hd__and3_4
XANTENNA_fanout567_A fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1245 _4078_/A VGND VGND VPWR VPWR _4406_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1256 hold3148/X VGND VGND VPWR VPWR hold3149/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1267 hold3121/X VGND VGND VPWR VPWR _7423_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1278 hold3100/X VGND VGND VPWR VPWR hold3101/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5038_ _5038_/A _5038_/B _5038_/C VGND VGND VPWR VPWR _5039_/B sky130_fd_sc_hd__and3_1
Xhold1289 _5741_/X VGND VGND VPWR VPWR _7351_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5011__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6989_ _7409_/CLK _6989_/D fanout577/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4850__C _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6148__B1 _6116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4859__A _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3482__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5123__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6320__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR input110/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR _4945_/A sky130_fd_sc_hd__clkbuf_8
Xhold3170 _6919_/Q VGND VGND VPWR VPWR hold3170/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6800_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input30_A mask_rev_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3181 _7106_/Q VGND VGND VPWR VPWR _4425_/C sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6803_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3192 _7643_/Q VGND VGND VPWR VPWR _6819_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6806_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6793_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2480 hold658/X VGND VGND VPWR VPWR _4261_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5426__A2 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2491 _4186_/X VGND VGND VPWR VPWR hold964/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4634__B1 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1790 _5797_/X VGND VGND VPWR VPWR hold403/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6387__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3673__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2065_A _7528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4340_ _4340_/A _5902_/B VGND VGND VPWR VPWR _4345_/S sky130_fd_sc_hd__nand2_4
XANTENNA__3912__A2 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4271_ _4551_/C _4491_/C _4352_/A _4551_/D VGND VGND VPWR VPWR _4276_/S sky130_fd_sc_hd__and4_4
XANTENNA__6311__B1 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6010_ _7585_/Q _7584_/Q VGND VGND VPWR VPWR _6010_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6912_ _6926_/CLK _6912_/D fanout565/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_77_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6843_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6843_/X sky130_fd_sc_hd__and2_1
XFILLER_0_175_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4443__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2866_A _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6774_ _6758_/X _6774_/B _6774_/C VGND VGND VPWR VPWR _6774_/Y sky130_fd_sc_hd__nand3b_4
X_3986_ _7415_/Q _3544_/X _3565_/X _7463_/Q _3925_/X VGND VGND VPWR VPWR _3986_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6393__A3 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5725_ _5725_/A0 _5896_/A0 _5730_/S VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5656_ _5863_/A0 _5656_/A1 _5656_/S VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_142_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4607_ _4887_/D _4747_/B _4887_/B _4879_/C VGND VGND VPWR VPWR _4645_/D sky130_fd_sc_hd__o211a_4
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6550__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5587_ hold36/X _5722_/A _5587_/C _5640_/D VGND VGND VPWR VPWR _5589_/S sky130_fd_sc_hd__and4_1
XFILLER_0_115_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold320 hold320/A VGND VGND VPWR VPWR hold320/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7326_ _7478_/CLK _7326_/D fanout583/X VGND VGND VPWR VPWR _7326_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold331 _5897_/X VGND VGND VPWR VPWR _7490_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3903__A2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4538_ _5586_/A0 _4538_/A1 _4538_/S VGND VGND VPWR VPWR _4538_/X sky130_fd_sc_hd__mux2_1
Xhold342 hold342/A VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold353 _4530_/X VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold364 hold364/A VGND VGND VPWR VPWR hold364/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold375 _4403_/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6302__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7257_ _7578_/CLK _7257_/D fanout595/X VGND VGND VPWR VPWR _7257_/Q sky130_fd_sc_hd__dfrtp_4
Xhold386 hold386/A VGND VGND VPWR VPWR hold386/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4469_ _5940_/A1 _4469_/A1 _4472_/S VGND VGND VPWR VPWR _4469_/X sky130_fd_sc_hd__mux2_1
Xhold397 _3455_/X VGND VGND VPWR VPWR _3456_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6208_ _7427_/Q _6110_/A _6074_/X _6100_/X _7475_/Q VGND VGND VPWR VPWR _6208_/X
+ sky130_fd_sc_hd__a32o_1
X_7188_ _7190_/CLK _7188_/D fanout574/X VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _7400_/Q _6091_/X _6116_/B _7312_/Q _6116_/X VGND VGND VPWR VPWR _6139_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 _4353_/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_175_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1031 hold2907/X VGND VGND VPWR VPWR hold2908/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4845__C _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5408__A2 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1042 _5931_/X VGND VGND VPWR VPWR _7520_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 hold2774/X VGND VGND VPWR VPWR hold2775/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1064 hold2821/X VGND VGND VPWR VPWR hold2822/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 _4480_/X VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 hold2866/X VGND VGND VPWR VPWR hold2867/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 hold2894/X VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_169_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5022__B _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1799_A _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6369__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6384__A3 _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5592__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3082_A _7527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input78_A spi_csb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5344__A1 _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6541__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7212_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_output234_A _4146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4607__B1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3668__A _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3840_ _7184_/Q _4533_/A _4497_/A _7154_/Q _3839_/X VGND VGND VPWR VPWR _3840_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3771_ _7498_/Q _5902_/A _5581_/A _7212_/Q _3770_/X VGND VGND VPWR VPWR _3771_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ _5510_/A _5510_/B _5510_/C VGND VGND VPWR VPWR _5548_/A sky130_fd_sc_hd__and3_1
XFILLER_0_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6490_ _7496_/Q _6447_/C _6429_/X _6419_/C _7560_/Q VGND VGND VPWR VPWR _6490_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6127__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5441_ _5343_/B _5343_/A _5441_/C _5506_/D VGND VGND VPWR VPWR _5441_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__6532__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5372_ _5252_/A _5370_/Y _5371_/X _4854_/X VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_100_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7111_ _7207_/CLK _7111_/D _4309_/B VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_4
X_4323_ _5714_/A0 _4323_/A1 _4327_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5822__S _5829_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7042_ _7201_/CLK _7042_/D _6833_/A VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_4
X_4254_ _4254_/A0 _5987_/A1 _4258_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4946__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4185_ _4185_/A0 _7639_/Q _4429_/B VGND VGND VPWR VPWR _4185_/X sky130_fd_sc_hd__mux2_4
XANTENNA__7369__RESET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3821__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3821__B2 _7449_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6826_ _7109_/Q _6824_/C _6795_/B _6825_/X VGND VGND VPWR VPWR _6826_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout432_A _6404_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6366__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6757_ _7181_/Q _6058_/X _6755_/X _6756_/X VGND VGND VPWR VPWR _6757_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_163_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_77_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3969_ _7026_/Q _3669_/C _5632_/B _3659_/X _7006_/Q VGND VGND VPWR VPWR _3969_/X
+ sky130_fd_sc_hd__a32o_1
Xwire508 _4058_/Y VGND VGND VPWR VPWR wire508/X sky130_fd_sc_hd__buf_4
XANTENNA__6771__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5708_ _5951_/A1 _5708_/A1 _5712_/S VGND VGND VPWR VPWR _5708_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6688_ _7153_/Q _6467_/X _6683_/X _6685_/X _6687_/X VGND VGND VPWR VPWR _6698_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5639_ hold464/X _5639_/A1 _5639_/S VGND VGND VPWR VPWR _5639_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3888__A1 _7512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6120__C _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold150 hold150/A VGND VGND VPWR VPWR hold150/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7309_ _7309_/CLK _7309_/D fanout579/X VGND VGND VPWR VPWR _7309_/Q sky130_fd_sc_hd__dfrtp_4
Xhold161 hold161/A VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold172 hold172/A VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold183 hold183/A VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5732__S _5739_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6826__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold194 hold194/A VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4856__B _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4575__C _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input132_A wb_dat_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3488__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3812__B2 _6969_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4083__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6762__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5907__S _5910_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3591__A3 _3519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3654__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6817__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6817__B2 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3670__B hold36/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6293__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6045__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5990_ _5990_/A0 hold61/X _5991_/S VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4941_ _4941_/A _4941_/B _4941_/C VGND VGND VPWR VPWR _4944_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4932__D _4940_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7660_ _7660_/A VGND VGND VPWR VPWR _7660_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4872_ _4856_/A _5399_/A _5058_/D VGND VGND VPWR VPWR _4956_/B sky130_fd_sc_hd__nand3b_4
XANTENNA__6348__A3 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6611_ _7437_/Q _6747_/B _6747_/C _6408_/A _7557_/Q VGND VGND VPWR VPWR _6611_/X
+ sky130_fd_sc_hd__a32o_1
X_3823_ _7465_/Q _3565_/X _3651_/X _7048_/Q _3822_/X VGND VGND VPWR VPWR _3828_/C
+ sky130_fd_sc_hd__a221o_1
X_7591_ _7593_/CLK _7591_/D fanout568/X VGND VGND VPWR VPWR _7591_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6753__B1 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5817__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6542_ _7474_/Q _6424_/C _6441_/X _6452_/X _7346_/Q VGND VGND VPWR VPWR _6542_/X
+ sky130_fd_sc_hd__a32o_1
X_3754_ _7514_/Q _5920_/A _3673_/X _7200_/Q _3753_/X VGND VGND VPWR VPWR _3759_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7599__622 VGND VGND VPWR VPWR _7599_/D _7599__622/LO sky130_fd_sc_hd__conb_1
XFILLER_0_113_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6473_ _6472_/X _6775_/B1 _6931_/Q _6777_/S _6473_/B2 VGND VGND VPWR VPWR _6473_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6505__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3685_ _7161_/Q hold56/A _5632_/B _3684_/X VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_112_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2829_A _7439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3564__C _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5424_ _4956_/A _4687_/Y _4726_/Y _4880_/Y VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__o22a_1
Xoutput200 _3413_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput211 _3437_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _4155_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_23_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput233 _7649_/X VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
XFILLER_0_112_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput244 _7653_/X VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
X_5355_ _5355_/A _5355_/B _5355_/C _5355_/D VGND VGND VPWR VPWR _5361_/A sky130_fd_sc_hd__and4_1
Xoutput255 _7232_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
XFILLER_0_100_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput266 _7229_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
XANTENNA__6808__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput277 _7236_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XANTENNA__6808__B2 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4306_ _4306_/A0 _5950_/A1 _4308_/S VGND VGND VPWR VPWR _4306_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput288 _6922_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_0_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput299 _3929_/Y VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
XANTENNA__7496__CLK _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5286_ _5222_/A _5107_/A _5342_/A _5285_/X VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__a31o_1
X_7025_ _7409_/CLK _7025_/D fanout568/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_4
X_4237_ _4237_/A0 _4236_/X _4249_/S VGND VGND VPWR VPWR _4237_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout382_A _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4295__A1 _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6823__A4 _4428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4168_ _7084_/Q _7257_/Q _7306_/Q _4168_/D VGND VGND VPWR VPWR _4168_/Y sky130_fd_sc_hd__nor4_2
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4692__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4099_ _4099_/A _7586_/Q _7587_/Q _4099_/D VGND VGND VPWR VPWR _4099_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_78_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6809_ _7109_/Q _6809_/A2 _6809_/B1 wire463/A _6808_/X VGND VGND VPWR VPWR _6809_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6744__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5727__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6412__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire349 _6118_/Y VGND VGND VPWR VPWR _6122_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7239_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1929_A _6916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3730__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3490__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6275__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4286__A1 _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout471 _5863_/A0 VGND VGND VPWR VPWR _5953_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout482 _5735_/A1 VGND VGND VPWR VPWR _5996_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout493 hold43/X VGND VGND VPWR VPWR _5940_/A1 sky130_fd_sc_hd__buf_6
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5786__A1 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3649__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7471_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4210__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3665__B _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7575_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold908 _4361_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold919 hold919/A VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3470_ _3469_/X _3470_/A1 _4429_/B VGND VGND VPWR VPWR _3470_/X sky130_fd_sc_hd__mux2_4
X_5140_ _4956_/A _4687_/Y _4761_/Y _4741_/Y _4706_/Y VGND VGND VPWR VPWR _5140_/X
+ sky130_fd_sc_hd__o32a_1
Xhold2309 _7092_/Q VGND VGND VPWR VPWR hold547/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_leaf_25_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6266__A2 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5071_ _5071_/A _5071_/B _5071_/C _4825_/A VGND VGND VPWR VPWR _5072_/D sky130_fd_sc_hd__nor4b_4
Xhold1608 _5905_/X VGND VGND VPWR VPWR hold276/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_193_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1619 _7482_/Q VGND VGND VPWR VPWR hold231/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2312_A _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4022_ _4014_/B _4017_/Y _4021_/X _4040_/D VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6671__C1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5226__B1 _5102_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5973_ _5973_/A0 hold17/X hold13/X VGND VGND VPWR VPWR _5973_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4924_ _5339_/A _4929_/A _5053_/C _5342_/B VGND VGND VPWR VPWR _4925_/C sky130_fd_sc_hd__nand4_2
XFILLER_0_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7643_ _7644_/CLK _7643_/D _4309_/B VGND VGND VPWR VPWR _7643_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4855_ _4644_/Y _4646_/Y _5222_/C _5404_/D _4966_/A VGND VGND VPWR VPWR _4855_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_118_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3806_ _7529_/Q _3529_/X _3670_/X _7134_/Q _3805_/X VGND VGND VPWR VPWR _3806_/X
+ sky130_fd_sc_hd__a221o_4
X_7574_ _7580_/CLK _7574_/D fanout597/X VGND VGND VPWR VPWR _7574_/Q sky130_fd_sc_hd__dfrtp_2
X_4786_ _4740_/D _4772_/A _4786_/C _4795_/C VGND VGND VPWR VPWR _4790_/C sky130_fd_sc_hd__and4bb_4
XFILLER_0_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6525_ _7498_/Q _6447_/C _6429_/X _6467_/X _7418_/Q VGND VGND VPWR VPWR _6525_/X
+ sky130_fd_sc_hd__a32o_1
X_3737_ _7522_/Q _5785_/B _5938_/C VGND VGND VPWR VPWR _3737_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6456_ _7487_/Q _6454_/X _6455_/X _7455_/Q _6453_/X VGND VGND VPWR VPWR _6456_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3668_ _4509_/A _4449_/B _4388_/B VGND VGND VPWR VPWR _4545_/A sky130_fd_sc_hd__and3_4
XFILLER_0_30_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5407_ _4887_/B _4945_/A _5399_/B _5404_/D VGND VGND VPWR VPWR _5410_/C sky130_fd_sc_hd__a31o_1
XANTENNA__5701__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6387_ _7146_/Q _6144_/C _6097_/B _6144_/B VGND VGND VPWR VPWR _6387_/X sky130_fd_sc_hd__o211a_1
X_3599_ _7317_/Q _5983_/A _5731_/B _3503_/X input32/X VGND VGND VPWR VPWR _3599_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout597_A fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5338_ _5203_/B _5329_/X _5337_/X VGND VGND VPWR VPWR _5340_/B sky130_fd_sc_hd__a21oi_1
Xhold2810 hold2810/A VGND VGND VPWR VPWR hold2810/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2821 _7031_/Q VGND VGND VPWR VPWR hold2821/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2832 _7041_/Q VGND VGND VPWR VPWR hold2832/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2843 _4182_/X VGND VGND VPWR VPWR hold2843/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4268__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5269_ _4698_/Y _5255_/X _5563_/A1 _5254_/X _5268_/X VGND VGND VPWR VPWR _5269_/X
+ sky130_fd_sc_hd__o311a_1
Xhold2854 _6947_/Q VGND VGND VPWR VPWR hold2854/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7008_ _7189_/CLK _7008_/D fanout572/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfstp_2
Xhold2865 hold2865/A VGND VGND VPWR VPWR _4492_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2876 _6980_/Q VGND VGND VPWR VPWR _4291_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold175_A _7246_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2887 _7488_/Q VGND VGND VPWR VPWR hold2887/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2898 hold2898/A VGND VGND VPWR VPWR _4252_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6407__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3491__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5768__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3779__B1 _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4440__A1 _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5965__B hold12/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6717__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3546__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5940__A1 _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input60_A mgmt_gpio_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6496__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__D _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6036__B _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6751__S _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5875__B _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3785__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4640_ _4733_/A _4733_/B _4641_/B VGND VGND VPWR VPWR _4778_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_21_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6184__A1 _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6184__B2 _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4571_ _4887_/B _4879_/C VGND VGND VPWR VPWR _4571_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6310_ _6963_/Q _6072_/B _6144_/B _6379_/B1 _7123_/Q VGND VGND VPWR VPWR _6310_/X
+ sky130_fd_sc_hd__a32o_1
Xmax_cap402 _4811_/A VGND VGND VPWR VPWR _5295_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3522_ hold27/A _5875_/A _5983_/A _3521_/X _7318_/Q VGND VGND VPWR VPWR _3522_/X
+ sky130_fd_sc_hd__a32o_1
Xhold705 _4529_/X VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7290_ _7501_/CLK _7290_/D fanout581/X VGND VGND VPWR VPWR _7290_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_123_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold716 hold716/A VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap424 _5216_/A VGND VGND VPWR VPWR _5553_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold727 _5754_/X VGND VGND VPWR VPWR _7363_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_97_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold738 hold738/A VGND VGND VPWR VPWR hold738/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold749 hold749/A VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6241_ _7293_/Q _6144_/A _6136_/C _6074_/X _7301_/Q VGND VGND VPWR VPWR _6241_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6487__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3453_ _3452_/X hold528/X _4429_/B VGND VGND VPWR VPWR _3453_/X sky130_fd_sc_hd__mux2_1
X_6172_ _7362_/Q _6332_/C _6379_/B1 _7394_/Q _6171_/X VGND VGND VPWR VPWR _6172_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2106 hold158/X VGND VGND VPWR VPWR _4502_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2117 _4222_/X VGND VGND VPWR VPWR hold800/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6239__A2 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5123_ _4605_/Y _4703_/Y _4826_/Y _4428_/B VGND VGND VPWR VPWR _5123_/X sky130_fd_sc_hd__o31a_1
Xhold2128 _4466_/X VGND VGND VPWR VPWR hold150/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2139 _7563_/Q VGND VGND VPWR VPWR hold145/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1405 hold1405/A VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1416 hold45/X VGND VGND VPWR VPWR _4179_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1427 hold221/X VGND VGND VPWR VPWR _5878_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1438 _7297_/Q VGND VGND VPWR VPWR hold191/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5054_ _5342_/A wire536/X _5260_/D _5058_/C _5180_/B VGND VGND VPWR VPWR _5056_/B
+ sky130_fd_sc_hd__a32oi_2
XANTENNA__5998__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1449 _5899_/X VGND VGND VPWR VPWR hold188/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4005_ _4005_/A _7071_/Q _4005_/C _7073_/Q VGND VGND VPWR VPWR _4006_/B sky130_fd_sc_hd__nor4_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4446__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5214__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6411__A2 _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5956_ _5965_/A _5956_/B hold48/X VGND VGND VPWR VPWR _5956_/X sky130_fd_sc_hd__and3_1
XANTENNA__4422__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5785__B _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4907_ _4933_/B _5213_/C _5260_/D VGND VGND VPWR VPWR _4907_/X sky130_fd_sc_hd__and3_1
XANTENNA__3776__A3 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4973__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5887_ hold213/X _5986_/A1 _5892_/S VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4181__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7626_ _7627_/CLK _7626_/D fanout569/X VGND VGND VPWR VPWR _7626_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6175__A1 _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4838_ _5058_/D _4856_/A _5282_/A _4839_/B VGND VGND VPWR VPWR _4841_/B sky130_fd_sc_hd__and4_1
XFILLER_0_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3528__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7557_ _7577_/CLK _7557_/D fanout584/X VGND VGND VPWR VPWR _7557_/Q sky130_fd_sc_hd__dfrtp_4
X_4769_ _5404_/C _5410_/B VGND VGND VPWR VPWR _4769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6508_ _7593_/Q _7577_/Q _6408_/C _6507_/X VGND VGND VPWR VPWR _6508_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_43_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7488_ _7560_/CLK _7488_/D fanout599/X VGND VGND VPWR VPWR _7488_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6478__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6439_ _7399_/Q _6409_/X _6437_/X _6438_/X VGND VGND VPWR VPWR _6439_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1627_A _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3700__A3 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__buf_4
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2640 hold637/X VGND VGND VPWR VPWR _5781_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2651 _7663_/A VGND VGND VPWR VPWR hold887/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2662 hold734/X VGND VGND VPWR VPWR _5934_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__buf_12
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__buf_2
XANTENNA__5989__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2673 _5880_/X VGND VGND VPWR VPWR hold743/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4864__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2684 hold893/X VGND VGND VPWR VPWR _4232_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2695 _7483_/Q VGND VGND VPWR VPWR hold781/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1950 hold476/X VGND VGND VPWR VPWR _4465_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1961 hold553/X VGND VGND VPWR VPWR _5752_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1972 _7029_/Q VGND VGND VPWR VPWR hold314/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1983 _7185_/Q VGND VGND VPWR VPWR hold434/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1994 hold478/X VGND VGND VPWR VPWR _4501_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_86_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6901__CLK _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4880__A _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5695__B _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3927__C _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6705__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5913__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_163_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_7 _3801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6469__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4758__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3662__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5429__B1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6641__A2 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_187_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5810_ _5810_/A0 _5954_/A1 _5811_/S VGND VGND VPWR VPWR _5810_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4790__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6790_ _3643_/Y _6790_/A1 _6792_/S VGND VGND VPWR VPWR _7634_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_119_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4404__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5741_ _5741_/A0 _5993_/A1 _5748_/S VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4955__A2 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5672_ _5951_/A1 _5672_/A1 _5676_/S VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__mux2_1
X_7411_ _7499_/CLK _7411_/D fanout578/X VGND VGND VPWR VPWR _7411_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4623_ _5127_/A _5222_/A _5107_/A VGND VGND VPWR VPWR _4841_/A sky130_fd_sc_hd__and3_1
XANTENNA__5825__S _5829_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3915__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7342_ _7555_/CLK _7342_/D fanout594/X VGND VGND VPWR VPWR _7342_/Q sky130_fd_sc_hd__dfrtp_4
X_4554_ _5914_/A1 _4554_/A1 _4556_/S VGND VGND VPWR VPWR _4554_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5380__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold502 hold502/A VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold513 _4306_/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold524 hold524/A VGND VGND VPWR VPWR hold524/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3505_ _3576_/B _3576_/C _3505_/C _3505_/D VGND VGND VPWR VPWR _3505_/Y sky130_fd_sc_hd__nor4_1
X_7273_ _7278_/CLK _7273_/D fanout580/X VGND VGND VPWR VPWR _7273_/Q sky130_fd_sc_hd__dfrtp_1
Xhold535 _5955_/X VGND VGND VPWR VPWR _7542_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold546 hold546/A VGND VGND VPWR VPWR _7226_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4485_ _4485_/A _5902_/B VGND VGND VPWR VPWR _4490_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2811_A _7287_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold557 hold557/A VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold568 hold568/A VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold579 hold579/A VGND VGND VPWR VPWR _7252_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2909_A _7399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6224_ _7468_/Q _6087_/X _6220_/X _6221_/X _6223_/X VGND VGND VPWR VPWR _6224_/X
+ sky130_fd_sc_hd__a2111o_2
X_3436_ _7354_/Q VGND VGND VPWR VPWR _3436_/Y sky130_fd_sc_hd__inv_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _7321_/Q _6116_/B _6081_/X _6075_/X _7425_/Q VGND VGND VPWR VPWR _6155_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3694__A2 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1202 hold1202/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5563_/A1 _4814_/Y _4844_/Y _5104_/Y VGND VGND VPWR VPWR _5111_/C sky130_fd_sc_hd__o31ai_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1213 hold2896/X VGND VGND VPWR VPWR hold1213/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _5714_/X VGND VGND VPWR VPWR _7327_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6086_ _7589_/Q _7588_/Q _6120_/B VGND VGND VPWR VPWR _6086_/X sky130_fd_sc_hd__and3_2
Xhold1235 _5993_/X VGND VGND VPWR VPWR _7575_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1246 hold3084/X VGND VGND VPWR VPWR hold3085/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1257 _5975_/X VGND VGND VPWR VPWR _7559_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5037_ _5037_/A _5037_/B _5037_/C VGND VGND VPWR VPWR _5039_/C sky130_fd_sc_hd__nand3_1
XANTENNA__6632__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1268 hold3098/X VGND VGND VPWR VPWR hold3099/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1279 _4504_/X VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_189_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6396__A1 _7025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6988_ _7409_/CLK _6988_/D fanout568/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6396__B2 _7201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5939_ _5939_/A0 _5993_/A1 hold23/X VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4850__D _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7609_ _7621_/CLK _7609_/D fanout575/X VGND VGND VPWR VPWR _7609_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6699__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5735__S _5739_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6420__A _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5371__A2 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1911_A _7231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input162_A wb_dat_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3482__C _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6320__A1 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5123__A2 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4564_/D sky130_fd_sc_hd__clkbuf_2
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _5071_/A sky130_fd_sc_hd__buf_12
Xhold3160 _7001_/Q VGND VGND VPWR VPWR hold3160/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3171 hold3171/A VGND VGND VPWR VPWR _4204_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3685__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6805_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3182 _7219_/Q VGND VGND VPWR VPWR _3645_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6812_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3193 _7616_/Q VGND VGND VPWR VPWR _6522_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6817_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6825_/A3 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2470 hold631/X VGND VGND VPWR VPWR _5670_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2481 _4261_/X VGND VGND VPWR VPWR hold659/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input23_A mask_rev_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6623__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2492 _7007_/Q VGND VGND VPWR VPWR hold696/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4634__A1 _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1780 _7098_/Q VGND VGND VPWR VPWR hold378/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1791 _7565_/Q VGND VGND VPWR VPWR hold1791/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6387__A1 _7146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4398__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__C _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6139__A1 _7400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6139__B2 _6116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5645__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5898__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5362__A2 _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3673__B _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A0 _5586_/A0 _4270_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5114__A2 _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3676__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4873__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2225_A _3564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6614__A2 _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6911_ _6926_/CLK _6911_/D fanout565/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6842_ _6873_/A _6869_/B VGND VGND VPWR VPWR _6842_/X sky130_fd_sc_hd__and2_1
XFILLER_0_77_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4389__A0 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6773_ _6773_/A _6773_/B _6773_/C _6773_/D VGND VGND VPWR VPWR _6774_/C sky130_fd_sc_hd__nor4_2
X_3985_ _7648_/A _3933_/A _5612_/B _3984_/X VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5724_ hold586/X _5967_/A1 _5730_/S VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3600__A2 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5655_ hold84/X _5655_/A1 _5656_/S VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3864__A hold36/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7157__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4606_ _4887_/D _4747_/B VGND VGND VPWR VPWR _5387_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5353__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5586_ _5586_/A0 _5586_/A1 _5586_/S VGND VGND VPWR VPWR _5586_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6550__A1 _7451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold310 hold310/A VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7325_ _7429_/CLK _7325_/D fanout583/X VGND VGND VPWR VPWR _7325_/Q sky130_fd_sc_hd__dfrtp_4
Xhold321 hold321/A VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4537_ _5852_/A0 _4537_/A1 _4538_/S VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__mux2_1
Xhold332 hold332/A VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold343 hold343/A VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_159_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold354 hold354/A VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7256_ _7266_/CLK _7256_/D fanout567/X VGND VGND VPWR VPWR _7256_/Q sky130_fd_sc_hd__dfrtp_4
Xhold365 hold365/A VGND VGND VPWR VPWR _7554_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold376 hold376/A VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4468_ _5840_/A1 _4468_/A1 _4472_/S VGND VGND VPWR VPWR _4468_/X sky130_fd_sc_hd__mux2_1
Xhold387 hold387/A VGND VGND VPWR VPWR _7570_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold398 _3456_/X VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_110_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6207_ _6204_/X _6205_/X _6206_/X _6116_/B VGND VGND VPWR VPWR _6207_/X sky130_fd_sc_hd__o31a_1
X_3419_ _7490_/Q VGND VGND VPWR VPWR _3419_/Y sky130_fd_sc_hd__inv_2
X_7187_ _7268_/CLK _7187_/D _6871_/A VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfrtp_4
X_4399_ _5754_/A1 _4399_/A1 _4399_/S VGND VGND VPWR VPWR _4399_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_73_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _7368_/Q _6084_/X _6136_/X _6137_/X _6135_/X VGND VGND VPWR VPWR _6138_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold1010 hold2756/X VGND VGND VPWR VPWR hold2757/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1021 hold2884/X VGND VGND VPWR VPWR hold2885/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _5976_/X VGND VGND VPWR VPWR _7560_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6605__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1043 hold2887/X VGND VGND VPWR VPWR hold2888/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6649_/S _4117_/B _6067_/X VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__a21o_1
Xhold1054 hold2776/X VGND VGND VPWR VPWR _7172_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 _4359_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 hold2813/X VGND VGND VPWR VPWR hold2814/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _4498_/X VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1098 hold2874/X VGND VGND VPWR VPWR hold2875/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6415__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6369__B2 _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4580__D _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6384__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6541__A1 _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6541__B2 _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4552__A0 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__B _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4607__A1 _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6028__C _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3830__A2 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3668__B _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6044__B _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3770_ _7029_/Q _3669_/C _5632_/B _3649_/X _7069_/Q VGND VGND VPWR VPWR _3770_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5440_ _5199_/C _5058_/C _5439_/X VGND VGND VPWR VPWR _5506_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__6532__A1 _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6532__B2 _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5371_ _5059_/B _5404_/D _4966_/A _5248_/A VGND VGND VPWR VPWR _5371_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_22_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7110_ _7644_/CLK _7110_/D _4309_/B VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfrtp_4
X_4322_ _4322_/A _5902_/B VGND VGND VPWR VPWR _4327_/S sky130_fd_sc_hd__nand2_4
XANTENNA__5107__C _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7041_ _7201_/CLK _7041_/D _6839_/A VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_4
X_4253_ _4253_/A0 _5986_/A1 _4258_/S VGND VGND VPWR VPWR _4253_/X sky130_fd_sc_hd__mux2_1
X_4184_ _4184_/A0 _5583_/A0 _4190_/S VGND VGND VPWR VPWR _4184_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3821__A2 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_6825_ _7110_/Q _6824_/C _6825_/A3 _6824_/X VGND VGND VPWR VPWR _6825_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3968_ _7279_/Q _3558_/X _4394_/A _7061_/Q _3967_/X VGND VGND VPWR VPWR _3968_/X
+ sky130_fd_sc_hd__a221o_1
X_6756_ _7065_/Q _6574_/B _6441_/X _6419_/D _7005_/Q VGND VGND VPWR VPWR _6756_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6771__B2 _7141_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5707_ _5896_/A0 _5707_/A1 _5712_/S VGND VGND VPWR VPWR _5707_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6687_ _6968_/Q _6420_/A _6457_/X _7062_/Q _6686_/X VGND VGND VPWR VPWR _6687_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_61_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3899_ _7488_/Q _3569_/X _5581_/A _7210_/Q _3898_/X VGND VGND VPWR VPWR _3899_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5638_ _5996_/A1 _5638_/A1 _5639_/S VGND VGND VPWR VPWR _5638_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4534__A0 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5569_ _5569_/A _5569_/B _5569_/C VGND VGND VPWR VPWR _5569_/X sky130_fd_sc_hd__and3_1
XANTENNA__3888__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold140 hold140/A VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7308_ _7542_/CLK _7308_/D fanout581/X VGND VGND VPWR VPWR _7308_/Q sky130_fd_sc_hd__dfrtp_4
Xhold151 hold151/A VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold162 hold162/A VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold173 hold173/A VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6287__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold184 hold184/A VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold195 hold195/A VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7239_ _7239_/CLK _7239_/D fanout566/X VGND VGND VPWR VPWR _7239_/Q sky130_fd_sc_hd__dfstp_1
Xfanout620 _4887_/D VGND VGND VPWR VPWR _4743_/A sky130_fd_sc_hd__buf_8
XANTENNA__4575__D _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A wb_adr_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__B _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5262__A1 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5262__B2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3488__B _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7079__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6762__B2 _7146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input90_A spimemio_flash_io2_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6514__A1 _7441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__1111_ clkbuf_0__1111_/X VGND VGND VPWR VPWR _6789_/A2 sky130_fd_sc_hd__clkbuf_16
XANTENNA__6278__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3670__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5253__A1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4940_ _4954_/A _5453_/A _4940_/C _4940_/D VGND VGND VPWR VPWR _4941_/B sky130_fd_sc_hd__and4_1
XANTENNA__3803__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4871_ _4747_/B _4879_/C _4887_/B _4887_/D VGND VGND VPWR VPWR _4937_/C sky130_fd_sc_hd__and4bb_4
XFILLER_0_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6610_ _7365_/Q _6462_/X _6607_/X _6609_/X VGND VGND VPWR VPWR _6610_/X sky130_fd_sc_hd__a211o_1
X_3822_ _7159_/Q hold56/A _5632_/B _3647_/X _7169_/Q VGND VGND VPWR VPWR _3822_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_21_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7590_ _7593_/CLK _7590_/D fanout567/X VGND VGND VPWR VPWR _7590_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3567__A1 _7334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6541_ _7394_/Q _6420_/C _6421_/X _7322_/Q _6540_/X VGND VGND VPWR VPWR _6544_/C
+ sky130_fd_sc_hd__a221o_1
X_3753_ input95/X _5785_/B _5659_/B _3526_/X _7506_/Q VGND VGND VPWR VPWR _3753_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_171_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4303__A _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6472_ wire348/X _6471_/Y _7279_/Q _6431_/Y VGND VGND VPWR VPWR _6472_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3684_ _7283_/Q _3590_/C _5659_/B _5848_/A _7451_/Q VGND VGND VPWR VPWR _3684_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5423_ _5423_/A _5423_/B VGND VGND VPWR VPWR _5438_/C sky130_fd_sc_hd__and2_1
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 _3412_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
XFILLER_0_112_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5833__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput212 _3436_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
Xoutput223 _7660_/X VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
Xoutput234 _4146_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
X_5354_ _5213_/B _5077_/B _5248_/C _5213_/X _5350_/X VGND VGND VPWR VPWR _5355_/D
+ sky130_fd_sc_hd__a311oi_4
Xoutput245 _4151_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
XFILLER_0_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput256 _7233_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
Xoutput267 _7230_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
XANTENNA__6269__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4305_ _4305_/A0 _5805_/A1 _4308_/S VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3861__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput278 _7237_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
Xoutput289 _6923_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
X_5285_ _5395_/A1 _5059_/B _5118_/B _5284_/X VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__a31o_1
X_7024_ _7024_/CLK _7024_/D fanout568/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_4
X_4236_ _5652_/A1 _5967_/A1 _4248_/S VGND VGND VPWR VPWR _4236_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4295__A2 _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4167_ _7601_/Q _7251_/Q _7255_/Q VGND VGND VPWR VPWR _4167_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_A _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4098_ _4098_/A1 _4011_/X _4123_/C _7071_/Q _4010_/Y VGND VGND VPWR VPWR _7071_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4692__B _4758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7170_/CLK sky130_fd_sc_hd__clkbuf_16
X_6808_ _7111_/Q _6808_/A2 _6808_/B1 _7110_/Q VGND VGND VPWR VPWR _6808_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6744__A1 _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6744__B2 _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6739_ _7145_/Q _6468_/X _6734_/X _6736_/X _6738_/X VGND VGND VPWR VPWR _6749_/A
+ sky130_fd_sc_hd__a2111o_2
XANTENNA__6412__B _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5743__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3730__B2 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3490__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout472 _4256_/A1 VGND VGND VPWR VPWR _5863_/A0 sky130_fd_sc_hd__clkbuf_16
XANTENNA__6680__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout483 _5735_/A1 VGND VGND VPWR VPWR _5852_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4883__A _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout494 hold1724/X VGND VGND VPWR VPWR hold1725/A sky130_fd_sc_hd__buf_6
XANTENNA__6432__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4107__B _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3665__C _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6499__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold909 hold909/A VGND VGND VPWR VPWR hold909/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5171__B1 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3721__A1 input16/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5070_ _4706_/A _5072_/C _4940_/C _5134_/A VGND VGND VPWR VPWR _5070_/X sky130_fd_sc_hd__a22o_1
Xhold1609 _7382_/Q VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4021_ _6905_/Q _6904_/Q _4025_/B hold51/A VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_79_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5972_ _5972_/A0 _5999_/A1 hold13/X VGND VGND VPWR VPWR _5972_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_176_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4923_ _5453_/A _4954_/C _4929_/A _4937_/C VGND VGND VPWR VPWR _5444_/C sky130_fd_sc_hd__nand4_1
XFILLER_0_74_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5828__S _5829_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2674_A _7467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7642_ _7646_/CLK _7642_/D _4309_/B VGND VGND VPWR VPWR _7642_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4854_ _4622_/Y _4654_/Y _4748_/Y _7111_/Q VGND VGND VPWR VPWR _4854_/X sky130_fd_sc_hd__o31a_2
XFILLER_0_16_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3856__B _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3805_ input97/X _5785_/B _5659_/B _5634_/A _7258_/Q VGND VGND VPWR VPWR _3805_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_172_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7573_ _7580_/CLK _7573_/D fanout597/X VGND VGND VPWR VPWR _7573_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4785_ _4700_/Y _4707_/Y _4784_/Y _4781_/Y VGND VGND VPWR VPWR _4791_/B sky130_fd_sc_hd__o211ai_1
XANTENNA_hold2841_A _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2939_A _7648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3736_ _7218_/Q _3996_/A _3734_/Y _3735_/X VGND VGND VPWR VPWR _7218_/D sky130_fd_sc_hd__a22o_2
X_6524_ _7530_/Q _6058_/X _6409_/X _7402_/Q VGND VGND VPWR VPWR _6524_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3960__A1 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3667_ _5640_/B _5612_/C _4346_/C VGND VGND VPWR VPWR _3667_/X sky130_fd_sc_hd__and3_4
X_6455_ _6463_/A _6455_/B _6600_/B VGND VGND VPWR VPWR _6455_/X sky130_fd_sc_hd__and3_4
XFILLER_0_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5406_ _4879_/C _5011_/B _5113_/A VGND VGND VPWR VPWR _5406_/Y sky130_fd_sc_hd__a21oi_2
X_6386_ _6878_/Q _6112_/X _6121_/X _6992_/Q VGND VGND VPWR VPWR _6386_/X sky130_fd_sc_hd__a22o_1
X_3598_ _5590_/A _5612_/B _3931_/D VGND VGND VPWR VPWR _3598_/X sky130_fd_sc_hd__and3_1
XFILLER_0_140_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3712__A1 _7515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5337_ _5038_/B _5053_/C _5328_/X _5336_/X VGND VGND VPWR VPWR _5337_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4179__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2800 _6981_/Q VGND VGND VPWR VPWR _4293_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2811 _7287_/Q VGND VGND VPWR VPWR hold2811/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5268_ _5255_/X _4774_/Y _5267_/X _5266_/Y VGND VGND VPWR VPWR _5268_/X sky130_fd_sc_hd__o211a_1
Xhold2822 hold2822/A VGND VGND VPWR VPWR _4359_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2833 hold2833/A VGND VGND VPWR VPWR _4371_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5465__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2844 _7651_/A VGND VGND VPWR VPWR hold594/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2855 hold2855/A VGND VGND VPWR VPWR _4247_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7007_ _7191_/CLK _7007_/D fanout572/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_4
X_4219_ _4252_/A0 _5985_/A1 _4231_/S VGND VGND VPWR VPWR _4219_/X sky130_fd_sc_hd__mux2_1
Xhold2866 _7152_/Q VGND VGND VPWR VPWR hold2866/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2877 hold2877/A VGND VGND VPWR VPWR hold2877/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5199_ _5282_/A _5342_/A _5199_/C _5342_/C VGND VGND VPWR VPWR _5200_/B sky130_fd_sc_hd__nand4b_2
Xhold2888 hold2888/A VGND VGND VPWR VPWR _5895_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2899 _4252_/X VGND VGND VPWR VPWR hold2899/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_97_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6407__B _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3779__B2 _7145_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5738__S _5739_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4440__A2 hold284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5965__C hold48/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_176_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6423__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6717__B2 _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3951__A1 _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3951__B2 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3155_A _6988_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4597__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input53_A mgmt_gpio_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3703__B2 _7116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6248__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6653__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7094__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6317__B _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5208__A1 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output307_A _4134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6036__C _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5648__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5875__C _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6184__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4195__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4570_ _4795_/C _4772_/A _4805_/B VGND VGND VPWR VPWR _4570_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_181_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3521_ _5590_/A _4449_/B _5731_/B VGND VGND VPWR VPWR _3521_/X sky130_fd_sc_hd__and3_4
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3942__A1 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold706 hold706/A VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold717 _5718_/X VGND VGND VPWR VPWR _7331_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold728 hold728/A VGND VGND VPWR VPWR hold728/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6240_ _7333_/Q _6136_/B _6116_/A _6112_/C VGND VGND VPWR VPWR _6240_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold739 hold739/A VGND VGND VPWR VPWR _7228_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3452_ _4028_/A0 _4025_/A hold51/X VGND VGND VPWR VPWR _3452_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6171_ _7298_/Q _6136_/B _6144_/B _6079_/X _7330_/Q VGND VGND VPWR VPWR _6171_/X
+ sky130_fd_sc_hd__a32o_1
X_5122_ _5061_/X _5122_/B _5122_/C VGND VGND VPWR VPWR _5122_/Y sky130_fd_sc_hd__nand3b_1
Xhold2107 _4502_/X VGND VGND VPWR VPWR hold159/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2118 _7093_/Q VGND VGND VPWR VPWR hold2118/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2129 hold150/X VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1406 _6884_/Q VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6644__B1 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5053_ _5339_/D _5342_/A _5053_/C VGND VGND VPWR VPWR _5058_/C sky130_fd_sc_hd__and3_4
Xhold1417 _4179_/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1428 _5878_/X VGND VGND VPWR VPWR hold222/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1439 hold191/X VGND VGND VPWR VPWR _5680_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4004_ _4004_/A _4006_/A VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__xor2_1
XANTENNA__4670__A2 _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2889_A _7260_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5955_ _5955_/A0 _5955_/A1 _5955_/S VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4970__B _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4906_ _4906_/A _4906_/B _5185_/C _4906_/D VGND VGND VPWR VPWR _4906_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3630__B1 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5886_ _5886_/A0 _5985_/A1 _5892_/S VGND VGND VPWR VPWR _7480_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_158_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7625_ _7627_/CLK _7625_/D fanout566/X VGND VGND VPWR VPWR _7625_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4837_ _4837_/A _4837_/B _4837_/C VGND VGND VPWR VPWR _4841_/C sky130_fd_sc_hd__nand3_1
XANTENNA__6175__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4186__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7556_ _7556_/CLK _7556_/D fanout597/X VGND VGND VPWR VPWR _7556_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout505_A hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4768_ _4740_/D _4768_/B VGND VGND VPWR VPWR _4768_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_71_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6507_ _7433_/Q _6747_/B _6747_/C _6408_/A _7553_/Q VGND VGND VPWR VPWR _6507_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3719_ _7146_/Q _5803_/A _5938_/B _4551_/C _3718_/X VGND VGND VPWR VPWR _3719_/X
+ sky130_fd_sc_hd__a41o_1
X_4699_ _4743_/A _4856_/A _4888_/B VGND VGND VPWR VPWR _5282_/B sky130_fd_sc_hd__nor3_4
X_7487_ _7487_/CLK _7487_/D fanout597/X VGND VGND VPWR VPWR _7487_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_141_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6438_ _7391_/Q _6420_/C _6419_/A _7543_/Q VGND VGND VPWR VPWR _6438_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_140_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6369_ _7004_/Q _6097_/B _6120_/B _6379_/B1 _7125_/Q VGND VGND VPWR VPWR _6369_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_22_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7415_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2630 _7254_/Q VGND VGND VPWR VPWR hold866/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6635__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__clkbuf_2
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2641 _7379_/Q VGND VGND VPWR VPWR hold710/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2652 hold887/X VGND VGND VPWR VPWR _4423_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__buf_4
Xhold2663 _7403_/Q VGND VGND VPWR VPWR hold728/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2674 _7467_/Q VGND VGND VPWR VPWR hold740/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1940 _5798_/X VGND VGND VPWR VPWR hold361/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2685 _4232_/X VGND VGND VPWR VPWR hold894/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4110__A1 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1951 _4465_/X VGND VGND VPWR VPWR hold477/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2696 hold781/X VGND VGND VPWR VPWR _5889_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1962 _5752_/X VGND VGND VPWR VPWR hold554/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1973 hold314/X VGND VGND VPWR VPWR _4356_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_37_csclk _7267_/CLK VGND VGND VPWR VPWR _7578_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4661__A2 _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1984 hold434/X VGND VGND VPWR VPWR _4537_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1995 _4501_/X VGND VGND VPWR VPWR hold479/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_39_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5610__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5695__C _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3621__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3927__D _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6166__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_68_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5992__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6600__B _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 _3894_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6469__A3 _6429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5216__B _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output257_A _7234_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5429__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6626__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7204__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6047__B _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5601__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5740_ _5785_/A _5884_/B _5992_/D VGND VGND VPWR VPWR _5748_/S sky130_fd_sc_hd__and3_4
XANTENNA__3612__B1 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4955__A3 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5671_ _5896_/A0 hold197/X _5676_/S VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7410_ _7412_/CLK _7410_/D fanout581/X VGND VGND VPWR VPWR _7410_/Q sky130_fd_sc_hd__dfrtp_4
X_4622_ _4947_/C _4657_/A VGND VGND VPWR VPWR _4622_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_25_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4553_ _5940_/A1 _4553_/A1 _4556_/S VGND VGND VPWR VPWR _4553_/X sky130_fd_sc_hd__mux2_1
X_7341_ _7478_/CLK _7341_/D fanout580/X VGND VGND VPWR VPWR _7341_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5380__A3 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold503 hold503/A VGND VGND VPWR VPWR _7462_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold514 hold514/A VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold525 hold525/A VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3504_ _3505_/C hold34/X VGND VGND VPWR VPWR _3504_/Y sky130_fd_sc_hd__nor2_4
X_4484_ _4484_/A0 _5586_/A0 _4484_/S VGND VGND VPWR VPWR _4484_/X sky130_fd_sc_hd__mux2_1
Xhold536 hold536/A VGND VGND VPWR VPWR hold536/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7272_ _7278_/CLK _7272_/D fanout580/X VGND VGND VPWR VPWR _7272_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6314__C1 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold547 hold547/A VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4668__D _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold558 hold558/A VGND VGND VPWR VPWR _7454_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold569 hold569/A VGND VGND VPWR VPWR _7472_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6223_ _7532_/Q _6092_/X _6112_/X _7484_/Q _6222_/X VGND VGND VPWR VPWR _6223_/X
+ sky130_fd_sc_hd__a221o_1
X_3435_ _7362_/Q VGND VGND VPWR VPWR _3435_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _7353_/Q _6099_/X _6110_/X _7433_/Q _6153_/X VGND VGND VPWR VPWR _6157_/B
+ sky130_fd_sc_hd__a221oi_2
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6617__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3694__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 hold2853/X VGND VGND VPWR VPWR hold1203/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5105_ _5387_/C _5399_/C _5453_/C VGND VGND VPWR VPWR _5105_/X sky130_fd_sc_hd__and3_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6119_/B _6121_/A _6332_/B _6112_/D VGND VGND VPWR VPWR _6085_/X sky130_fd_sc_hd__and4b_4
Xhold1214 hold1214/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xhold1225 hold3067/X VGND VGND VPWR VPWR hold3068/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1236 hold3074/X VGND VGND VPWR VPWR hold3075/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5036_ _4821_/Y _4862_/X _4865_/Y _4992_/Y _5035_/Y VGND VGND VPWR VPWR _5037_/A
+ sky130_fd_sc_hd__o311a_1
Xhold1247 _5984_/X VGND VGND VPWR VPWR _7567_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1258 hold3116/X VGND VGND VPWR VPWR hold3117/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1269 _4329_/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5840__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6987_ _7206_/CLK _6987_/D VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6396__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3603__B1 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5938_ hold22/X _5938_/B _5938_/C _5992_/D VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__and4_1
XFILLER_0_180_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5869_ _5869_/A0 _5986_/A1 _5874_/S VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7608_ _7621_/CLK _7608_/D fanout579/X VGND VGND VPWR VPWR _7608_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3906__A1 input15/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7539_ _7539_/CLK hold93/X fanout578/X VGND VGND VPWR VPWR _7539_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3906__B2 _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6420__B _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6320__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4331__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input155_A wb_dat_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4875__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4564_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3150 _7187_/Q VGND VGND VPWR VPWR hold3150/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _4825_/A sky130_fd_sc_hd__buf_12
Xhold3161 hold3161/A VGND VGND VPWR VPWR _4323_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6608__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3172 _7407_/Q VGND VGND VPWR VPWR hold3172/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3685__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6808_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3183 _3645_/X VGND VGND VPWR VPWR _7219_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6814_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3194 _6498_/X VGND VGND VPWR VPWR _7616_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2460 hold656/X VGND VGND VPWR VPWR _4214_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6820_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6795_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2471 _6920_/Q VGND VGND VPWR VPWR hold664/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2482 _7225_/Q VGND VGND VPWR VPWR hold678/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2493 hold696/X VGND VGND VPWR VPWR _4330_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1770 _4396_/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5292__C1 _4428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5831__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4634__A2 _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input16_A mask_rev_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1781 hold378/X VGND VGND VPWR VPWR _4446_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1792 hold1792/A VGND VGND VPWR VPWR _5981_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6387__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6139__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4131__A _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3673__C _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6311__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4428__A_N _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3676__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6614__A3 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5822__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6910_ _7075_/CLK _6910_/D _6860_/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3833__B1 _3675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6841_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6841_/X sky130_fd_sc_hd__and2_1
XANTENNA__5586__A0 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6772_ _6971_/Q _6420_/A _6422_/X _6966_/Q _6771_/X VGND VGND VPWR VPWR _6773_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3984_ input4/X _3503_/X _3675_/X _7187_/Q VGND VGND VPWR VPWR _3984_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5723_ _5723_/A0 _5903_/A0 _5730_/S VGND VGND VPWR VPWR _5723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5836__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5654_ _5951_/A1 _5654_/A1 _5656_/S VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5889__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3864__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4605_ _5260_/A _5260_/B VGND VGND VPWR VPWR _4605_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5353__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5585_ _5951_/A1 _5585_/A1 _5586_/S VGND VGND VPWR VPWR _5585_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6550__A2 _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_170_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold300 hold300/A VGND VGND VPWR VPWR hold300/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold311 hold311/A VGND VGND VPWR VPWR _7449_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7324_ _7412_/CLK _7324_/D fanout580/X VGND VGND VPWR VPWR _7324_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4536_ _5914_/A1 _4536_/A1 _4538_/S VGND VGND VPWR VPWR _4536_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold322 hold322/A VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold333 hold333/A VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold344 hold344/A VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold355 hold355/A VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7255_ _7255_/CLK _7255_/D fanout569/X VGND VGND VPWR VPWR _7255_/Q sky130_fd_sc_hd__dfrtp_4
Xhold366 hold366/A VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6302__A2 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4467_ _4467_/A _4551_/D VGND VGND VPWR VPWR _4472_/S sky130_fd_sc_hd__nand2_4
Xhold377 hold377/A VGND VGND VPWR VPWR _7175_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold388 hold388/A VGND VGND VPWR VPWR hold388/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold399 _3457_/X VGND VGND VPWR VPWR _3557_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6206_ _7299_/Q _6022_/X _6035_/Y _6073_/X _7387_/Q VGND VGND VPWR VPWR _6206_/X
+ sky130_fd_sc_hd__a32o_1
X_3418_ _7498_/Q VGND VGND VPWR VPWR _3418_/Y sky130_fd_sc_hd__inv_2
X_4398_ _5647_/A0 _4398_/A1 _4399_/S VGND VGND VPWR VPWR _4398_/X sky130_fd_sc_hd__mux2_1
X_7186_ _7186_/CLK _7186_/D fanout589/X VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4187__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A mask_rev_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 hold2405/X VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6137_ _7288_/Q _6144_/A _6136_/C _6079_/X _7328_/Q VGND VGND VPWR VPWR _6137_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _5678_/X VGND VGND VPWR VPWR _7295_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 hold2886/X VGND VGND VPWR VPWR _7464_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1033 hold2904/X VGND VGND VPWR VPWR hold2905/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6605__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1044 _5895_/X VGND VGND VPWR VPWR _7488_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6751_/S _4117_/B _6067_/X VGND VGND VPWR VPWR _6573_/S sky130_fd_sc_hd__a21oi_4
XFILLER_0_175_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1055 hold2772/X VGND VGND VPWR VPWR hold2773/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 hold2811/X VGND VGND VPWR VPWR hold2812/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5813__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 _4456_/X VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5019_ _5024_/A1 _4669_/X _4974_/B _5180_/A _5158_/A VGND VGND VPWR VPWR _5021_/C
+ sky130_fd_sc_hd__o2111ai_1
Xhold1088 hold2929/X VGND VGND VPWR VPWR hold2930/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 _4468_/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6415__B _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6369__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5746__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6541__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__C _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4886__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4304__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4607__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5804__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2290 _5820_/X VGND VGND VPWR VPWR hold601/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3830__A3 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4126__A _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3668__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3594__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6532__A2 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4543__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5370_ _4659_/Y _4844_/Y _5457_/B _5512_/A _5367_/Y VGND VGND VPWR VPWR _5370_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4321_ _3570_/Y _4321_/A1 _4321_/S VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7040_ _7189_/CLK _7040_/D fanout572/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfrtp_4
X_4252_ _4252_/A0 _5985_/A1 _4258_/S VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4183_ _4183_/A0 _7638_/Q _4429_/B VGND VGND VPWR VPWR _4183_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5256__C1 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6599__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3859__B hold36/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3821__A3 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6824_ _7111_/Q _6824_/B _6824_/C VGND VGND VPWR VPWR _6824_/X sky130_fd_sc_hd__and3_1
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6755_ _7166_/Q _6463_/X _6466_/X _7213_/Q _6754_/X VGND VGND VPWR VPWR _6755_/X
+ sky130_fd_sc_hd__a221o_1
X_3967_ _7051_/Q _4509_/A _5619_/B _3966_/X VGND VGND VPWR VPWR _3967_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_57_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6771__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5706_ _5967_/A1 _5706_/A1 _5712_/S VGND VGND VPWR VPWR _5706_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3585__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6686_ _7173_/Q _6747_/B _6747_/C _6425_/X _7017_/Q VGND VGND VPWR VPWR _6686_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout418_A hold21/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3898_ _7173_/Q _5866_/B _4521_/B _3647_/X _7168_/Q VGND VGND VPWR VPWR _3898_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5637_ _5985_/A1 _5637_/A1 _5639_/S VGND VGND VPWR VPWR _5637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5568_ _5568_/A _5568_/B _5568_/C VGND VGND VPWR VPWR _5569_/C sky130_fd_sc_hd__and3_1
XFILLER_0_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold130 hold130/A VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__clkbuf_2
Xhold141 hold141/A VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7307_ _7359_/CLK hold89/X fanout576/X VGND VGND VPWR VPWR _7307_/Q sky130_fd_sc_hd__dfrtp_4
X_4519_ _4519_/A0 _5647_/A0 _4520_/S VGND VGND VPWR VPWR _4519_/X sky130_fd_sc_hd__mux2_1
Xhold152 hold152/A VGND VGND VPWR VPWR _7275_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold163 _5916_/X VGND VGND VPWR VPWR _7507_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5499_ _5499_/A _5499_/B _5433_/C VGND VGND VPWR VPWR _5572_/A sky130_fd_sc_hd__nor3b_1
Xhold174 hold174/A VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold185 hold185/A VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6287__B2 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7238_ _7239_/CLK _7238_/D fanout566/X VGND VGND VPWR VPWR _7238_/Q sky130_fd_sc_hd__dfstp_2
Xfanout610 _4831_/A VGND VGND VPWR VPWR _4795_/C sky130_fd_sc_hd__buf_12
Xhold196 hold196/A VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout621 input110/X VGND VGND VPWR VPWR _4887_/D sky130_fd_sc_hd__buf_12
XANTENNA__5495__C1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7169_ _7170_/CLK _7169_/D fanout573/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6039__A1 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1602_A _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5798__A0 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A wb_adr_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4470__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3488__C _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6762__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input83_A spimemio_flash_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6514__A2 _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4525__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4289__A0 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6450__A1 _7559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3803__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4870_ _4947_/C _5213_/B _5213_/C VGND VGND VPWR VPWR _4877_/A sky130_fd_sc_hd__and3_4
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3821_ _7028_/Q _3669_/C _5603_/B _5848_/A _7449_/Q VGND VGND VPWR VPWR _3828_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_156_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6753__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3567__A2 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6540_ _7378_/Q _6408_/B _6460_/X _7386_/Q VGND VGND VPWR VPWR _6540_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_144_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3752_ _7530_/Q _3529_/X _3535_/X _7482_/Q _3751_/X VGND VGND VPWR VPWR _3759_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6471_ _6471_/A _6471_/B _6471_/C _6471_/D VGND VGND VPWR VPWR _6471_/Y sky130_fd_sc_hd__nor4_2
X_3683_ _7228_/Q hold12/A _5640_/C _5630_/S _7250_/Q VGND VGND VPWR VPWR _3683_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__4303__B _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6505__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2452_A _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4516__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5422_ _5422_/A _5422_/B _5496_/A _5422_/D VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__and4_1
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput202 _3411_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
XFILLER_0_23_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput213 _4156_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
Xoutput224 _7661_/X VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
Xoutput235 _4147_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
X_5353_ _4622_/Y _4726_/Y _4946_/Y _4898_/Y _5352_/Y VGND VGND VPWR VPWR _5355_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput246 _4128_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput257 _7234_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
X_4304_ _4304_/A0 _5948_/A1 _4308_/S VGND VGND VPWR VPWR _4304_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3861__C _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput268 _7231_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
XANTENNA__6269__B2 _7310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput279 _7238_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
X_5284_ _5399_/B _5081_/A _5115_/X _5281_/X VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__a31o_1
X_7023_ _7024_/CLK _7023_/D fanout568/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfstp_2
X_4235_ _4235_/A0 _4234_/X _4249_/S VGND VGND VPWR VPWR _4235_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4166_ _7599_/Q _7252_/Q _7255_/Q VGND VGND VPWR VPWR _4166_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4097_ _4171_/B _4084_/X _4096_/X _4114_/B VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__a22o_1
XANTENNA_fanout368_A _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4692__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout535_A _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6807_ _6806_/X _6807_/A1 _6822_/S VGND VGND VPWR VPWR _7639_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4999_ _5183_/A _5203_/B _5018_/B VGND VGND VPWR VPWR _5026_/A sky130_fd_sc_hd__and3_1
XANTENNA__6744__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6738_ _7019_/Q _6425_/X _6457_/X _7064_/Q _6737_/X VGND VGND VPWR VPWR _6738_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6412__C _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6669_ _7122_/Q _6420_/C _6467_/X _7152_/Q _6668_/X VGND VGND VPWR VPWR _6669_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1552_A _7508_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4507__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5028__C _5028_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3730__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout440 _6056_/X VGND VGND VPWR VPWR _6447_/C sky130_fd_sc_hd__buf_8
XANTENNA__5483__A2 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout473 _4256_/A1 VGND VGND VPWR VPWR _5998_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout484 _5995_/A1 VGND VGND VPWR VPWR _5950_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout495 _5714_/A0 VGND VGND VPWR VPWR _5948_/A1 sky130_fd_sc_hd__buf_12
XFILLER_0_69_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6432__A1 _7527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5171__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3721__A2 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2033_A _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4020_ _4019_/X _4018_/X _4040_/A _3450_/B VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5971_ _5971_/A0 _5998_/A1 hold13/X VGND VGND VPWR VPWR _5971_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4922_ _4922_/A _4922_/B _4922_/C VGND VGND VPWR VPWR _4925_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7641_ _7646_/CLK _7641_/D _4309_/B VGND VGND VPWR VPWR _7641_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6187__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4853_ _5248_/A _5094_/A VGND VGND VPWR VPWR _4853_/Y sky130_fd_sc_hd__nand2_1
X_3804_ _7521_/Q _5929_/A _5776_/A _7385_/Q _3803_/X VGND VGND VPWR VPWR _3804_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5934__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7572_ _7572_/CLK _7572_/D fanout596/X VGND VGND VPWR VPWR _7572_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4784_ _5113_/A _4784_/B VGND VGND VPWR VPWR _4784_/Y sky130_fd_sc_hd__nand2_1
X_6523_ _6522_/X _6523_/A1 _6573_/S VGND VGND VPWR VPWR _7617_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3735_ _3797_/A1 _3856_/A _7073_/Q _6893_/Q VGND VGND VPWR VPWR _3735_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6454_ _7595_/Q _6463_/A _6600_/B _7596_/Q VGND VGND VPWR VPWR _6454_/X sky130_fd_sc_hd__and4b_4
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmgmt_gpio_31_buff_inst _4163_/X VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3666_ hold36/A _5612_/C _4346_/C VGND VGND VPWR VPWR _3666_/X sky130_fd_sc_hd__and3_4
X_5405_ _4756_/X _5134_/X _5405_/C _5405_/D VGND VGND VPWR VPWR _5538_/B sky130_fd_sc_hd__and4bb_1
XANTENNA__5162__A1 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6385_ _7065_/Q _6032_/Y _6081_/X _7196_/Q _6384_/X VGND VGND VPWR VPWR _6385_/X
+ sky130_fd_sc_hd__a221o_1
X_3597_ hold76/A _5983_/A _5938_/C _3535_/X _7485_/Q VGND VGND VPWR VPWR _3597_/X
+ sky130_fd_sc_hd__a32o_4
X_5336_ _4996_/A _5038_/B _5328_/X _5335_/X VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3712__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2801 hold2801/A VGND VGND VPWR VPWR hold2801/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2812 hold2812/A VGND VGND VPWR VPWR _5669_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5267_ _4803_/A _4775_/C _4946_/Y _4717_/Y VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__o2bb2a_1
Xhold2823 _7631_/Q VGND VGND VPWR VPWR _6784_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2834 _7094_/Q VGND VGND VPWR VPWR hold2834/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout485_A _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2845 hold594/X VGND VGND VPWR VPWR _4243_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7006_ _7170_/CLK _7006_/D fanout573/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6662__A1 _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2856 _4247_/X VGND VGND VPWR VPWR hold2856/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4218_ _4218_/A0 _4217_/X _4232_/S VGND VGND VPWR VPWR _4218_/X sky130_fd_sc_hd__mux2_1
Xhold2867 hold2867/A VGND VGND VPWR VPWR _4498_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5198_ _4672_/X _4893_/Y _4873_/X _5423_/A _5196_/X VGND VGND VPWR VPWR _5200_/A
+ sky130_fd_sc_hd__o311a_1
Xhold2878 _7520_/Q VGND VGND VPWR VPWR hold2878/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2889 _7260_/Q VGND VGND VPWR VPWR hold2889/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4149_ _6935_/Q _4076_/B _6899_/Q VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6407__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5217__A2 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5622__C1 _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4976__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7393__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4440__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6717__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5925__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6193__A3 _6093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7214__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3951__A2 _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3782__B _3782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6350__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3050_A _7229_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5055__A _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4900__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3703__A2 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3148_A _7559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input46_A mgmt_gpio_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4894__A _4932_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_csclk_A _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3467__A1 _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6317__C _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6169__B1 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6708__A2 _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3449__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3520_ _5590_/A _4509_/A _4449_/B VGND VGND VPWR VPWR _3520_/X sky130_fd_sc_hd__and3_4
XFILLER_0_80_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap404 _5956_/B VGND VGND VPWR VPWR _5884_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold707 _5763_/X VGND VGND VPWR VPWR _7371_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap426 _4884_/B VGND VGND VPWR VPWR _4954_/C sky130_fd_sc_hd__clkbuf_8
Xhold718 hold718/A VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold729 _5799_/X VGND VGND VPWR VPWR _7403_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3451_ hold51/X _4025_/A _3450_/X VGND VGND VPWR VPWR _3451_/Y sky130_fd_sc_hd__a21oi_1
Xmax_cap459 _4667_/Y VGND VGND VPWR VPWR _5024_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_122_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6170_ _6170_/A1 _4116_/X _6067_/X _6169_/X VGND VGND VPWR VPWR _7604_/D sky130_fd_sc_hd__o31a_1
XFILLER_0_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7190_/CLK sky130_fd_sc_hd__clkbuf_16
X_5121_ _4722_/Y _4880_/Y _4826_/Y _4605_/Y VGND VGND VPWR VPWR _5122_/C sky130_fd_sc_hd__a211o_1
Xhold2108 hold159/X VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2119 hold2119/A VGND VGND VPWR VPWR _4441_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5447__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1407 hold7/X VGND VGND VPWR VPWR _4185_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5052_ _5052_/A _5052_/B _5052_/C VGND VGND VPWR VPWR _5056_/A sky130_fd_sc_hd__nor3_1
Xhold1418 hold46/X VGND VGND VPWR VPWR hold1418/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1429 hold222/X VGND VGND VPWR VPWR _7473_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3458__A1 _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4003_ _4003_/A _4003_/B VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5954_ _5954_/A0 _5954_/A1 _5955_/S VGND VGND VPWR VPWR _5954_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4970__C _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4905_ _5213_/B _4954_/C _5213_/C _5260_/D VGND VGND VPWR VPWR _4906_/B sky130_fd_sc_hd__nand4_2
XFILLER_0_8_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5885_ _5885_/A0 hold464/X _5892_/S VGND VGND VPWR VPWR _5885_/X sky130_fd_sc_hd__mux2_1
X_7624_ _7627_/CLK _7624_/D fanout569/X VGND VGND VPWR VPWR _7624_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5907__A0 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4836_ _4836_/A _5260_/B _4836_/C _5094_/A VGND VGND VPWR VPWR _4837_/C sky130_fd_sc_hd__nand4_1
XFILLER_0_63_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3918__C1 _3917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7555_ _7555_/CLK _7555_/D fanout594/X VGND VGND VPWR VPWR _7555_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4767_ _4860_/A _4767_/B VGND VGND VPWR VPWR _5410_/B sky130_fd_sc_hd__nor2_8
XANTENNA__6580__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6506_ _7329_/Q _6423_/X _6503_/X _6505_/X VGND VGND VPWR VPWR _6506_/X sky130_fd_sc_hd__a211o_1
X_3718_ _7030_/Q _3669_/C _5632_/B _3520_/X _7443_/Q VGND VGND VPWR VPWR _3718_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7486_ _7578_/CLK _7486_/D fanout603/X VGND VGND VPWR VPWR _7486_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4698__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4698_ _4772_/A _4797_/B _4814_/C VGND VGND VPWR VPWR _4698_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_114_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6437_ _7551_/Q _6408_/A _6434_/X _7463_/Q _6436_/X VGND VGND VPWR VPWR _6437_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5135__B2 _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3649_ _4551_/C hold56/A _4491_/C VGND VGND VPWR VPWR _3649_/X sky130_fd_sc_hd__and3_2
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6368_ _6970_/Q _6136_/B _6144_/B _6032_/Y _7024_/Q VGND VGND VPWR VPWR _6368_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5319_ _5319_/A _5531_/B _5491_/C VGND VGND VPWR VPWR _5319_/X sky130_fd_sc_hd__and3_1
X_6299_ _7056_/Q _6332_/B _6084_/X _6097_/X _7182_/Q VGND VGND VPWR VPWR _6299_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5603__A _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2620 _7373_/Q VGND VGND VPWR VPWR hold883/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_hold1515_A _7513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2631 hold866/X VGND VGND VPWR VPWR _5628_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__buf_4
Xhold2642 hold710/X VGND VGND VPWR VPWR _5772_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2653 _4423_/X VGND VGND VPWR VPWR hold888/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__buf_2
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6418__B _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__clkbuf_4
Xhold2664 hold728/X VGND VGND VPWR VPWR _5799_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2675 hold740/X VGND VGND VPWR VPWR _5871_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1930 hold354/X VGND VGND VPWR VPWR _4198_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2686 _7653_/A VGND VGND VPWR VPWR hold874/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1941 _7212_/Q VGND VGND VPWR VPWR hold416/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2697 _7244_/Q VGND VGND VPWR VPWR hold969/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1952 hold477/X VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1963 hold554/X VGND VGND VPWR VPWR _7361_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1974 _7014_/Q VGND VGND VPWR VPWR hold450/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7574__RESET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4661__A3 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1985 _4537_/X VGND VGND VPWR VPWR hold435/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6399__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1996 hold479/X VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_97_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input100_A wb_adr_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3621__B2 _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5374__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6571__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6600__C _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_9 _3902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5429__A2 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6626__B2 _7406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3612__A1 _7240_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3612__B2 _7436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2198_A _7350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5670_ _5967_/A1 _5670_/A1 _5670_/S VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__mux2_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5365__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4621_ _4947_/C _4954_/A VGND VGND VPWR VPWR _4966_/A sky130_fd_sc_hd__and2_4
XANTENNA__4799__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6562__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7340_ _7581_/CLK _7340_/D fanout584/X VGND VGND VPWR VPWR _7340_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4552_ _5840_/A1 _4552_/A1 _4556_/S VGND VGND VPWR VPWR _4552_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3915__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold504 hold504/A VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3503_ _4449_/B _5612_/B _4388_/B VGND VGND VPWR VPWR _3503_/X sky130_fd_sc_hd__and3_4
Xhold515 hold515/A VGND VGND VPWR VPWR _7310_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7271_ _7333_/CLK _7271_/D fanout582/X VGND VGND VPWR VPWR _7271_/Q sky130_fd_sc_hd__dfrtp_1
Xhold526 hold526/A VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4483_ _4483_/A0 _5852_/A0 _4484_/S VGND VGND VPWR VPWR _4483_/X sky130_fd_sc_hd__mux2_1
Xhold537 hold537/A VGND VGND VPWR VPWR _7296_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold548 _4439_/X VGND VGND VPWR VPWR _7092_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold559 hold559/A VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6222_ _7428_/Q _6094_/A _6074_/X _6094_/X _7508_/Q VGND VGND VPWR VPWR _6222_/X
+ sky130_fd_sc_hd__a32o_1
X_3434_ _7370_/Q VGND VGND VPWR VPWR _3434_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_122_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _7457_/Q _6112_/C _6079_/X _6119_/X _7401_/Q VGND VGND VPWR VPWR _6153_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6617__A1 _7565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5104_ _4888_/B _5091_/A _4817_/X _5103_/Y VGND VGND VPWR VPWR _5104_/Y sky130_fd_sc_hd__a31oi_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6617__B2 hold76/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6106_/B _6119_/A _7588_/Q _7589_/Q VGND VGND VPWR VPWR _6084_/X sky130_fd_sc_hd__and4b_4
Xhold1204 hold1204/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_0_148_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1215 hold3081/X VGND VGND VPWR VPWR hold1215/X sky130_fd_sc_hd__dlygate4sd1_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _4220_/X VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1237 _5858_/X VGND VGND VPWR VPWR _7455_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5035_ _5035_/A _5035_/B _5035_/C _5035_/D VGND VGND VPWR VPWR _5035_/Y sky130_fd_sc_hd__nor4_1
Xhold1248 hold3093/X VGND VGND VPWR VPWR hold3094/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1259 hold3118/X VGND VGND VPWR VPWR _7431_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4981__B _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3851__B2 _4174_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6986_ _7633_/CLK _6986_/D VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5937_ hold17/X _5937_/A1 _5937_/S VGND VGND VPWR VPWR _5937_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_180_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3603__A1 _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3603__B2 _7517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_12_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5868_ _5868_/A0 _5985_/A1 _5874_/S VGND VGND VPWR VPWR _5868_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6148__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7607_ _7621_/CLK _7607_/D fanout579/X VGND VGND VPWR VPWR _7607_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4819_ _4888_/B _4856_/A _5058_/D VGND VGND VPWR VPWR _5011_/B sky130_fd_sc_hd__and3b_4
XANTENNA__5356__A1 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5799_ _5997_/A1 _5799_/A1 _5802_/S VGND VGND VPWR VPWR _5799_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_145_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7538_ _7542_/CLK _7538_/D fanout581/X VGND VGND VPWR VPWR _7538_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3906__A2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6420__C _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5108__A1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6305__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7469_ _7510_/CLK _7469_/D fanout603/X VGND VGND VPWR VPWR _7469_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6320__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3140 hold3140/A VGND VGND VPWR VPWR _4528_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4563_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3151 hold3151/A VGND VGND VPWR VPWR _4540_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _5071_/C sky130_fd_sc_hd__buf_8
Xhold3162 _7535_/Q VGND VGND VPWR VPWR hold3162/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6608__B2 _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR input124/X sky130_fd_sc_hd__clkbuf_4
Xhold3173 hold3173/A VGND VGND VPWR VPWR _5804_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input148_A wb_dat_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6811_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3184 _7103_/Q VGND VGND VPWR VPWR _4425_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6818_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3195 _7610_/Q VGND VGND VPWR VPWR _6330_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2450 _7315_/Q VGND VGND VPWR VPWR hold137/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6809_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2461 _4214_/X VGND VGND VPWR VPWR hold657/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6824_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2472 hold664/X VGND VGND VPWR VPWR _4205_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2483 hold678/X VGND VGND VPWR VPWR _5592_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2494 _7223_/Q VGND VGND VPWR VPWR hold676/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1760 _5994_/X VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1771 _7290_/Q VGND VGND VPWR VPWR hold294/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4634__A3 _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1782 _4446_/X VGND VGND VPWR VPWR hold379/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1793 _5981_/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3842__A1 _7505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_168_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5595__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6792__A0 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6139__A3 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4131__B _4131_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5243__A _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7425__RESET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6614__A4 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4293__S _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6840_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6840_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6771_ _7055_/Q _6434_/B _6771_/A3 _6419_/C _7141_/Q VGND VGND VPWR VPWR _6771_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6783__A0 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3983_ _7343_/Q _3545_/X _3980_/X _3981_/X _3982_/X VGND VGND VPWR VPWR _3983_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_175_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5722_ _5722_/A _5938_/B _5731_/B _5902_/B VGND VGND VPWR VPWR _5730_/S sky130_fd_sc_hd__and4_4
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7151_/CLK sky130_fd_sc_hd__clkbuf_16
X_5653_ _5896_/A0 _5653_/A1 _5653_/S VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4604_ _4795_/C _4740_/D _4772_/A _4805_/B VGND VGND VPWR VPWR _4604_/Y sky130_fd_sc_hd__nor4_2
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3864__C _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5584_ _5815_/A1 _5584_/A1 _5586_/S VGND VGND VPWR VPWR _5584_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6550__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7323_ _7499_/CLK hold99/X fanout578/X VGND VGND VPWR VPWR _7323_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_csclk _7267_/CLK VGND VGND VPWR VPWR _6956_/CLK sky130_fd_sc_hd__clkbuf_16
X_4535_ _5583_/A0 _4535_/A1 _4538_/S VGND VGND VPWR VPWR _4535_/X sky130_fd_sc_hd__mux2_1
Xhold301 hold301/A VGND VGND VPWR VPWR _7458_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold312 hold312/A VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5852__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold323 hold323/A VGND VGND VPWR VPWR _7465_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold334 hold334/A VGND VGND VPWR VPWR hold334/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold345 hold345/A VGND VGND VPWR VPWR _7314_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7254_ _7264_/CLK _7254_/D fanout565/X VGND VGND VPWR VPWR _7254_/Q sky130_fd_sc_hd__dfrtp_1
Xhold356 _7058_/Q VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4466_ _4466_/A0 _5979_/A0 _4466_/S VGND VGND VPWR VPWR _4466_/X sky130_fd_sc_hd__mux2_1
Xhold367 hold367/A VGND VGND VPWR VPWR _7418_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold378 hold378/A VGND VGND VPWR VPWR hold378/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold389 _5721_/X VGND VGND VPWR VPWR _7334_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6205_ _7291_/Q _6072_/B _6144_/B _6032_/Y _7347_/Q VGND VGND VPWR VPWR _6205_/X
+ sky130_fd_sc_hd__a32o_1
X_3417_ _7506_/Q VGND VGND VPWR VPWR _3417_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7185_ _7186_/CLK _7185_/D _6833_/A VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_4
X_4397_ _5815_/A1 _4397_/A1 _4399_/S VGND VGND VPWR VPWR _4397_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout398_A _4932_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _7296_/Q _6136_/B _6136_/C VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__and3_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 hold2418/X VGND VGND VPWR VPWR hold2419/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1012 hold2603/X VGND VGND VPWR VPWR hold2604/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 hold2834/X VGND VGND VPWR VPWR hold2835/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6067_/A _6931_/Q VGND VGND VPWR VPWR _6067_/X sky130_fd_sc_hd__and2_4
XFILLER_0_84_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4992__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1034 hold2906/X VGND VGND VPWR VPWR _7544_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1045 hold2854/X VGND VGND VPWR VPWR hold2855/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout565_A fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1056 _4474_/X VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 _5669_/X VGND VGND VPWR VPWR _7287_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5018_ _5034_/C _5018_/B VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__nand2_1
Xhold1078 hold2926/X VGND VGND VPWR VPWR hold2927/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _4451_/X VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6369__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6415__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6969_ _7196_/CLK _6969_/D fanout589/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_76_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6526__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5762__S _5766_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold890 _5674_/X VGND VGND VPWR VPWR _7292_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5063__A _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5213__D _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4068__B2 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2280 _5856_/X VGND VGND VPWR VPWR hold558/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2291 _7414_/Q VGND VGND VPWR VPWR hold602/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1590 hold239/X VGND VGND VPWR VPWR _5770_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5280__A3 _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6765__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3579__B1 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4240__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6517__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3594__A3 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4142__A _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4320_ _3607_/Y _4320_/A1 _4321_/S VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_140_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4796__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6296__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4288__S _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4251_ _4251_/A0 hold464/X _4258_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
X_4182_ _4182_/A0 _5840_/A1 _4190_/S VGND VGND VPWR VPWR _4182_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6048__A2 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7432__SET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3806__A1 _7529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3806__B2 _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2697_A _7244_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4317__A _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3859__C _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5008__B1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6823_ _4114_/B _7105_/D _6823_/A3 _4428_/Y _4430_/B VGND VGND VPWR VPWR _7645_/D
+ sky130_fd_sc_hd__o41ai_2
XANTENNA__6756__B1 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6220__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6754_ _7176_/Q _6747_/B _6747_/C _6443_/X _7196_/Q VGND VGND VPWR VPWR _6754_/X
+ sky130_fd_sc_hd__a32o_1
X_3966_ _6911_/Q _5612_/B _5947_/A _5713_/A _7327_/Q VGND VGND VPWR VPWR _3966_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4231__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6771__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5705_ _5903_/A0 _5705_/A1 _5712_/S VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3585__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6685_ _7042_/Q _6408_/B _6462_/X _7032_/Q _6684_/X VGND VGND VPWR VPWR _6685_/X
+ sky130_fd_sc_hd__a221o_2
X_3897_ _7002_/Q _4322_/A _3889_/X _3892_/X _3896_/X VGND VGND VPWR VPWR _3897_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3990__B1 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5636_ _5979_/A0 _5636_/A1 _5639_/S VGND VGND VPWR VPWR _5636_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5567_ _4778_/A _5410_/X _5308_/C _5148_/C _5308_/A VGND VGND VPWR VPWR _5568_/C
+ sky130_fd_sc_hd__a2111oi_1
X_7306_ _7501_/CLK _7306_/D fanout580/X VGND VGND VPWR VPWR _7306_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3742__B1 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold120 hold120/A VGND VGND VPWR VPWR hold120/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold131 _3496_/A VGND VGND VPWR VPWR _3511_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4518_ hold318/X _5815_/A1 _4520_/S VGND VGND VPWR VPWR _4518_/X sky130_fd_sc_hd__mux2_1
Xhold142 hold142/A VGND VGND VPWR VPWR _7451_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold153 _6900_/Q VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5498_ _5053_/C _5553_/A1 _5328_/X _5497_/X VGND VGND VPWR VPWR _5499_/B sky130_fd_sc_hd__a31o_1
Xhold164 hold164/A VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7237_ _7239_/CLK _7237_/D fanout566/X VGND VGND VPWR VPWR _7237_/Q sky130_fd_sc_hd__dfstp_2
Xhold175 _7246_/Q VGND VGND VPWR VPWR hold175/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6287__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold186 hold186/A VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4449_ _4473_/A _4449_/B _4455_/C _4551_/D VGND VGND VPWR VPWR _4454_/S sky130_fd_sc_hd__and4_2
Xfanout600 fanout601/X VGND VGND VPWR VPWR fanout600/X sky130_fd_sc_hd__buf_12
Xhold197 _7289_/Q VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout611 _4909_/D VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__buf_12
XFILLER_0_95_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7168_ _7213_/CLK _7168_/D fanout590/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6119_/A _6119_/B _6121_/A _6121_/C VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__and4_4
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7505_/CLK _7099_/D fanout601/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1797_A _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6762__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5970__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3981__B1 _7447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6514__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input76_A qspi_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6278__A2 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5789__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6450__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6738__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6202__A2 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3820_ _6876_/Q _4509_/A _5603_/B _3564_/X _7361_/Q VGND VGND VPWR VPWR _3828_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4213__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3751_ _6877_/Q _5866_/B _5632_/B _4497_/A _7155_/Q VGND VGND VPWR VPWR _3751_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_156_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5961__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_59_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2180_A _7292_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6470_ _7503_/Q _6466_/X _6467_/X _7415_/Q _6469_/X VGND VGND VPWR VPWR _6471_/D
+ sky130_fd_sc_hd__a221o_1
X_3682_ _5590_/A _3931_/D _5640_/C VGND VGND VPWR VPWR _3682_/X sky130_fd_sc_hd__and3_2
XANTENNA__4303__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5421_ _4595_/Y _4605_/Y _4956_/A _4834_/Y _4583_/B VGND VGND VPWR VPWR _5422_/B
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6498__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput203 wire365/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3724__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput214 _4149_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
X_5352_ _5213_/C _4940_/D _5346_/X _5217_/X _5213_/B VGND VGND VPWR VPWR _5352_/Y
+ sky130_fd_sc_hd__a32oi_4
Xoutput225 _7662_/X VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
Xoutput236 _7670_/X VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput247 _4125_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
X_4303_ _4346_/C _5623_/B _5640_/D VGND VGND VPWR VPWR _4308_/S sky130_fd_sc_hd__and3_2
Xoutput258 _7243_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
XANTENNA__3861__D _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput269 _6919_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
X_5283_ _5059_/B _5115_/X _5282_/X VGND VGND VPWR VPWR _5481_/A sky130_fd_sc_hd__a21oi_1
X_7022_ _7409_/CLK _7022_/D fanout568/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfrtp_4
X_4234_ _5651_/A1 _5903_/A0 _4248_/S VGND VGND VPWR VPWR _4234_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4165_ _6938_/Q input93/X _7262_/Q VGND VGND VPWR VPWR _4165_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_156_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4096_ input123/X input122/X _4096_/C _4096_/D VGND VGND VPWR VPWR _4096_/X sky130_fd_sc_hd__and4bb_2
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4452__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6729__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6806_ _7109_/Q _6806_/A2 _6806_/B1 wire463/A _6805_/X VGND VGND VPWR VPWR _6806_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout430_A _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4204__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4998_ _5024_/A1 _4669_/X _5038_/A _4974_/B VGND VGND VPWR VPWR _5018_/B sky130_fd_sc_hd__o211a_2
XANTENNA__6744__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5952__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3949_ _7016_/Q _4346_/C _5619_/B _3948_/X VGND VGND VPWR VPWR _3949_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3465__A_N _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6737_ _6991_/Q _6420_/B _6462_/X _7034_/Q VGND VGND VPWR VPWR _6737_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_190_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6668_ _7056_/Q _6600_/B _6651_/C _6452_/X _7021_/Q VGND VGND VPWR VPWR _6668_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5619_ _5619_/A _5619_/B _5640_/D VGND VGND VPWR VPWR _5620_/S sky130_fd_sc_hd__and3_1
XFILLER_0_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6599_ _6599_/A1 _4116_/X _6067_/X _6598_/X VGND VGND VPWR VPWR _7620_/D sky130_fd_sc_hd__o31a_1
XANTENNA__3715__B1 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7181__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3730__A3 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5468__B1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout430 _6574_/C VGND VGND VPWR VPWR _6771_/A3 sky130_fd_sc_hd__buf_12
Xfanout441 _6424_/C VGND VGND VPWR VPWR _6574_/B sky130_fd_sc_hd__buf_12
XANTENNA__6680__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout474 hold84/X VGND VGND VPWR VPWR _5754_/A1 sky130_fd_sc_hd__buf_12
Xfanout485 _5995_/A1 VGND VGND VPWR VPWR _5815_/A1 sky130_fd_sc_hd__buf_6
XANTENNA__4883__C _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout496 _5903_/A0 VGND VGND VPWR VPWR _5714_/A0 sky130_fd_sc_hd__clkbuf_16
XANTENNA_input130_A wb_adr_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6904__CLK _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6432__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4443__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6196__A1 _7443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__B2 _7307_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5943__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_60_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6499__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6671__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3470__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5226__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5970_ _5970_/A0 _5997_/A1 hold13/X VGND VGND VPWR VPWR _5970_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4434__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4921_ _5213_/A _4932_/B _4929_/A _5260_/D VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__and4_1
XFILLER_0_176_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7640_ _7646_/CLK _7640_/D _4309_/B VGND VGND VPWR VPWR _7640_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6082__A _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6187__A1 _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4852_ _4583_/B _4595_/Y _4695_/Y _7110_/Q VGND VGND VPWR VPWR _5294_/A sky130_fd_sc_hd__o31a_4
XANTENNA__6187__B2 _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3803_ _7353_/Q _5803_/A _4212_/A _5758_/A _7369_/Q VGND VGND VPWR VPWR _3803_/X
+ sky130_fd_sc_hd__a32o_1
X_7571_ _7575_/CLK _7571_/D fanout596/X VGND VGND VPWR VPWR _7571_/Q sky130_fd_sc_hd__dfrtp_4
X_4783_ _4772_/A _4801_/B _5410_/A _5410_/B VGND VGND VPWR VPWR _4783_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_0_90_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6522_ _6521_/X _6522_/A1 _6649_/S VGND VGND VPWR VPWR _6522_/X sky130_fd_sc_hd__mux2_1
X_3734_ _3923_/S _3734_/B VGND VGND VPWR VPWR _3734_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6453_ _7479_/Q _6447_/C _6459_/C _6452_/X _7343_/Q VGND VGND VPWR VPWR _6453_/X
+ sky130_fd_sc_hd__a32o_1
X_3665_ _4473_/A _4551_/A _4551_/C VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__and3_2
XFILLER_0_113_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5404_ _5410_/A _5404_/B _5404_/C _5404_/D VGND VGND VPWR VPWR _5405_/C sky130_fd_sc_hd__nand4_1
X_6384_ _7191_/Q _6119_/A _6106_/B _6136_/B _6144_/C VGND VGND VPWR VPWR _6384_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5162__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3596_ _7293_/Q _3543_/X _3592_/X _3593_/X _3595_/X VGND VGND VPWR VPWR _3606_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5335_ _5038_/B _5030_/C _5339_/B _5334_/X VGND VGND VPWR VPWR _5335_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5860__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2802 hold2802/A VGND VGND VPWR VPWR hold2802/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5266_ _5266_/A _5266_/B _5256_/X VGND VGND VPWR VPWR _5266_/Y sky130_fd_sc_hd__nor3b_1
Xhold2813 _7117_/Q VGND VGND VPWR VPWR hold2813/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2824 hold2824/A VGND VGND VPWR VPWR hold2824/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2835 hold2835/A VGND VGND VPWR VPWR _4442_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7005_ _7212_/CLK _7005_/D fanout574/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5465__A3 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2846 _4243_/X VGND VGND VPWR VPWR hold595/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6662__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4217_ _4251_/A0 hold464/X _4231_/S VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
Xhold2857 _7415_/Q VGND VGND VPWR VPWR hold2857/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout380_A _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5197_ _4858_/Y _5528_/A3 _4873_/X _4672_/X _5046_/A VGND VGND VPWR VPWR _5423_/A
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout478_A hold2072/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2868 _7635_/Q VGND VGND VPWR VPWR _6791_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2879 hold2879/A VGND VGND VPWR VPWR _5931_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4148_ _7268_/Q input81/X _4174_/B VGND VGND VPWR VPWR _4148_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_183_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4079_ _6865_/A _6869_/B VGND VGND VPWR VPWR _4079_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6178__A1 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6423__C _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5689__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3951__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4878__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6350__A1 _7199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6350__B2 _7154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5055__B _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5770__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6653__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input39_A mgmt_gpio_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5861__A0 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3210_A _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5208__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4416__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_761 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6708__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7399__SET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5392__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap405 wire406/X VGND VGND VPWR VPWR _5956_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold708 hold708/A VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_80_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold719 _5675_/X VGND VGND VPWR VPWR _7293_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3450_ _4025_/A _3450_/B VGND VGND VPWR VPWR _3450_/X sky130_fd_sc_hd__and2b_1
XANTENNA__6341__A1 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap449 _5399_/D VGND VGND VPWR VPWR _4846_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5120_ _4845_/X _5180_/B _5119_/X VGND VGND VPWR VPWR _5122_/B sky130_fd_sc_hd__a21oi_1
Xhold2109 _7355_/Q VGND VGND VPWR VPWR hold139/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5051_ _5051_/A _5051_/B _5051_/C VGND VGND VPWR VPWR _5052_/C sky130_fd_sc_hd__nand3_1
XANTENNA__6644__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1408 _4185_/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1419 _5614_/X VGND VGND VPWR VPWR _5618_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4655__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5852__A0 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4002_ _6910_/Q _4002_/B _4006_/A VGND VGND VPWR VPWR _4003_/B sky130_fd_sc_hd__and3_1
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4407__A1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7220__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5953_ _5953_/A0 _5953_/A1 _5955_/S VGND VGND VPWR VPWR _5953_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5080__B2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2777_A _7141_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4904_ _4904_/A _4904_/B VGND VGND VPWR VPWR _4906_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5884_ _5938_/C _5884_/B _5992_/D VGND VGND VPWR VPWR _5884_/X sky130_fd_sc_hd__and3_4
XANTENNA__3630__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7623_ _7623_/CLK _7623_/D fanout575/X VGND VGND VPWR VPWR _7623_/Q sky130_fd_sc_hd__dfrtp_1
X_4835_ _4583_/B _4595_/Y _4832_/Y _4834_/Y _4956_/A VGND VGND VPWR VPWR _4837_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_173_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5855__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4766_ _4766_/A _4766_/B VGND VGND VPWR VPWR _4766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6580__A1 _7292_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7554_ _7575_/CLK _7554_/D fanout595/X VGND VGND VPWR VPWR _7554_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_172_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6505_ _7297_/Q _6420_/A _6421_/X _7321_/Q _6504_/X VGND VGND VPWR VPWR _6505_/X
+ sky130_fd_sc_hd__a221o_1
X_3717_ _7459_/Q _5857_/A _3713_/X _3714_/X _3716_/X VGND VGND VPWR VPWR _3717_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_16_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7485_ _7565_/CLK hold81/X fanout603/X VGND VGND VPWR VPWR _7485_/Q sky130_fd_sc_hd__dfrtp_4
X_4697_ _4772_/A _4797_/B _4814_/C VGND VGND VPWR VPWR _5091_/C sky130_fd_sc_hd__and3_4
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4698__C _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3648_ _5803_/A _4388_/B _3931_/D VGND VGND VPWR VPWR _3648_/X sky130_fd_sc_hd__and3_2
X_6436_ _7319_/Q _6421_/X _6435_/X _7511_/Q VGND VGND VPWR VPWR _6436_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4343__A0 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6367_ _7115_/Q _6317_/C _6332_/C _7034_/Q _6366_/X VGND VGND VPWR VPWR _6367_/X
+ sky130_fd_sc_hd__a221o_1
X_3579_ _5640_/C _5623_/B _3578_/X _4248_/S input69/X VGND VGND VPWR VPWR _3579_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3697__A2 _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5318_ _4583_/B _4821_/Y _4802_/Y _4595_/Y VGND VGND VPWR VPWR _5531_/B sky130_fd_sc_hd__a211o_1
X_6298_ _7172_/Q _6110_/X _6112_/X _6874_/Q _6297_/X VGND VGND VPWR VPWR _6303_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2610 _7341_/Q VGND VGND VPWR VPWR hold876/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2621 hold883/X VGND VGND VPWR VPWR _5765_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__B1 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5603__B _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__6635__A2 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2632 _5628_/X VGND VGND VPWR VPWR hold867/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5249_ _4659_/Y _4946_/Y _5247_/X VGND VGND VPWR VPWR _5249_/Y sky130_fd_sc_hd__o21ai_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2643 _7547_/Q VGND VGND VPWR VPWR hold680/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2654 _7459_/Q VGND VGND VPWR VPWR hold692/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1920 _7226_/Q VGND VGND VPWR VPWR hold545/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6418__C _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2665 _7371_/Q VGND VGND VPWR VPWR hold706/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2676 _5871_/X VGND VGND VPWR VPWR hold741/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1931 _4198_/X VGND VGND VPWR VPWR hold355/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__clkbuf_4
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1942 hold416/X VGND VGND VPWR VPWR _5585_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2687 hold874/X VGND VGND VPWR VPWR _4249_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2698 hold969/X VGND VGND VPWR VPWR _5615_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1953 _7034_/Q VGND VGND VPWR VPWR hold446/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1964 _7409_/Q VGND VGND VPWR VPWR hold518/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1975 hold450/X VGND VGND VPWR VPWR _4338_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1986 _7049_/Q VGND VGND VPWR VPWR hold370/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1997 _7023_/Q VGND VGND VPWR VPWR hold504/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6399__A1 _6961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6434__B _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3621__A2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5765__S _5766_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3909__B1 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6571__A1 _7283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold3160_A _7001_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4689__B1_N _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3688__A2 _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6626__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5429__A3 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4129__B _4129_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4627__B1_N _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5062__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5062__B2 _4744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3612__A2 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4620_ _4616_/Y _4617_/Y _4618_/Y _4615_/Y VGND VGND VPWR VPWR _4657_/A sky130_fd_sc_hd__a22oi_4
XFILLER_0_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6562__A1 _7315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6562__B2 _7483_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4551_ _4551_/A _5866_/B _4551_/C _4551_/D VGND VGND VPWR VPWR _4556_/S sky130_fd_sc_hd__nand4_4
XANTENNA__3915__A3 _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3502_ _3576_/C _3576_/B VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__and2_4
X_7270_ _7530_/CLK _7270_/D fanout602/X VGND VGND VPWR VPWR _7270_/Q sky130_fd_sc_hd__dfrtp_1
Xhold505 _4349_/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4482_ _4482_/A0 _5914_/A1 _4484_/S VGND VGND VPWR VPWR _4482_/X sky130_fd_sc_hd__mux2_1
Xhold516 hold516/A VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold527 hold527/A VGND VGND VPWR VPWR _7502_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4325__A0 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold538 hold538/A VGND VGND VPWR VPWR hold538/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6221_ _7324_/Q _6116_/B _6081_/X _6090_/X _7380_/Q VGND VGND VPWR VPWR _6221_/X
+ sky130_fd_sc_hd__a32o_1
Xhold549 hold549/A VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3433_ _7378_/Q VGND VGND VPWR VPWR _3433_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3679__A2 _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5704__A _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _7481_/Q _6112_/X _6151_/X _6150_/X _6149_/X VGND VGND VPWR VPWR _6152_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5103_ _5563_/A1 _4806_/Y _4844_/Y _5102_/Y _5101_/Y VGND VGND VPWR VPWR _5103_/Y
+ sky130_fd_sc_hd__o311ai_2
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6617__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _7455_/Q _6094_/A _6079_/X _6082_/X _7319_/Q VGND VGND VPWR VPWR _6083_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 hold2871/X VGND VGND VPWR VPWR hold1205/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1216 hold1216/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 hold3001/X VGND VGND VPWR VPWR hold3002/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5038_/A _5038_/B _5034_/C VGND VGND VPWR VPWR _5035_/C sky130_fd_sc_hd__and3_1
Xhold1238 hold2957/X VGND VGND VPWR VPWR hold2958/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1249 _5894_/X VGND VGND VPWR VPWR _7487_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_164_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3851__A2 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6985_ _7633_/CLK _6985_/D VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6250__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5936_ hold61/X _5936_/A1 _5937_/S VGND VGND VPWR VPWR _5936_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_193_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5867_ _5867_/A0 _5993_/A1 _5874_/S VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7606_ _7623_/CLK _7606_/D fanout576/X VGND VGND VPWR VPWR _7606_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout510_A _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4818_ _4818_/A _4818_/B _4818_/C VGND VGND VPWR VPWR _4824_/A sky130_fd_sc_hd__nor3_1
XANTENNA__5356__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A input164/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5798_ _5987_/A1 _5798_/A1 _5802_/S VGND VGND VPWR VPWR _5798_/X sky130_fd_sc_hd__mux2_1
X_7537_ _7537_/CLK _7537_/D fanout577/X VGND VGND VPWR VPWR _7537_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4749_ _4814_/C _4608_/Y _4657_/C VGND VGND VPWR VPWR _4884_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7468_ _7565_/CLK _7468_/D fanout599/X VGND VGND VPWR VPWR _7468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_160_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6419_ _6419_/A _6419_/B _6419_/C _6419_/D VGND VGND VPWR VPWR _6419_/Y sky130_fd_sc_hd__nor4_1
X_7399_ _7457_/CLK _7399_/D fanout586/X VGND VGND VPWR VPWR _7399_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5614__A _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3130 _7256_/Q VGND VGND VPWR VPWR hold3130/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3141 _7051_/Q VGND VGND VPWR VPWR hold3141/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4563_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3152 _7471_/Q VGND VGND VPWR VPWR hold3152/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _5071_/B sky130_fd_sc_hd__buf_8
Xhold3163 hold3163/A VGND VGND VPWR VPWR _5948_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR _4786_/C sky130_fd_sc_hd__buf_4
Xhold3174 _7220_/Q VGND VGND VPWR VPWR _3609_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6815_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4619__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2440 _5605_/X VGND VGND VPWR VPWR hold646/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3185 _7104_/Q VGND VGND VPWR VPWR _4425_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2451 hold137/X VGND VGND VPWR VPWR _5700_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6821_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3196 _6307_/X VGND VGND VPWR VPWR _7610_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6812_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2462 _7043_/Q VGND VGND VPWR VPWR hold981/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput169 wb_stb_i VGND VGND VPWR VPWR _4093_/B sky130_fd_sc_hd__buf_4
Xhold2473 _7114_/Q VGND VGND VPWR VPWR hold983/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2484 _5592_/X VGND VGND VPWR VPWR hold679/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2495 hold676/X VGND VGND VPWR VPWR _5589_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1750 _7485_/Q VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1761 _7546_/Q VGND VGND VPWR VPWR hold302/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1772 hold294/X VGND VGND VPWR VPWR _5672_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4634__A4 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1783 _7211_/Q VGND VGND VPWR VPWR hold418/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1794 _7554_/Q VGND VGND VPWR VPWR hold364/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3842__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3006_A _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6241__B1 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_168_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7191_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6529__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4555__A0 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output262_A _7226_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6058__C _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6480__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3833__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7465__RESET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6074__B _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6232__B1 _6116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3982_ _7244_/Q _3590_/C _3519_/B _3569_/X _7487_/Q VGND VGND VPWR VPWR _3982_/X
+ sky130_fd_sc_hd__a32o_1
X_6770_ _7126_/Q _6420_/C _6455_/X _7201_/Q _6769_/X VGND VGND VPWR VPWR _6773_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3597__A1 hold76/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5721_ _5955_/A1 _5721_/A1 _5721_/S VGND VGND VPWR VPWR _5721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3597__B2 _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2475_A _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6090__A _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4603__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5652_ _5967_/A1 _5652_/A1 _5658_/S VGND VGND VPWR VPWR _5652_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6535__A1 _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4546__A0 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4603_ _4795_/C _4740_/D VGND VGND VPWR VPWR _5260_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4322__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5583_ _5583_/A0 _5583_/A1 _5586_/S VGND VGND VPWR VPWR _5583_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7455__SET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7322_ _7429_/CLK _7322_/D fanout583/X VGND VGND VPWR VPWR _7322_/Q sky130_fd_sc_hd__dfrtp_4
X_4534_ _5840_/A1 _4534_/A1 _4538_/S VGND VGND VPWR VPWR _4534_/X sky130_fd_sc_hd__mux2_1
Xhold302 hold302/A VGND VGND VPWR VPWR hold302/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold313 hold313/A VGND VGND VPWR VPWR _7529_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold324 hold324/A VGND VGND VPWR VPWR hold324/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6299__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold335 hold335/A VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7253_ _7264_/CLK _7253_/D fanout565/X VGND VGND VPWR VPWR _7253_/Q sky130_fd_sc_hd__dfrtp_1
Xhold346 hold346/A VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4465_ _4465_/A0 _5852_/A0 _4466_/S VGND VGND VPWR VPWR _4465_/X sky130_fd_sc_hd__mux2_1
Xhold357 hold357/A VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold368 hold368/A VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2907_A _7560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3416_ _7514_/Q VGND VGND VPWR VPWR _3416_/Y sky130_fd_sc_hd__inv_2
Xhold379 hold379/A VGND VGND VPWR VPWR _7098_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6204_ _7363_/Q _6093_/X _6106_/X _7395_/Q _6203_/X VGND VGND VPWR VPWR _6204_/X
+ sky130_fd_sc_hd__a221o_1
X_7184_ _7186_/CLK _7184_/D fanout588/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfstp_4
X_4396_ hold43/X _4396_/A1 _4399_/S VGND VGND VPWR VPWR _4396_/X sky130_fd_sc_hd__mux2_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _7344_/Q _6032_/Y _6317_/C _7384_/Q _6134_/X VGND VGND VPWR VPWR _6135_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _4489_/X VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1013 hold2743/X VGND VGND VPWR VPWR hold2744/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1024 hold2836/X VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6066_ _4099_/D _7584_/Q _6065_/Y _6062_/X _6066_/B2 VGND VGND VPWR VPWR _6066_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1035 hold2737/X VGND VGND VPWR VPWR hold2738/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__C1 _3806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1046 hold2856/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1057 hold2570/X VGND VGND VPWR VPWR hold2571/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5017_ _5006_/Y _5008_/X _5016_/Y VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__a21oi_1
Xhold1068 hold2841/X VGND VGND VPWR VPWR hold2842/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1079 hold2928/X VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_169_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3824__A2 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6223__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6968_ _7196_/CLK _6968_/D fanout588/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_177_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5919_ _5919_/A0 _5991_/A1 _5919_/S VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__mux2_1
X_6899_ _7075_/CLK _6899_/D _6849_/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5329__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6526__A1 _7562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6526__B2 _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4537__A0 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5328__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3760__A1 _6991_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3760__B2 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input160_A wb_dat_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold880 hold880/A VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold891 hold891/A VGND VGND VPWR VPWR hold891/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2270 _7472_/Q VGND VGND VPWR VPWR hold568/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input21_A mask_rev_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2281 _7291_/Q VGND VGND VPWR VPWR hold2281/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2292 hold602/X VGND VGND VPWR VPWR _5811_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1580 _7484_/Q VGND VGND VPWR VPWR hold227/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1591 _5770_/X VGND VGND VPWR VPWR hold240/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_58_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6765__A1 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6765__B2 _7116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3579__A1 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3751__B2 _7155_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4250_ _4250_/A1 hold284/X _4168_/D _4231_/S hold48/X VGND VGND VPWR VPWR _4258_/S
+ sky130_fd_sc_hd__o311a_4
XFILLER_0_129_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4181_ _4076_/B _4181_/A1 _4429_/B VGND VGND VPWR VPWR _4181_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5404__D _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7646__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5256__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6453__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3806__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5008__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6205__B1 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6822_ _6821_/X _6822_/A1 _6822_/S VGND VGND VPWR VPWR _7644_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_77_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6753_ _7131_/Q _6424_/X _6427_/X _7121_/Q VGND VGND VPWR VPWR _6753_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_161_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3965_ _7455_/Q _5785_/B _5866_/B _3964_/X VGND VGND VPWR VPWR _3965_/X sky130_fd_sc_hd__a31o_2
XFILLER_0_190_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5704_ _5704_/A _5902_/B VGND VGND VPWR VPWR _5712_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_70_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6508__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3896_ _7424_/Q _3537_/X _3862_/X _3893_/X _3895_/X VGND VGND VPWR VPWR _3896_/X
+ sky130_fd_sc_hd__a2111o_1
X_6684_ _7027_/Q _6459_/B _6459_/C _6460_/X _7113_/Q VGND VGND VPWR VPWR _6684_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3990__B2 _7303_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5635_ _5986_/A1 _5635_/A1 _5639_/S VGND VGND VPWR VPWR _5635_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5863__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5566_ _5566_/A1 wire462/X _5565_/X _5557_/X VGND VGND VPWR VPWR _7207_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_13_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold110 hold110/A VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7305_ _7359_/CLK _7305_/D fanout576/X VGND VGND VPWR VPWR _7305_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3742__A1 _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold121 hold121/A VGND VGND VPWR VPWR _7453_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold132 _3519_/B VGND VGND VPWR VPWR _5614_/B sky130_fd_sc_hd__buf_4
X_4517_ _4517_/A0 _5583_/A0 _4520_/S VGND VGND VPWR VPWR _4517_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5497_ _5203_/B _5553_/A1 _5425_/X _5172_/X VGND VGND VPWR VPWR _5497_/X sky130_fd_sc_hd__a31o_1
Xhold143 hold143/A VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold154 _3466_/X VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold165 hold165/A VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold176 hold176/A VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7236_ _7363_/CLK _7236_/D fanout575/X VGND VGND VPWR VPWR _7236_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6287__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4448_ _4448_/A0 _5991_/A1 _4448_/S VGND VGND VPWR VPWR _4448_/X sky130_fd_sc_hd__mux2_1
Xfanout601 fanout602/X VGND VGND VPWR VPWR fanout601/X sky130_fd_sc_hd__buf_12
Xhold187 _7492_/Q VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout612 _4909_/D VGND VGND VPWR VPWR _4772_/A sky130_fd_sc_hd__buf_12
Xhold198 hold198/A VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5495__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6692__B1 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7167_ _7170_/CLK _7167_/D fanout573/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_4
X_4379_ _4379_/A0 _5914_/A1 _4381_/S VGND VGND VPWR VPWR _4379_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_95_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6110_/A _6115_/X _6117_/X _6114_/X _6108_/X VGND VGND VPWR VPWR _6118_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_7098_ _7197_/CLK _7098_/D fanout601/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6444__B1 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6047_/Y _6048_/X _6051_/C _6019_/Y _6435_/B VGND VGND VPWR VPWR _7595_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3412__A _7546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6426__C _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5058__B _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3981__B2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5773__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input69_A mgmt_gpio_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5074__A _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6278__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7186_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5238__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_csclk _7267_/CLK VGND VGND VPWR VPWR _7096_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_188_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ _7378_/Q _3498_/X _3745_/X _3747_/X _3749_/X VGND VGND VPWR VPWR _3750_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6071__C _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6070__A_N _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3681_ _7065_/Q _4394_/A _3676_/X _3677_/X _3680_/X VGND VGND VPWR VPWR _3681_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_171_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5174__B1 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5420_ _4595_/Y _4956_/A _4730_/Y _5529_/A _5419_/X VGND VGND VPWR VPWR _5422_/A
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3724__A1 _6923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput204 _4143_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
X_5351_ _4601_/Y _4956_/B _4726_/Y _4622_/Y VGND VGND VPWR VPWR _5355_/B sky130_fd_sc_hd__a211o_1
XANTENNA__3724__B2 _7323_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput215 _7654_/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
Xoutput226 _7663_/X VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
Xoutput237 _4148_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
Xoutput248 _4126_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
X_4302_ _3570_/Y _4302_/A1 _4302_/S VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__mux2_1
Xoutput259 _7223_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
XANTENNA__6269__A3 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5282_ _5282_/A _5282_/B _5399_/D _5282_/D VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__and4_1
XANTENNA__5477__A1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7021_ _7409_/CLK _7021_/D fanout568/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6674__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4233_ _6839_/B _3541_/Y _4248_/S _4215_/X hold48/X VGND VGND VPWR VPWR _4249_/S
+ sky130_fd_sc_hd__o221a_4
X_4164_ _7091_/Q _4164_/A1 _7259_/Q VGND VGND VPWR VPWR _4164_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5229__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4095_ _5115_/A _4095_/B _4095_/C _4095_/D VGND VGND VPWR VPWR _4096_/D sky130_fd_sc_hd__and4_1
XANTENNA__4328__A _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5858__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6729__B2 _6965_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6805_ _7111_/Q _6805_/A2 _6805_/B1 _7110_/Q VGND VGND VPWR VPWR _6805_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_175_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4997_ _5158_/A _4997_/B _5404_/C _5410_/B VGND VGND VPWR VPWR _5028_/C sky130_fd_sc_hd__nand4_4
XFILLER_0_58_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout423_A _6073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6736_ _7044_/Q _6408_/B _6460_/X _7115_/Q _6735_/X VGND VGND VPWR VPWR _6736_/X
+ sky130_fd_sc_hd__a221o_1
X_3948_ _5587_/C _5623_/B _3864_/X _7222_/Q _3947_/X VGND VGND VPWR VPWR _3948_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_190_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3963__A1 _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3963__B2 _6967_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6667_ _7197_/Q _6463_/A _6771_/A3 _6463_/X _7162_/Q VGND VGND VPWR VPWR _6667_/X
+ sky130_fd_sc_hd__a32o_1
X_3879_ _3879_/A _3879_/B _3879_/C _3879_/D VGND VGND VPWR VPWR _3922_/A sky130_fd_sc_hd__nor4_4
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5618_ _5618_/A0 _5951_/A1 _5618_/S VGND VGND VPWR VPWR _5618_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6598_ _6649_/S _6598_/A2 _6777_/S _6597_/X VGND VGND VPWR VPWR _6598_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5549_ _5342_/A _5094_/A wire536/X _5343_/A _5343_/B VGND VGND VPWR VPWR _5550_/D
+ sky130_fd_sc_hd__a311oi_4
XFILLER_0_131_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5468__A1 _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6665__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7219_ _4150_/A1 _7219_/D _6871_/X VGND VGND VPWR VPWR _7219_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__3479__B1 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout420 hold36/X VGND VGND VPWR VPWR _4551_/A sky130_fd_sc_hd__buf_12
Xfanout431 _6429_/X VGND VGND VPWR VPWR _6651_/C sky130_fd_sc_hd__buf_12
Xfanout442 _6144_/B VGND VGND VPWR VPWR _6136_/C sky130_fd_sc_hd__buf_12
XANTENNA_hold1705_A _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6680__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout475 hold2072/X VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__buf_6
Xfanout486 _5995_/A1 VGND VGND VPWR VPWR _5896_/A0 sky130_fd_sc_hd__buf_12
Xfanout497 hold464/X VGND VGND VPWR VPWR _5903_/A0 sky130_fd_sc_hd__buf_12
XANTENNA_input123_A wb_adr_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5768__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__A2 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3954__A1 _7511_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3954__B2 _7182_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4701__A _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6353__C1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6499__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3706__B2 _7483_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5171__A3 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__5459__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6656__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3890__B1 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4920_ _5213_/A _5213_/B _5183_/C _4929_/A VGND VGND VPWR VPWR _4922_/A sky130_fd_sc_hd__and4_1
XFILLER_0_157_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6082__B _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4851_ _4851_/A _4851_/B _5294_/C VGND VGND VPWR VPWR _4851_/Y sky130_fd_sc_hd__nand3_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4198__A1 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ input5/X _3486_/X _3490_/X input13/X _3801_/X VGND VGND VPWR VPWR _3802_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_145_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7570_ _7572_/CLK _7570_/D fanout596/X VGND VGND VPWR VPWR _7570_/Q sky130_fd_sc_hd__dfrtp_4
X_4782_ _4772_/A _4801_/B _5410_/A _5410_/B VGND VGND VPWR VPWR _4784_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6521_ _6501_/X _6511_/X _6520_/X _6431_/Y _7281_/Q VGND VGND VPWR VPWR _6521_/X
+ sky130_fd_sc_hd__o32a_1
X_3733_ _3686_/X _3689_/X _3733_/C _3733_/D VGND VGND VPWR VPWR _3733_/X sky130_fd_sc_hd__and4bb_2
XFILLER_0_16_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6452_ _7595_/Q _6574_/B _6651_/B _7596_/Q VGND VGND VPWR VPWR _6452_/X sky130_fd_sc_hd__and4b_4
X_3664_ _5803_/A _5640_/B _5612_/C VGND VGND VPWR VPWR _4485_/A sky130_fd_sc_hd__and3_4
XANTENNA__5698__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5403_ _5402_/X _5345_/Y _5322_/Y hold33/A _4428_/Y VGND VGND VPWR VPWR _7204_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_113_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3595_ _7453_/Q _5848_/A _3529_/X _7533_/Q _3594_/X VGND VGND VPWR VPWR _3595_/X
+ sky130_fd_sc_hd__a221o_1
X_6383_ _6971_/Q _6074_/X _6110_/A _6382_/X _6380_/X VGND VGND VPWR VPWR _6383_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_140_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5334_ _5203_/B _5553_/A1 _5328_/X _5333_/X VGND VGND VPWR VPWR _5334_/X sky130_fd_sc_hd__a31o_1
X_5265_ _5265_/A _5265_/B _5564_/A _5265_/D VGND VGND VPWR VPWR _5266_/B sky130_fd_sc_hd__nand4_1
Xhold2803 _7137_/Q VGND VGND VPWR VPWR hold2803/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2814 hold2814/A VGND VGND VPWR VPWR _4456_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2825 _7665_/A VGND VGND VPWR VPWR hold2825/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4984__C _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7004_ _7212_/CLK _7004_/D fanout573/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2836 _4442_/X VGND VGND VPWR VPWR hold2836/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4216_ _6839_/B _3481_/Y _4231_/S _4215_/X _5992_/D VGND VGND VPWR VPWR _4232_/S
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6662__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2847 _6985_/Q VGND VGND VPWR VPWR _4300_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5196_ _4672_/X _4858_/Y _4980_/X _5044_/C _5195_/X VGND VGND VPWR VPWR _5196_/X
+ sky130_fd_sc_hd__o311a_1
Xhold2858 hold2858/A VGND VGND VPWR VPWR _5813_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2869 hold2869/A VGND VGND VPWR VPWR hold2869/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5870__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4147_ _7266_/Q input78/X _4174_/B VGND VGND VPWR VPWR _4147_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_183_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4078_ _4078_/A _4078_/B _4168_/D VGND VGND VPWR VPWR _4078_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_78_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6719_ _7048_/Q _6435_/X _6446_/X _7189_/Q _6718_/X VGND VGND VPWR VPWR _6719_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4521__A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6350__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4361__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4900__A3 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6638__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4894__C _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4664__A2 _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5613__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3624__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output292_A _6926_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5392__A3 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4431__A _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold709 _4393_/X VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7419__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap428 _4657_/A VGND VGND VPWR VPWR _4954_/A sky130_fd_sc_hd__buf_6
XANTENNA__5144__A3 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6629__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5050_ _5113_/A _5399_/C _5399_/D VGND VGND VPWR VPWR _5052_/B sky130_fd_sc_hd__and3_1
XANTENNA__6644__A3 _6429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1409 hold8/X VGND VGND VPWR VPWR _5995_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4655__A2 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4001_ _6910_/Q _6909_/Q VGND VGND VPWR VPWR _4001_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__6792__S _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4700__A_N _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_189_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5604__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4606__A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5952_ _5952_/A0 hold84/X _5955_/S VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__mux2_1
XANTENNA__3615__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4903_ _5213_/B _5213_/C _5260_/D _4940_/D VGND VGND VPWR VPWR _4903_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_75_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5883_ _5883_/A0 _5955_/A1 _5883_/S VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_164_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3630__A3 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7622_ _7623_/CLK _7622_/D fanout575/X VGND VGND VPWR VPWR _7622_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4834_ _5127_/A _4834_/B VGND VGND VPWR VPWR _4834_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__3918__A1 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7553_ _7577_/CLK hold14/X fanout585/X VGND VGND VPWR VPWR _7553_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_172_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4765_ _5260_/C _4765_/B _4790_/B VGND VGND VPWR VPWR _4766_/A sky130_fd_sc_hd__and3_1
XFILLER_0_133_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6580__A2 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4979__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6504_ _7385_/Q _6413_/C _6426_/X _6451_/X _7481_/Q VGND VGND VPWR VPWR _6504_/X
+ sky130_fd_sc_hd__a32o_1
X_3716_ _7411_/Q _3493_/X _5902_/A _7499_/Q _3715_/X VGND VGND VPWR VPWR _3716_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_172_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7484_ _7510_/CLK _7484_/D fanout603/X VGND VGND VPWR VPWR _7484_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4696_ _5297_/A _4850_/B VGND VGND VPWR VPWR _5531_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6435_ _6462_/D _6435_/B _6467_/A _6600_/B VGND VGND VPWR VPWR _6435_/X sky130_fd_sc_hd__and4_4
X_3647_ _5938_/B _4551_/C hold56/A VGND VGND VPWR VPWR _3647_/X sky130_fd_sc_hd__and3_2
XFILLER_0_24_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6366_ _6965_/Q _6072_/B _6144_/B _6079_/X _7014_/Q VGND VGND VPWR VPWR _6366_/X
+ sky130_fd_sc_hd__a32o_1
X_3578_ _7627_/Q _7254_/Q _7255_/Q VGND VGND VPWR VPWR _3578_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3697__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5317_ _5317_/A _5317_/B _5317_/C _5531_/A VGND VGND VPWR VPWR _5319_/A sky130_fd_sc_hd__nor4b_1
XANTENNA_fanout490_A hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6297_ _7066_/Q _6332_/B _6332_/C _6119_/X _7132_/Q VGND VGND VPWR VPWR _6297_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2600 _5922_/X VGND VGND VPWR VPWR _7512_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2611 hold876/X VGND VGND VPWR VPWR _5729_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__B2 _7527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2622 _6933_/Q VGND VGND VPWR VPWR hold879/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2633 _7269_/Q VGND VGND VPWR VPWR hold626/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5603__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5248_ _5248_/A _5248_/B _5248_/C VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__and3_1
Xhold2644 hold680/X VGND VGND VPWR VPWR _5961_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1910 _5816_/X VGND VGND VPWR VPWR hold367/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__buf_12
XANTENNA__5843__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2655 hold692/X VGND VGND VPWR VPWR _5862_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__buf_12
Xhold1921 hold545/X VGND VGND VPWR VPWR _5593_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2666 hold706/X VGND VGND VPWR VPWR _5763_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2677 _6942_/Q VGND VGND VPWR VPWR hold881/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1932 _7195_/Q VGND VGND VPWR VPWR hold406/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1943 _7450_/Q VGND VGND VPWR VPWR hold428/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2688 _4249_/X VGND VGND VPWR VPWR hold875/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5179_ _5177_/Y _4986_/Y _5173_/X _5176_/X VGND VGND VPWR VPWR _5179_/Y sky130_fd_sc_hd__o211ai_2
Xhold2699 _7060_/Q VGND VGND VPWR VPWR hold708/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1954 hold446/X VGND VGND VPWR VPWR _4362_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1965 hold518/X VGND VGND VPWR VPWR _5806_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1976 _6959_/Q VGND VGND VPWR VPWR hold488/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6399__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1987 hold370/X VGND VGND VPWR VPWR _4380_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1998 hold504/X VGND VGND VPWR VPWR _4349_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_79_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3420__A _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6434__C _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3909__B2 _7400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6571__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5066__B _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6323__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5781__S hold49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input51_A mgmt_gpio_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3688__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5834__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3845__B1 hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4426__A _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output305_A _4166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3612__A3 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6011__B2 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6562__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4550_ _5586_/A0 _4550_/A1 _4550_/S VGND VGND VPWR VPWR _4550_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_170_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3501_ _4551_/A _5722_/A _5992_/C VGND VGND VPWR VPWR _3501_/X sky130_fd_sc_hd__and3_4
XFILLER_0_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold506 hold506/A VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6314__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5117__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4481_ _4481_/A0 _5940_/A1 _4484_/S VGND VGND VPWR VPWR _4481_/X sky130_fd_sc_hd__mux2_1
Xhold517 _5991_/X VGND VGND VPWR VPWR _7574_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold528 _7208_/Q VGND VGND VPWR VPWR hold528/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6220_ _7348_/Q _6070_/X _6218_/X _6219_/X _6217_/X VGND VGND VPWR VPWR _6220_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold539 hold539/A VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3432_ _7386_/Q VGND VGND VPWR VPWR _3432_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5704__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3679__A3 _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _7409_/Q _6121_/C _6116_/C _6136_/C VGND VGND VPWR VPWR _6151_/X sky130_fd_sc_hd__o211a_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2420_A _7119_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5453_/B _5102_/B VGND VGND VPWR VPWR _5102_/Y sky130_fd_sc_hd__nand2_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6144_/A _6116_/A _6121_/C VGND VGND VPWR VPWR _6082_/X sky130_fd_sc_hd__and3_4
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 hold1206/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XANTENNA__5825__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 hold2753/X VGND VGND VPWR VPWR hold2754/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1228 _4432_/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5033_/B _5033_/C _5033_/D VGND VGND VPWR VPWR _5035_/D sky130_fd_sc_hd__nand4_1
Xhold1239 hold2949/X VGND VGND VPWR VPWR hold2950/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3836__B1 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7415__SET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3851__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2887_A _7488_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6984_ _7633_/CLK _6984_/D VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6250__B2 _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5935_ _5998_/A1 _5935_/A1 _5937_/S VGND VGND VPWR VPWR _5935_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5866_ hold22/X _5866_/B _5938_/B _5992_/D VGND VGND VPWR VPWR _5874_/S sky130_fd_sc_hd__and4_4
XFILLER_0_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7605_ _7623_/CLK _7605_/D fanout576/X VGND VGND VPWR VPWR _7605_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4817_ _5399_/C _5089_/B _4823_/C VGND VGND VPWR VPWR _4817_/X sky130_fd_sc_hd__and3_1
XFILLER_0_146_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5797_ _5896_/A0 _5797_/A1 _5802_/S VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6553__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7536_ _7539_/CLK _7536_/D fanout578/X VGND VGND VPWR VPWR _7536_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5761__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4748_ _4887_/B _4879_/C _4748_/C VGND VGND VPWR VPWR _4748_/Y sky130_fd_sc_hd__nand3_4
XANTENNA_fanout503_A hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7467_ _7505_/CLK _7467_/D fanout601/X VGND VGND VPWR VPWR _7467_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4679_ _4679_/A _5089_/C _4679_/C VGND VGND VPWR VPWR _4679_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__6305__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4316__A1 _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6418_ _6455_/B _6424_/C _6459_/B VGND VGND VPWR VPWR _6419_/D sky130_fd_sc_hd__and3_4
XFILLER_0_141_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7398_ _7582_/CLK _7398_/D fanout585/X VGND VGND VPWR VPWR _7398_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5614__B _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6349_ _7023_/Q _6070_/X _6090_/X _7043_/Q _6348_/X VGND VGND VPWR VPWR _6349_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3120 hold3120/A VGND VGND VPWR VPWR _5822_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3415__A _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3131 hold3131/A VGND VGND VPWR VPWR _5630_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6429__C _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3142 hold3142/A VGND VGND VPWR VPWR _4383_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4563_/D sky130_fd_sc_hd__clkbuf_2
Xhold3153 hold3153/A VGND VGND VPWR VPWR _5876_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _4091_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3164 _7343_/Q VGND VGND VPWR VPWR hold3164/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR input126/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3175 _3609_/X VGND VGND VPWR VPWR _7220_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5816__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5277__C1 _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2430 _4536_/X VGND VGND VPWR VPWR hold938/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6817_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2441 _7316_/Q VGND VGND VPWR VPWR hold997/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3186 _7102_/Q VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6799_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3197 _7639_/Q VGND VGND VPWR VPWR _6807_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2452 _7255_/Q VGND VGND VPWR VPWR hold649/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6815_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2463 hold981/X VGND VGND VPWR VPWR _4373_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2474 hold983/X VGND VGND VPWR VPWR _4452_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1740 hold237/X VGND VGND VPWR VPWR _5870_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2485 _7268_/Q VGND VGND VPWR VPWR hold949/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2496 _5589_/X VGND VGND VPWR VPWR hold677/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1751 hold80/X VGND VGND VPWR VPWR _5891_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1762 hold302/X VGND VGND VPWR VPWR _5960_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1773 _7394_/Q VGND VGND VPWR VPWR hold334/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1784 hold418/X VGND VGND VPWR VPWR _5584_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1795 hold364/X VGND VGND VPWR VPWR _5969_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3842__A3 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input99_A wb_adr_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5077__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3763__C1 _3762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4307__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5807__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3833__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6232__A1 _7436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6232__B2 _7316_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3981_ _7056_/Q _5947_/B _5623_/B _7447_/Q _5848_/A VGND VGND VPWR VPWR _3981_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5720_ _5954_/A1 _5720_/A1 _5721_/S VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3597__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5651_ _5903_/A0 _5651_/A1 _5658_/S VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4603__B _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6535__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4602_ _4772_/A _4805_/B VGND VGND VPWR VPWR _5260_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_41_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5582_ _5714_/A0 _5582_/A1 _5586_/S VGND VGND VPWR VPWR _5582_/X sky130_fd_sc_hd__mux2_1
X_7321_ _7457_/CLK _7321_/D fanout586/X VGND VGND VPWR VPWR _7321_/Q sky130_fd_sc_hd__dfrtp_2
X_4533_ _4533_/A _4551_/D VGND VGND VPWR VPWR _4538_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold303 hold303/A VGND VGND VPWR VPWR _7546_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold314 hold314/A VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold325 hold325/A VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6299__B2 _7182_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7252_ _7264_/CLK _7252_/D fanout565/X VGND VGND VPWR VPWR _7252_/Q sky130_fd_sc_hd__dfrtp_4
Xhold336 hold336/A VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3793__A_N _3764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4464_ _4464_/A0 _5914_/A1 _4466_/S VGND VGND VPWR VPWR _4464_/X sky130_fd_sc_hd__mux2_1
Xhold347 hold347/A VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold358 hold358/A VGND VGND VPWR VPWR hold358/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold369 hold369/A VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6203_ _7331_/Q _6022_/X _6116_/A _6084_/X _7371_/Q VGND VGND VPWR VPWR _6203_/X
+ sky130_fd_sc_hd__a32o_1
X_3415_ _7522_/Q VGND VGND VPWR VPWR _3415_/Y sky130_fd_sc_hd__inv_2
X_7183_ _7186_/CLK _7183_/D fanout588/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_159_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4395_ _5714_/A0 _4395_/A1 _4399_/S VGND VGND VPWR VPWR _4395_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _7360_/Q _6332_/C _6379_/B1 _7392_/Q VGND VGND VPWR VPWR _6134_/X sky130_fd_sc_hd__a22o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1003 hold2422/X VGND VGND VPWR VPWR hold2423/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _7586_/Q _7587_/Q _6065_/C VGND VGND VPWR VPWR _6065_/Y sky130_fd_sc_hd__nor3_1
Xhold1014 _5750_/X VGND VGND VPWR VPWR _7359_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 hold2770/X VGND VGND VPWR VPWR hold2771/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1036 _5705_/X VGND VGND VPWR VPWR _7319_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 hold2559/X VGND VGND VPWR VPWR hold2560/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1058 hold2572/X VGND VGND VPWR VPWR _7476_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5016_ _4956_/A _5012_/Y _5014_/Y _5011_/Y VGND VGND VPWR VPWR _5016_/Y sky130_fd_sc_hd__o211ai_1
Xhold1069 hold2843/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3824__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6223__A1 _7532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6223__B2 _7484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _7196_/CLK _6967_/D fanout589/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5918_ hold76/X hold61/X _5919_/S VGND VGND VPWR VPWR _5918_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3588__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5982__A0 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6898_ _7075_/CLK _6898_/D _6848_/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5849_ hold464/X _5849_/A1 _5856_/S VGND VGND VPWR VPWR _5849_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5329__A3 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6526__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7519_ _7563_/CLK _7519_/D fanout602/X VGND VGND VPWR VPWR _7519_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3760__A2 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold870 hold870/A VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold881 hold881/A VGND VGND VPWR VPWR hold881/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold892 _5719_/X VGND VGND VPWR VPWR _7332_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5063__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input153_A wb_dat_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2260 _7358_/Q VGND VGND VPWR VPWR hold590/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2271 hold568/X VGND VGND VPWR VPWR _5877_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2282 hold2282/A VGND VGND VPWR VPWR _5673_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2293 _7272_/Q VGND VGND VPWR VPWR hold500/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1570 _7498_/Q VGND VGND VPWR VPWR hold241/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input14_A mask_rev_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1581 hold227/X VGND VGND VPWR VPWR _5890_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1592 hold240/X VGND VGND VPWR VPWR _7377_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_58_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6765__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3579__A2 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6517__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4528__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3751__A2 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6150__B1 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4180_ _5866_/B _5938_/B _4388_/B _4551_/D VGND VGND VPWR VPWR _4190_/S sky130_fd_sc_hd__and4_4
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2216_A _7503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5256__A2 _4744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6453__B2 _7343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6085__B _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6205__A1 _7291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6205__B2 _7347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6821_ _7109_/Q _6821_/A2 _6821_/B1 wire463/A _6820_/X VGND VGND VPWR VPWR _6821_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4216__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6756__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6752_ _6751_/X _6776_/A2 _6777_/S VGND VGND VPWR VPWR _7626_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_70_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3964_ _7431_/Q _3525_/X _3537_/X _7423_/Q _3963_/X VGND VGND VPWR VPWR _3964_/X
+ sky130_fd_sc_hd__a221o_1
X_5703_ _5703_/A0 _5955_/A1 _5703_/S VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6683_ _7057_/Q _6447_/C _6651_/C _6447_/X _7183_/Q VGND VGND VPWR VPWR _6683_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_161_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3895_ _7472_/Q _3494_/X _5857_/A _7456_/Q _3894_/X VGND VGND VPWR VPWR _3895_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5716__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4519__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5634_ _5634_/A _5992_/D VGND VGND VPWR VPWR _5639_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3990__A2 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5565_ _5562_/Y _5564_/Y _5560_/X VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold100 hold100/A VGND VGND VPWR VPWR hold100/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4987__C _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7304_ _7542_/CLK _7304_/D fanout577/X VGND VGND VPWR VPWR _7304_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4516_ _4516_/A0 _5714_/A0 _4520_/S VGND VGND VPWR VPWR _4516_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3742__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold111 hold111/A VGND VGND VPWR VPWR _7531_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold122 hold122/A VGND VGND VPWR VPWR hold122/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold133 _5956_/X VGND VGND VPWR VPWR _5964_/S sky130_fd_sc_hd__buf_4
X_5496_ _5496_/A _5496_/B _5496_/C VGND VGND VPWR VPWR _5529_/C sky130_fd_sc_hd__and3_1
Xhold144 hold144/A VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7235_ _7239_/CLK _7235_/D fanout566/X VGND VGND VPWR VPWR _7235_/Q sky130_fd_sc_hd__dfstp_2
Xhold155 _3468_/X VGND VGND VPWR VPWR _3576_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_4447_ _4447_/A0 hold61/X _4448_/S VGND VGND VPWR VPWR _4447_/X sky130_fd_sc_hd__mux2_1
Xhold166 _7641_/Q VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6141__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold177 hold177/A VGND VGND VPWR VPWR hold177/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold188 hold188/A VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6692__A1 _7123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold199 hold199/A VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout602 fanout606/X VGND VGND VPWR VPWR fanout602/X sky130_fd_sc_hd__buf_12
Xfanout613 input126/X VGND VGND VPWR VPWR _4909_/D sky130_fd_sc_hd__buf_8
XANTENNA__6692__B2 _7158_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7166_ _7213_/CLK _7166_/D fanout590/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfrtp_4
X_4378_ _4378_/A0 _5583_/A0 _4381_/S VGND VGND VPWR VPWR _4378_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_1_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7268_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_input6_A mask_rev_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6116_/B _6097_/B _6144_/B _6116_/X _7311_/Q VGND VGND VPWR VPWR _6117_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout570_A _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7097_ _7197_/CLK _7097_/D fanout601/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5180__A _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6444__A1 _7447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _7594_/Q _7593_/Q _6435_/B VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__a21o_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5707__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3981__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6132__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6683__B2 _7183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2090 _6926_/Q VGND VGND VPWR VPWR hold628/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_59_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6738__A2 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4749__A1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3972__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3680_ _7363_/Q _3564_/X _3648_/X _7040_/Q _3679_/X VGND VGND VPWR VPWR _3680_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5174__A1 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5350_ _5094_/A _5183_/C _4891_/D _5453_/A VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3724__A2 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput205 _4141_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_0_11_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput216 _7655_/X VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
Xoutput227 _7664_/X VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
Xoutput238 _4139_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
X_4301_ _3607_/Y _4301_/A1 _4302_/S VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__mux2_1
Xoutput249 _4133_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
XFILLER_0_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6123__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5281_ _4836_/A _5282_/D _5134_/C _5280_/X VGND VGND VPWR VPWR _5281_/X sky130_fd_sc_hd__a31o_1
XANTENNA_hold2333_A _7307_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7020_ _7170_/CLK _7020_/D fanout573/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_4
X_4232_ _4232_/A0 _4231_/X _4232_/S VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold22_A hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4163_ _7092_/Q _4163_/A1 _7261_/Q VGND VGND VPWR VPWR _4163_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4094_ _4825_/A _5071_/A _4564_/A _4564_/B VGND VGND VPWR VPWR _4095_/D sky130_fd_sc_hd__a211oi_1
XFILLER_0_179_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4328__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6824__A _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6729__A2 _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6804_ _6803_/X _6804_/A1 _6822_/S VGND VGND VPWR VPWR _7638_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5937__A0 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4996_ _4996_/A _5183_/A _5295_/C _5038_/B VGND VGND VPWR VPWR _5033_/D sky130_fd_sc_hd__nand4_1
XANTENNA__5401__A2 _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6735_ _7029_/Q _6459_/B _6459_/C _6451_/X _6877_/Q VGND VGND VPWR VPWR _6735_/X
+ sky130_fd_sc_hd__a32o_1
X_3947_ _7235_/Q _5587_/C _5603_/B _3542_/X _6919_/Q VGND VGND VPWR VPWR _3947_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6666_ _7167_/Q _6408_/D _6657_/X _6662_/X _6665_/X VGND VGND VPWR VPWR _6666_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3963__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3878_ _7037_/Q _3648_/X _3659_/X _7007_/Q _3877_/X VGND VGND VPWR VPWR _3879_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5617_ hold175/X _5896_/A0 _5618_/S VGND VGND VPWR VPWR _5617_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5165__B2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6597_ _6595_/X _6430_/X _6587_/X _6596_/X VGND VGND VPWR VPWR _6597_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3715__A2 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5548_ _5548_/A _5548_/B _5575_/B VGND VGND VPWR VPWR _5548_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6114__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5479_ _4679_/Y _4814_/Y _4971_/X _5478_/Y VGND VGND VPWR VPWR _5482_/B sky130_fd_sc_hd__o31a_1
XANTENNA__6665__A1 _7001_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7218_ _4150_/A1 _7218_/D _6870_/X VGND VGND VPWR VPWR _7218_/Q sky130_fd_sc_hd__dfrtn_1
Xfanout410 _4491_/A VGND VGND VPWR VPWR _5612_/C sky130_fd_sc_hd__buf_12
Xfanout421 hold35/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__buf_12
Xfanout432 _6404_/Y VGND VGND VPWR VPWR _6651_/B sky130_fd_sc_hd__clkbuf_16
Xfanout443 _6035_/Y VGND VGND VPWR VPWR _6144_/B sky130_fd_sc_hd__buf_12
X_7149_ _7447_/CLK _7149_/D fanout598/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3423__A _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout465 hold17/X VGND VGND VPWR VPWR _5955_/A1 sky130_fd_sc_hd__buf_12
Xfanout476 _5979_/A0 VGND VGND VPWR VPWR _5586_/A0 sky130_fd_sc_hd__clkbuf_16
Xfanout487 _5986_/A1 VGND VGND VPWR VPWR _5914_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout498 _5840_/A1 VGND VGND VPWR VPWR _5993_/A1 sky130_fd_sc_hd__buf_12
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7190__RESET_B fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A wb_adr_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5928__A0 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5069__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5784__S hold49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3954__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input81_A spi_sdo VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4701__B _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5459__A2 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3890__A1 _7178_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7207__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_185_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4850_ _5295_/D _4850_/B _5138_/D _5295_/A VGND VGND VPWR VPWR _5294_/C sky130_fd_sc_hd__nand4_4
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6082__C _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6187__A3 _6093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3801_ _3485_/X _4491_/A _3931_/D _3501_/X _7577_/Q VGND VGND VPWR VPWR _3801_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_185_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4781_ _4781_/A _4781_/B VGND VGND VPWR VPWR _4781_/Y sky130_fd_sc_hd__nor2_1
X_6520_ _7409_/Q _6468_/X _6430_/X _6519_/X _6516_/X VGND VGND VPWR VPWR _6520_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3945__A2 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3732_ _3732_/A _3732_/B _3732_/C _3732_/D VGND VGND VPWR VPWR _3733_/D sky130_fd_sc_hd__nor4_2
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6451_ _7595_/Q _6467_/A _6600_/B _7596_/Q VGND VGND VPWR VPWR _6451_/X sky130_fd_sc_hd__and4b_4
XFILLER_0_113_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6344__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3663_ _4509_/A _4551_/C _3931_/D VGND VGND VPWR VPWR _3663_/X sky130_fd_sc_hd__and3_2
XFILLER_0_43_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2450_A _7315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3508__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5402_ _5374_/X _5401_/X _5580_/A2 _5372_/X VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__a211o_1
X_6382_ _7116_/Q _6317_/C _6089_/X _7045_/Q _6381_/X VGND VGND VPWR VPWR _6382_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3594_ _7397_/Q _5803_/A _3933_/A _3519_/X _7549_/Q VGND VGND VPWR VPWR _3594_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5333_ _5053_/C _5553_/A1 _5328_/X _5332_/X VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_140_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5264_ _4786_/C _5079_/B _5102_/B _5263_/X VGND VGND VPWR VPWR _5265_/D sky130_fd_sc_hd__a31oi_2
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2804 hold2804/A VGND VGND VPWR VPWR _4480_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7003_ _7144_/CLK _7003_/D fanout572/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfstp_2
Xhold2815 _6982_/Q VGND VGND VPWR VPWR _4294_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2826 hold2826/A VGND VGND VPWR VPWR _4433_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4215_ _4078_/A _4078_/B _4168_/D _5785_/B _5992_/C VGND VGND VPWR VPWR _4215_/X
+ sky130_fd_sc_hd__o311a_2
Xhold2837 _6983_/Q VGND VGND VPWR VPWR _4296_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2848 hold2848/A VGND VGND VPWR VPWR hold2848/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5195_ _4672_/X _5174_/Y _4986_/Y _5169_/X _5194_/Y VGND VGND VPWR VPWR _5195_/X
+ sky130_fd_sc_hd__o311a_1
Xhold2859 _5813_/X VGND VGND VPWR VPWR hold2859/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4146_ _7265_/Q input80/X _4174_/B VGND VGND VPWR VPWR _4146_/X sky130_fd_sc_hd__mux2_8
X_4077_ _3400_/Y _4076_/C _4076_/X VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__o21bai_1
XANTENNA__5083__B1 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5622__A2 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3633__A1 _7484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3633__B2 _7444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5386__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4979_ _4996_/A _5328_/A _5328_/B VGND VGND VPWR VPWR _5034_/C sky130_fd_sc_hd__and3_2
XANTENNA__6583__B1 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6718_ _7184_/Q _6574_/B _6771_/A3 _6443_/X _7194_/Q VGND VGND VPWR VPWR _6718_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3936__A2 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6649_ _6648_/X _6649_/A1 _6649_/S VGND VGND VPWR VPWR _6649_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6335__B1 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4521__B _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3418__A _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6350__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5310__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5310__B2 _4744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_csclk _7496_/CLK VGND VGND VPWR VPWR _7429_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__7371__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5779__S hold49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6326__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3560__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6629__A1 _7542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6629__B2 _7518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7459__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4159__A input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4000_ _4002_/B _4006_/A _6910_/Q VGND VGND VPWR VPWR _4003_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5951_ _5951_/A0 _5951_/A1 _5955_/S VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3615__A1 _7292_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4606__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3615__B2 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5080__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4902_ _4902_/A _4902_/B _5448_/D _5223_/D VGND VGND VPWR VPWR _4904_/B sky130_fd_sc_hd__nand4_1
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5882_ _5882_/A0 _5954_/A1 _5883_/S VGND VGND VPWR VPWR _5882_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_192_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7621_ _7621_/CLK _7621_/D fanout579/X VGND VGND VPWR VPWR _7621_/Q sky130_fd_sc_hd__dfrtp_1
X_4833_ _5295_/D _4834_/B _5295_/A VGND VGND VPWR VPWR _4839_/B sky130_fd_sc_hd__and3_1
XFILLER_0_145_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6565__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3918__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7552_ _7581_/CLK _7552_/D fanout584/X VGND VGND VPWR VPWR _7552_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_145_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4764_ _4700_/Y _4727_/Y _4718_/Y _4763_/Y VGND VGND VPWR VPWR _4766_/B sky130_fd_sc_hd__o211ai_1
XFILLER_0_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6503_ _7353_/Q _6413_/C _6459_/C _6408_/B _7377_/Q VGND VGND VPWR VPWR _6503_/X
+ sky130_fd_sc_hd__a32o_1
X_3715_ _6915_/Q _5612_/B _5947_/A _3515_/X _7239_/Q VGND VGND VPWR VPWR _3715_/X
+ sky130_fd_sc_hd__a32o_2
X_7483_ _7521_/CLK _7483_/D fanout600/X VGND VGND VPWR VPWR _7483_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4695_ _4802_/A _4794_/A VGND VGND VPWR VPWR _4695_/Y sky130_fd_sc_hd__nand2_2
XANTENNA_hold2832_A _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6434_ _6455_/B _6434_/B _6600_/B VGND VGND VPWR VPWR _6434_/X sky130_fd_sc_hd__and3_4
XFILLER_0_125_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3646_ _4449_/B _5612_/C _4346_/C VGND VGND VPWR VPWR _4322_/A sky130_fd_sc_hd__and3_4
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6365_ _7195_/Q _6072_/B _6120_/B _6364_/X VGND VGND VPWR VPWR _6365_/X sky130_fd_sc_hd__a31o_1
X_3577_ _4388_/B _5596_/B _5640_/C VGND VGND VPWR VPWR _5630_/S sky130_fd_sc_hd__and3_1
XFILLER_0_140_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4995__C _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3551__B1 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5316_ _4605_/Y _4956_/A _4731_/Y _4755_/Y _4814_/Y VGND VGND VPWR VPWR _5531_/A
+ sky130_fd_sc_hd__o32a_1
X_6296_ _7177_/Q _6092_/X _6295_/X _6294_/X _6293_/X VGND VGND VPWR VPWR _6303_/A
+ sky130_fd_sc_hd__a2111o_1
Xhold2601 _7241_/Q VGND VGND VPWR VPWR hold845/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2612 _5729_/X VGND VGND VPWR VPWR hold877/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__A2 _6090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7129__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5247_ _5419_/A _5247_/B _5247_/C VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__and3_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout483_A _5735_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2623 hold879/X VGND VGND VPWR VPWR _4218_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2634 hold626/X VGND VGND VPWR VPWR _5648_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1900 _5707_/X VGND VGND VPWR VPWR hold433/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2645 _5961_/X VGND VGND VPWR VPWR hold681/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__buf_4
Xhold1911 _7231_/Q VGND VGND VPWR VPWR hold520/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2656 _6971_/Q VGND VGND VPWR VPWR hold753/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1922 _5593_/X VGND VGND VPWR VPWR hold546/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_leaf_46_csclk_A _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2667 _7035_/Q VGND VGND VPWR VPWR hold747/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__clkbuf_16
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1933 hold406/X VGND VGND VPWR VPWR _4549_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5178_ _5295_/C _5183_/C _5216_/A VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__o21a_1
Xhold2678 hold881/X VGND VGND VPWR VPWR _4237_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1944 hold428/X VGND VGND VPWR VPWR _5852_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2689 _7196_/Q VGND VGND VPWR VPWR hold763/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1955 _4362_/X VGND VGND VPWR VPWR hold447/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1966 _5806_/X VGND VGND VPWR VPWR hold519/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4129_ _6897_/Q _4129_/B VGND VGND VPWR VPWR _4130_/A sky130_fd_sc_hd__nand2b_2
Xhold1977 hold488/X VGND VGND VPWR VPWR _4262_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1988 _7018_/Q VGND VGND VPWR VPWR hold572/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1999 _7434_/Q VGND VGND VPWR VPWR hold440/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_39_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6556__B1 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1765_A hold284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3909__A2 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6308__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6323__A3 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input44_A mgmt_gpio_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5598__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4426__B _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4270__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6547__B1 _6545_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5770__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5972__S hold13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3500_ _3511_/A hold53/X _3500_/C VGND VGND VPWR VPWR _3519_/B sky130_fd_sc_hd__and3_4
XFILLER_0_107_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_170_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4480_ _4480_/A0 _5840_/A1 _4484_/S VGND VGND VPWR VPWR _4480_/X sky130_fd_sc_hd__mux2_1
Xhold507 hold507/A VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold518 hold518/A VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold529 _3453_/X VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3431_ _7394_/Q VGND VGND VPWR VPWR _3431_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_150_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3533__B1 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3679__A4 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6150_ _7513_/Q _7592_/Q _6317_/C _6087_/X _7465_/Q VGND VGND VPWR VPWR _6150_/X
+ sky130_fd_sc_hd__a32o_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _4888_/B _5091_/A _5100_/X _5099_/Y VGND VGND VPWR VPWR _5101_/Y sky130_fd_sc_hd__a31oi_2
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7589_/Q _6119_/A _6106_/B _7588_/Q VGND VGND VPWR VPWR _6081_/X sky130_fd_sc_hd__and4bb_4
XFILLER_0_148_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 hold2869/X VGND VGND VPWR VPWR hold1207/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _4984_/B _4984_/A _4660_/Y _4862_/X _4759_/Y VGND VGND VPWR VPWR _5033_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 hold2755/X VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1229 hold3050/X VGND VGND VPWR VPWR hold3051/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_164_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3521__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_178_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5589__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6983_ _7633_/CLK _6983_/D VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5934_ _5997_/A1 _5934_/A1 _5937_/S VGND VGND VPWR VPWR _5934_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4261__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5865_ _5991_/A1 _5865_/A1 _5865_/S VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6538__B1 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7604_ _7623_/CLK _7604_/D fanout576/X VGND VGND VPWR VPWR _7604_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4816_ _5410_/A _5061_/B _5399_/C VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__and3_1
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5796_ _5967_/A1 _5796_/A1 _5802_/S VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4747_ _4887_/D _4747_/B _4887_/B _4879_/C VGND VGND VPWR VPWR _5094_/A sky130_fd_sc_hd__and4b_4
X_7535_ _7537_/CLK _7535_/D fanout577/X VGND VGND VPWR VPWR _7535_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5882__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7466_ _7530_/CLK _7466_/D fanout600/X VGND VGND VPWR VPWR _7466_/Q sky130_fd_sc_hd__dfrtp_4
X_4678_ _4679_/A _5089_/C _4679_/C VGND VGND VPWR VPWR _5342_/A sky130_fd_sc_hd__and3_4
XFILLER_0_98_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6417_ _6427_/A _6434_/B _6747_/C VGND VGND VPWR VPWR _6419_/C sky130_fd_sc_hd__and3_4
X_3629_ _7412_/Q _3493_/X _5686_/A _7308_/Q _3628_/X VGND VGND VPWR VPWR _3632_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4316__A2 _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5513__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6710__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7397_ _7581_/CLK _7397_/D fanout584/X VGND VGND VPWR VPWR _7397_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5614__C hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6348_ _7211_/Q _6332_/B _6089_/X _6100_/X _7063_/Q VGND VGND VPWR VPWR _6348_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3110 _5966_/X VGND VGND VPWR VPWR hold3110/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3121 _5822_/X VGND VGND VPWR VPWR hold3121/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3132 _5630_/X VGND VGND VPWR VPWR hold3132/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6069__A2 _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3143 _4383_/X VGND VGND VPWR VPWR hold3143/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4563_/C sky130_fd_sc_hd__clkbuf_2
X_6279_ _7350_/Q _6070_/X _6082_/X _7326_/Q _6278_/X VGND VGND VPWR VPWR _6280_/D
+ sky130_fd_sc_hd__a221o_1
Xhold3154 _5876_/X VGND VGND VPWR VPWR hold3154/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2420 _7119_/Q VGND VGND VPWR VPWR hold941/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3165 hold3165/A VGND VGND VPWR VPWR _5732_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR _4831_/A sky130_fd_sc_hd__clkbuf_4
Xhold2431 _7024_/Q VGND VGND VPWR VPWR hold951/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3176 _7215_/Q VGND VGND VPWR VPWR _3924_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5277__B1 _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5911__A _5911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6820_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2442 hold997/X VGND VGND VPWR VPWR _5701_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3187 _6792_/S VGND VGND VPWR VPWR _6789_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6802_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3198 _7641_/Q VGND VGND VPWR VPWR _6813_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2453 hold649/X VGND VGND VPWR VPWR _5629_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2464 _7251_/Q VGND VGND VPWR VPWR hold2464/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1730 _7276_/Q VGND VGND VPWR VPWR hold316/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2475 _7048_/Q VGND VGND VPWR VPWR hold905/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1741 _5870_/X VGND VGND VPWR VPWR hold238/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2486 hold949/X VGND VGND VPWR VPWR _5647_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1752 _7368_/Q VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2497 _7148_/Q VGND VGND VPWR VPWR hold670/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1763 _5960_/X VGND VGND VPWR VPWR hold303/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1774 hold334/X VGND VGND VPWR VPWR _5789_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3431__A _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1785 _7561_/Q VGND VGND VPWR VPWR hold308/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1796 _5969_/X VGND VGND VPWR VPWR hold365/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6241__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4252__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5752__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5792__S _5793_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3763__B1 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4840__A_N _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5821__A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6480__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6768__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5967__S hold13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6232__A2 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3980_ _7036_/Q _3648_/X _4545_/A _7192_/Q _3927_/X VGND VGND VPWR VPWR _3980_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3597__A3 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5991__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5650_ _7257_/Q hold284/X _4168_/D _4248_/S hold47/X VGND VGND VPWR VPWR _5653_/S
+ sky130_fd_sc_hd__o311ai_4
XFILLER_0_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6090__C _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4601_ _5091_/A _5399_/A VGND VGND VPWR VPWR _4601_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5743__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5581_ _5581_/A _5902_/B VGND VGND VPWR VPWR _5586_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_127_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7320_ _7499_/CLK _7320_/D fanout578/X VGND VGND VPWR VPWR _7320_/Q sky130_fd_sc_hd__dfstp_4
X_4532_ _4532_/A0 hold84/X _4532_/S VGND VGND VPWR VPWR _4532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold304 hold304/A VGND VGND VPWR VPWR hold304/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7251_ _7264_/CLK _7251_/D fanout565/X VGND VGND VPWR VPWR _7251_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6299__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7403__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold315 _4356_/X VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold326 hold326/A VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4463_ _4463_/A0 _5583_/A0 _4466_/S VGND VGND VPWR VPWR _4463_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold337 hold337/A VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold348 hold348/A VGND VGND VPWR VPWR hold348/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6202_ _7523_/Q _6379_/B1 _6200_/X _6201_/X VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3516__A hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3414_ _7530_/Q VGND VGND VPWR VPWR _3414_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold359 hold359/A VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7182_ _7186_/CLK _7182_/D fanout588/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_4
X_4394_ _4394_/A _5902_/B VGND VGND VPWR VPWR _4399_/S sky130_fd_sc_hd__nand2_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6133_ _6094_/A _6130_/X _6132_/X _6126_/X _6128_/X VGND VGND VPWR VPWR _6133_/X
+ sky130_fd_sc_hd__a2111o_4
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5731__A _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 _5737_/X VGND VGND VPWR VPWR _7348_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6064_ _6064_/A1 _6062_/X _6063_/X VGND VGND VPWR VPWR _7600_/D sky130_fd_sc_hd__a21bo_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 hold2464/X VGND VGND VPWR VPWR hold2465/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1026 _4272_/X VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1037 hold2734/X VGND VGND VPWR VPWR hold2735/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5015_ _5038_/A _5553_/A1 _5030_/C _5013_/X VGND VGND VPWR VPWR _5015_/X sky130_fd_sc_hd__a31o_1
Xhold1048 _5746_/X VGND VGND VPWR VPWR _7356_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1059 hold2591/X VGND VGND VPWR VPWR hold2592/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4482__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6759__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5877__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6223__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4234__A1 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A _6022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6966_ _7070_/CLK _6966_/D fanout590/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5431__B1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5917_ _5917_/A0 _5998_/A1 _5919_/S VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3588__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6897_ _7075_/CLK _6897_/D _6847_/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3993__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5848_ _5848_/A hold48/X VGND VGND VPWR VPWR _5856_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_146_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5734__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5779_ _5896_/A0 _5779_/A1 hold49/X VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7518_ _7565_/CLK _7518_/D fanout603/X VGND VGND VPWR VPWR _7518_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7449_ _7505_/CLK _7449_/D fanout601/X VGND VGND VPWR VPWR _7449_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3760__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold860 hold860/A VGND VGND VPWR VPWR hold860/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold871 hold871/A VGND VGND VPWR VPWR _7477_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold882 hold882/A VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold893 hold893/A VGND VGND VPWR VPWR hold893/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input146_A wb_dat_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2250 hold472/X VGND VGND VPWR VPWR _5616_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6907__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2261 hold590/X VGND VGND VPWR VPWR _5748_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2272 _5877_/X VGND VGND VPWR VPWR hold569/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2283 _7430_/Q VGND VGND VPWR VPWR hold580/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2294 hold500/X VGND VGND VPWR VPWR _5652_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5670__A0 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1560 hold223/X VGND VGND VPWR VPWR _5635_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1571 hold241/X VGND VGND VPWR VPWR _5906_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1582 _7203_/Q VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1593 _7063_/Q VGND VGND VPWR VPWR hold298/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5787__S _5793_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4225__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3579__A3 _3578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5973__A1 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3984__B1 _3675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6517__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5725__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3751__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6150__A1 _7513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6150__B2 _7465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6453__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6085__C _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4464__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6205__A2 _6072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__A3 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6820_ _7111_/Q _6820_/A2 _6820_/B1 _7110_/Q VGND VGND VPWR VPWR _6820_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4736__A_N _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4216__A1 _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6756__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6751_ _6750_/X _6751_/A1 _6751_/S VGND VGND VPWR VPWR _6751_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5964__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3963_ _7257_/Q _5965_/A _5632_/B _3669_/X _6967_/Q VGND VGND VPWR VPWR _3963_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_163_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5702_ _5702_/A0 _5954_/A1 _5703_/S VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__mux2_1
X_6682_ _7128_/Q _6424_/X _6677_/X _6681_/X _6430_/X VGND VGND VPWR VPWR _6682_/X
+ sky130_fd_sc_hd__a2111o_1
X_3894_ _7057_/Q _5938_/C _4521_/B _3663_/X _7163_/Q VGND VGND VPWR VPWR _3894_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__6508__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5633_ _5633_/A0 _5993_/A1 _5633_/S VGND VGND VPWR VPWR _5633_/X sky130_fd_sc_hd__mux2_1
X_5564_ _5564_/A _5564_/B _5564_/C VGND VGND VPWR VPWR _5564_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_41_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold101 hold101/A VGND VGND VPWR VPWR _7283_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7303_ _7309_/CLK _7303_/D fanout576/X VGND VGND VPWR VPWR _7303_/Q sky130_fd_sc_hd__dfstp_4
X_4515_ _5938_/B _4551_/C hold56/A _4551_/D VGND VGND VPWR VPWR _4520_/S sky130_fd_sc_hd__and4_4
Xhold112 hold112/A VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold123 hold123/A VGND VGND VPWR VPWR _7445_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3742__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5495_ _4956_/A _4956_/B _4595_/Y _4605_/Y VGND VGND VPWR VPWR _5529_/B sky130_fd_sc_hd__a211o_1
Xhold134 hold134/A VGND VGND VPWR VPWR _7549_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold145 hold145/A VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4446_ _4446_/A0 _5998_/A1 _4448_/S VGND VGND VPWR VPWR _4446_/X sky130_fd_sc_hd__mux2_1
X_7234_ _7255_/CLK _7234_/D fanout565/X VGND VGND VPWR VPWR _7234_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6141__A1 _7512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold156 _4455_/X VGND VGND VPWR VPWR _4460_/S sky130_fd_sc_hd__buf_2
Xhold167 hold167/A VGND VGND VPWR VPWR hold167/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold178 hold178/A VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4152__A0 _6947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold189 hold189/A VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout603 fanout605/X VGND VGND VPWR VPWR fanout603/X sky130_fd_sc_hd__buf_12
X_7165_ _7170_/CLK _7165_/D fanout573/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6692__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout614 _4786_/C VGND VGND VPWR VPWR _4805_/B sky130_fd_sc_hd__buf_12
X_4377_ _4377_/A0 _5840_/A1 _4381_/S VGND VGND VPWR VPWR _4377_/X sky130_fd_sc_hd__mux2_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6116_/A _6116_/B _6116_/C VGND VGND VPWR VPWR _6116_/X sky130_fd_sc_hd__and3_4
X_7096_ _7096_/CLK _7096_/D fanout605/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5180__B _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6047_ _6435_/B _6434_/B VGND VGND VPWR VPWR _6047_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6444__A2 _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5652__A0 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4207__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5955__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6949_ _6956_/CLK _6949_/D fanout604/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1580_A _7484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3966__B1 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3981__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1845_A _7465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4391__A0 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5074__C _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6132__B2 _7504_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4143__B1 _4142_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6683__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold690 hold690/A VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6467__A _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4446__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2080 _5636_/X VGND VGND VPWR VPWR hold109/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_188_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2091 hold628/X VGND VGND VPWR VPWR _4211_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1390 _6887_/Q VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6199__A1 _7483_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4715__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5946__A1 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7066__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3972__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6371__A1 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6371__B2 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput206 _3405_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
XFILLER_0_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput217 _4165_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
X_4300_ _3643_/Y _4300_/A1 _4302_/S VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__mux2_1
Xoutput228 _7665_/X VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
Xoutput239 _4138_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
XANTENNA__6123__A1 _7279_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5280_ _4836_/A _5061_/B _5399_/C _5279_/Y VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4231_ _4258_/A0 _5991_/A1 _4231_/S VGND VGND VPWR VPWR _4231_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6674__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4162_ _6939_/Q _4164_/A1 _7258_/Q VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
X_4093_ _4093_/A _4093_/B _4093_/C _4093_/D VGND VGND VPWR VPWR _4096_/C sky130_fd_sc_hd__and4_1
XANTENNA__4437__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4328__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2695_A _7483_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6729__A3 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6803_ _7110_/Q _6803_/A2 _6803_/B1 _4426_/Y _6802_/X VGND VGND VPWR VPWR _6803_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4995_ _4996_/A _5183_/A _5138_/D _5038_/B VGND VGND VPWR VPWR _5033_/C sky130_fd_sc_hd__nand4_1
XFILLER_0_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6734_ _7054_/Q _6434_/B _6771_/A3 _6420_/C _7125_/Q VGND VGND VPWR VPWR _6734_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3946_ _7295_/Q hold12/A _4346_/C _3666_/X _7011_/Q VGND VGND VPWR VPWR _3946_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3877_ _7027_/Q _4346_/C _5603_/B _3543_/X _7288_/Q VGND VGND VPWR VPWR _3877_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3963__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6665_ _7001_/Q _6419_/D _6424_/X _7127_/Q _6664_/X VGND VGND VPWR VPWR _6665_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5616_ _5616_/A0 _5967_/A1 _5618_/S VGND VGND VPWR VPWR _5616_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5165__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6596_ _7284_/Q _6431_/Y _6775_/B1 VGND VGND VPWR VPWR _6596_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout409_A _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4373__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5547_ _4741_/Y _5065_/Y _5352_/Y _5448_/B _5546_/X VGND VGND VPWR VPWR _5575_/B
+ sky130_fd_sc_hd__o2111a_2
XANTENNA__3715__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7671__A _7671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5478_ _5478_/A _5478_/B _5559_/B VGND VGND VPWR VPWR _5478_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4125__A0 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4429_ _4114_/B _4429_/B VGND VGND VPWR VPWR _4430_/D sky130_fd_sc_hd__nand2b_1
X_7217_ _7075_/CLK _7217_/D _6869_/X VGND VGND VPWR VPWR _7217_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__6665__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3479__A2 _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout411 _4491_/A VGND VGND VPWR VPWR _4551_/C sky130_fd_sc_hd__buf_12
Xfanout422 _6106_/X VGND VGND VPWR VPWR _6379_/B1 sky130_fd_sc_hd__buf_12
XFILLER_0_10_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout433 _6404_/Y VGND VGND VPWR VPWR _6413_/C sky130_fd_sc_hd__buf_4
Xfanout444 _6023_/Y VGND VGND VPWR VPWR _6116_/C sky130_fd_sc_hd__buf_12
X_7148_ _7395_/CLK _7148_/D fanout598/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout466 hold17/X VGND VGND VPWR VPWR _5991_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout477 _5979_/A0 VGND VGND VPWR VPWR _5997_/A1 sky130_fd_sc_hd__buf_12
X_7079_ _7096_/CLK _7079_/D fanout605/X VGND VGND VPWR VPWR _7659_/A sky130_fd_sc_hd__dfrtp_1
Xfanout488 _5995_/A1 VGND VGND VPWR VPWR _5986_/A1 sky130_fd_sc_hd__buf_12
Xfanout499 hold464/X VGND VGND VPWR VPWR _5840_/A1 sky130_fd_sc_hd__buf_12
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7506__RESET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input109_A wb_adr_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input74_A pad_flash_io1_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6105__A1 _7303_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6105__B2 _7287_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6656__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4429__B _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3890__A2 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5919__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ _7139_/Q _5965_/A _4521_/B _3798_/X VGND VGND VPWR VPWR _3800_/X sky130_fd_sc_hd__a31o_4
X_4780_ _5091_/C _5387_/C _4790_/B VGND VGND VPWR VPWR _4781_/A sky130_fd_sc_hd__and3_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__A1 _7468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5395__A2 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__B2 _7508_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3731_ _4177_/B _4231_/S _3727_/X _3729_/X _3730_/X VGND VGND VPWR VPWR _3732_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_184_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_0_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7189_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4180__A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3662_ _4509_/A _5640_/B _5612_/C VGND VGND VPWR VPWR _4394_/A sky130_fd_sc_hd__and3_4
X_6450_ _7559_/Q _6419_/C _6442_/X _6445_/X _6449_/X VGND VGND VPWR VPWR _6471_/A
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5147__A2 _4758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6344__B2 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5001__D1 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5401_ _4836_/A _5399_/A _5401_/A3 _5400_/Y VGND VGND VPWR VPWR _5401_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6381_ _6966_/Q _6072_/B _6144_/B _6332_/C _7035_/Q VGND VGND VPWR VPWR _6381_/X
+ sky130_fd_sc_hd__a32o_1
X_3593_ _7413_/Q _5803_/A _3590_/C _5713_/A _7333_/Q VGND VGND VPWR VPWR _3593_/X
+ sky130_fd_sc_hd__a32o_1
X_5332_ _5339_/A _5011_/A _5339_/B _5331_/Y VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5263_ _5222_/A _5260_/C _5387_/D _4756_/X VGND VGND VPWR VPWR _5263_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_11_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5855__A0 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2805 _6998_/Q VGND VGND VPWR VPWR _4319_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_167_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4214_ _4214_/A0 _5805_/A1 _4214_/S VGND VGND VPWR VPWR _4214_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7002_ _7212_/CLK _7002_/D fanout574/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2816 hold2816/A VGND VGND VPWR VPWR hold2816/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5194_ _5183_/A _5188_/X _5203_/B _5170_/X _5193_/X VGND VGND VPWR VPWR _5194_/Y
+ sky130_fd_sc_hd__a311oi_2
Xhold2827 _6975_/Q VGND VGND VPWR VPWR _4283_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2838 hold2838/A VGND VGND VPWR VPWR hold2838/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2849 _6996_/Q VGND VGND VPWR VPWR _4315_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4145_ _7562_/Q _4174_/B _4144_/Y VGND VGND VPWR VPWR _4145_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3881__A2 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4076_ _6909_/Q _4076_/B _4076_/C _6910_/Q VGND VGND VPWR VPWR _4076_/X sky130_fd_sc_hd__and4b_1
XANTENNA__5083__A1 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3633__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5386__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6583__A1 _7436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4978_ _5410_/A _5138_/D VGND VGND VPWR VPWR _4978_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_19_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6583__B2 _7556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6717_ _7159_/Q _6419_/A _6419_/C _7139_/Q _6716_/X VGND VGND VPWR VPWR _6717_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3929_ _3929_/A VGND VGND VPWR VPWR _3929_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3936__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6648_ _6631_/Y wire347/X _7286_/Q _6431_/Y VGND VGND VPWR VPWR _6648_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__6335__B2 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4521__C _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6579_ _7372_/Q _6413_/C _6651_/C _6058_/X _7532_/Q VGND VGND VPWR VPWR _6579_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6638__A2 _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3434__A _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3872__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6271__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4265__A _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3624__A2 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5795__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6629__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6262__B1 _6093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4175__A _4175_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5950_ _5950_/A0 _5950_/A1 _5955_/S VGND VGND VPWR VPWR _5950_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6093__C _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3615__A2 _3543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4901_ _4726_/Y _4899_/Y _4898_/Y _4894_/Y _4891_/Y VGND VGND VPWR VPWR _4902_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5881_ _5881_/A0 _5953_/A1 _5883_/S VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7620_ _7621_/CLK _7620_/D fanout582/X VGND VGND VPWR VPWR _7620_/Q sky130_fd_sc_hd__dfrtp_1
X_4832_ _5260_/B _4836_/C VGND VGND VPWR VPWR _4832_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6565__A1 _7307_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6565__B2 _7291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7551_ _7551_/CLK _7551_/D fanout595/X VGND VGND VPWR VPWR _7551_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_172_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4763_ _4763_/A _4763_/B _4763_/C VGND VGND VPWR VPWR _4763_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__3918__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3519__A hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2658_A _7448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6502_ _7401_/Q _6409_/X _6420_/B _7305_/Q _6499_/X VGND VGND VPWR VPWR _6502_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3714_ _6966_/Q _5632_/B _5659_/B _3663_/X _7166_/Q VGND VGND VPWR VPWR _3714_/X
+ sky130_fd_sc_hd__a32o_2
X_7482_ _7565_/CLK _7482_/D fanout605/X VGND VGND VPWR VPWR _7482_/Q sky130_fd_sc_hd__dfrtp_4
X_4694_ _4768_/B _4694_/B _4801_/B _4801_/C VGND VGND VPWR VPWR _5138_/C sky130_fd_sc_hd__nor4_4
XFILLER_0_126_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6433_ _6462_/D _7598_/Q _7597_/Q _6435_/B VGND VGND VPWR VPWR _6574_/C sky130_fd_sc_hd__and4bb_4
X_3645_ _3644_/X _3645_/A1 _3996_/A VGND VGND VPWR VPWR _3645_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6364_ _7212_/Q _6089_/X _6379_/B1 _7190_/Q _6363_/X VGND VGND VPWR VPWR _6364_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3576_ _4491_/C _3576_/B _3576_/C VGND VGND VPWR VPWR _3576_/X sky130_fd_sc_hd__and3_4
XANTENNA__3551__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3551__B2 _7518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5315_ _5038_/A _5410_/A _4823_/B _4809_/B _5160_/C VGND VGND VPWR VPWR _5317_/C
+ sky130_fd_sc_hd__a311o_1
X_6295_ _7142_/Q _6121_/C _6116_/C _6136_/C VGND VGND VPWR VPWR _6295_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2602 hold845/X VGND VGND VPWR VPWR _5610_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2613 _7413_/Q VGND VGND VPWR VPWR hold872/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5246_ _4622_/Y _4726_/Y _4748_/Y _4947_/Y _5245_/X VGND VGND VPWR VPWR _5247_/C
+ sky130_fd_sc_hd__o32a_1
Xhold2624 _4218_/X VGND VGND VPWR VPWR hold880/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2635 _7381_/Q VGND VGND VPWR VPWR hold862/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1901 _7354_/Q VGND VGND VPWR VPWR hold292/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4500__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2646 _7579_/Q VGND VGND VPWR VPWR hold651/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1912 hold520/X VGND VGND VPWR VPWR _5599_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5177_ _5295_/C _5183_/C _5553_/A1 VGND VGND VPWR VPWR _5177_/Y sky130_fd_sc_hd__o21ai_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__buf_6
Xhold2657 hold753/X VGND VGND VPWR VPWR _4276_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1923 _6913_/Q VGND VGND VPWR VPWR hold524/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2668 hold747/X VGND VGND VPWR VPWR _4363_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout476_A _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2679 _4237_/X VGND VGND VPWR VPWR hold882/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1934 _4549_/X VGND VGND VPWR VPWR hold407/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1945 _5852_/X VGND VGND VPWR VPWR hold429/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4128_ _6896_/Q _4128_/B VGND VGND VPWR VPWR _4128_/Y sky130_fd_sc_hd__nor2_1
Xhold1956 hold447/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1967 hold519/X VGND VGND VPWR VPWR _7409_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1978 _4262_/X VGND VGND VPWR VPWR hold489/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1989 hold572/X VGND VGND VPWR VPWR _4343_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6253__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4059_ _6892_/Q _6891_/Q _4123_/B _4058_/Y VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3909__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3429__A _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4319__A0 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6459__B _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6492__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input37_A mgmt_gpio_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3845__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6244__B1 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4426__C _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4723__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3781__A1 _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5507__C1 _5185_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold508 hold508/A VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold519 hold519/A VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3430_ _7402_/Q VGND VGND VPWR VPWR _3430_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3533__A1 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5100_/A _5260_/B _5387_/C VGND VGND VPWR VPWR _5100_/X sky130_fd_sc_hd__and3_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _6094_/A _6136_/B _6116_/A VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__and3_4
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5031_/B _5031_/C VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__nor3_1
XANTENNA__6483__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 hold1208/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
Xhold1219 hold3014/X VGND VGND VPWR VPWR hold3015/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3836__A2 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2406_A _7441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6235__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3521__B _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6982_ _7633_/CLK _6982_/D VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5933_ _5996_/A1 _5933_/A1 _5937_/S VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6250__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_csclk _7267_/CLK VGND VGND VPWR VPWR _7522_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_180_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5864_ _5999_/A1 _5864_/A1 _5865_/S VGND VGND VPWR VPWR _5864_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6538__A1 _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6538__B2 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4549__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7603_ _7623_/CLK _7603_/D fanout575/X VGND VGND VPWR VPWR _7603_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4815_ _5387_/C _4815_/B _5399_/C VGND VGND VPWR VPWR _4818_/A sky130_fd_sc_hd__and3_1
XANTENNA__4352__B _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5210__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5795_ _5903_/A0 _5795_/A1 _5802_/S VGND VGND VPWR VPWR _5795_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_133_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7534_ _7566_/CLK _7534_/D fanout596/X VGND VGND VPWR VPWR _7534_/Q sky130_fd_sc_hd__dfrtp_4
X_4746_ _4755_/A _5138_/B _4746_/C _5005_/A VGND VGND VPWR VPWR _4746_/Y sky130_fd_sc_hd__nand4_1
Xclkbuf_leaf_48_csclk _7496_/CLK VGND VGND VPWR VPWR _7577_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7465_ _7563_/CLK _7465_/D fanout602/X VGND VGND VPWR VPWR _7465_/Q sky130_fd_sc_hd__dfrtp_4
X_4677_ _5089_/B _4675_/Y _4673_/Y _4562_/Y VGND VGND VPWR VPWR _4758_/B sky130_fd_sc_hd__o2bb2ai_4
X_6416_ _6435_/B _6467_/A _6651_/B _6462_/D VGND VGND VPWR VPWR _6419_/B sky130_fd_sc_hd__and4bb_1
X_3628_ _7540_/Q _3590_/C _5947_/B _3544_/X _7420_/Q VGND VGND VPWR VPWR _3628_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7396_ _7581_/CLK _7396_/D fanout584/X VGND VGND VPWR VPWR _7396_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_114_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6347_ _7053_/Q _6087_/X _6344_/X _6346_/X VGND VGND VPWR VPWR _6347_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3559_ _7542_/Q _5947_/A _5947_/B _3558_/X _7286_/Q VGND VGND VPWR VPWR _3559_/X
+ sky130_fd_sc_hd__a32o_2
Xhold3100 _7157_/Q VGND VGND VPWR VPWR hold3100/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout593_A fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3111 _7167_/Q VGND VGND VPWR VPWR hold3111/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3122 _6957_/Q VGND VGND VPWR VPWR hold3122/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_9_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3133 _6927_/Q VGND VGND VPWR VPWR hold3133/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3144 _7351_/Q VGND VGND VPWR VPWR hold3144/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2410 hold618/X VGND VGND VPWR VPWR _5967_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6278_ _7374_/Q _6116_/B _6084_/X _6110_/X _7438_/Q VGND VGND VPWR VPWR _6278_/X
+ sky130_fd_sc_hd__a32o_1
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4562_/B sky130_fd_sc_hd__clkbuf_2
Xhold3155 _6988_/Q VGND VGND VPWR VPWR hold3155/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5277__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR _4089_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2421 hold941/X VGND VGND VPWR VPWR _4458_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3166 _6911_/Q VGND VGND VPWR VPWR hold3166/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6474__B1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR _4860_/A sky130_fd_sc_hd__buf_6
Xhold2432 hold951/X VGND VGND VPWR VPWR _4350_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3177 _3924_/X VGND VGND VPWR VPWR _7215_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5911__B _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6800_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
X_5229_ _5222_/A _5091_/C _5213_/B _4916_/B VGND VGND VPWR VPWR _5231_/B sky130_fd_sc_hd__a31o_1
Xhold2443 _7365_/Q VGND VGND VPWR VPWR hold732/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3188 _7216_/Q VGND VGND VPWR VPWR _3858_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2454 _5629_/X VGND VGND VPWR VPWR hold650/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3199 _7606_/Q VGND VGND VPWR VPWR _6237_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3827__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1720 _5996_/X VGND VGND VPWR VPWR hold278/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2465 hold2465/A VGND VGND VPWR VPWR _5625_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1731 hold316/X VGND VGND VPWR VPWR _5656_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2476 hold905/X VGND VGND VPWR VPWR _4379_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1742 _7059_/Q VGND VGND VPWR VPWR hold382/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2487 _7138_/Q VGND VGND VPWR VPWR hold635/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1753 hold74/X VGND VGND VPWR VPWR _5760_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2498 hold670/X VGND VGND VPWR VPWR _4493_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1764 _7306_/Q VGND VGND VPWR VPWR _4078_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4527__B _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6226__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1775 _5789_/X VGND VGND VPWR VPWR hold335/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1786 hold308/X VGND VGND VPWR VPWR _5977_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1797 _7490_/Q VGND VGND VPWR VPWR hold330/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6241__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6529__A1 _7578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5201__A1 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5201__B2 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3763__B2 _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6465__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5821__B hold12/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6480__A3 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6217__B1 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4172__B _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6090__D _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4600_ _4843_/A _5073_/A VGND VGND VPWR VPWR _5222_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5580_ _5580_/A1 _5580_/A2 _5579_/X _5577_/Y VGND VGND VPWR VPWR _7208_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3754__A1 _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4531_ _4531_/A0 _5647_/A0 _4532_/S VGND VGND VPWR VPWR _4531_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3754__B2 _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold305 hold305/A VGND VGND VPWR VPWR _7569_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7250_ _7255_/CLK _7250_/D fanout565/X VGND VGND VPWR VPWR _7250_/Q sky130_fd_sc_hd__dfrtp_2
Xhold316 hold316/A VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6299__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4462_ _4462_/A0 _5840_/A1 _4466_/S VGND VGND VPWR VPWR _4462_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_159_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4665__A_N _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold327 _4275_/X VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold338 hold338/A VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold349 hold349/A VGND VGND VPWR VPWR _7261_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6201_ _7451_/Q _6144_/A _6116_/A _6089_/X _7507_/Q VGND VGND VPWR VPWR _6201_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3516__B _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3413_ _7538_/Q VGND VGND VPWR VPWR _3413_/Y sky130_fd_sc_hd__inv_2
X_4393_ _5754_/A1 _4393_/A1 _4393_/S VGND VGND VPWR VPWR _4393_/X sky130_fd_sc_hd__mux2_1
X_7181_ _7190_/CLK _7181_/D _6871_/A VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2523_A _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _7320_/Q _6082_/X _6094_/X _7504_/Q _6131_/X VGND VGND VPWR VPWR _6132_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5731__B _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6456__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4628__A _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6063_ _6932_/Q _6061_/X _6775_/B1 _4117_/B VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__a211o_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 hold2477/X VGND VGND VPWR VPWR hold2478/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1016 hold2466/X VGND VGND VPWR VPWR _7251_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__A2 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3532__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 hold2897/X VGND VGND VPWR VPWR hold2898/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1038 hold2736/X VGND VGND VPWR VPWR _7279_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5014_ _5328_/A _5328_/B _5339_/C _5018_/B VGND VGND VPWR VPWR _5014_/Y sky130_fd_sc_hd__nand4_2
Xhold1049 hold2919/X VGND VGND VPWR VPWR hold2920/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6208__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2892_A _7197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7268_/CLK _6965_/D _6873_/A VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_95_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5431__A1 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5916_ _5916_/A0 _5979_/A0 _5919_/S VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6896_ _7075_/CLK _6896_/D _6846_/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3993__A1 _6988_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3993__B2 _7319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5847_ hold27/X hold17/X _5847_/S VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5778_ hold43/X _5778_/A1 hold49/X VGND VGND VPWR VPWR _5778_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3745__A1 _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7517_ _7565_/CLK hold62/X fanout605/X VGND VGND VPWR VPWR _7517_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3745__B2 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4729_ _4984_/B _4802_/A _4733_/B _4733_/A VGND VGND VPWR VPWR _4834_/B sky130_fd_sc_hd__and4b_2
XFILLER_0_133_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4302__S _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7448_ _7521_/CLK _7448_/D fanout600/X VGND VGND VPWR VPWR _7448_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_102_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6695__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold850 hold850/A VGND VGND VPWR VPWR hold850/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold861 _4484_/X VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7379_ _7487_/CLK _7379_/D fanout593/X VGND VGND VPWR VPWR _7379_/Q sky130_fd_sc_hd__dfrtp_4
Xhold872 hold872/A VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold883 hold883/A VGND VGND VPWR VPWR hold883/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold894 hold894/A VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3442__A _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2240 hold561/X VGND VGND VPWR VPWR _5733_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2251 _7404_/Q VGND VGND VPWR VPWR hold903/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2262 _7342_/Q VGND VGND VPWR VPWR hold598/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2273 _7390_/Q VGND VGND VPWR VPWR hold582/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input139_A wb_dat_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2284 hold580/X VGND VGND VPWR VPWR _5829_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2295 _5652_/X VGND VGND VPWR VPWR hold501/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1550 _5827_/X VGND VGND VPWR VPWR hold272/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1561 _5635_/X VGND VGND VPWR VPWR hold224/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1572 _5906_/X VGND VGND VPWR VPWR hold242/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1583 hold19/X VGND VGND VPWR VPWR _3470_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1594 hold298/X VGND VGND VPWR VPWR _4397_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_67_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3984__B2 _7187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3617__A _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5489__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6686__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6150__A2 _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6438__B1 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6453__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5661__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6205__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6750_ wire346/X _6749_/Y _6960_/Q _6431_/Y VGND VGND VPWR VPWR _6750_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3962_ _6962_/Q _5632_/B _5640_/C _5794_/A _7399_/Q VGND VGND VPWR VPWR _3962_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5701_ _5701_/A0 _5953_/A1 _5703_/S VGND VGND VPWR VPWR _5701_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3975__A1 _7407_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3975__B2 _7001_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6681_ _7118_/Q _6427_/X _6679_/X _6680_/X VGND VGND VPWR VPWR _6681_/X sky130_fd_sc_hd__a211o_1
X_3893_ _7536_/Q _3590_/C _5947_/B _3565_/X _7464_/Q VGND VGND VPWR VPWR _3893_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_162_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2473_A _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5632_ _5992_/C _5632_/B _5992_/D VGND VGND VPWR VPWR _5633_/S sky130_fd_sc_hd__and3_1
XANTENNA__3727__A1 _7315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5563_ _5563_/A1 _4722_/Y _4741_/Y _5084_/C _5379_/X VGND VGND VPWR VPWR _5564_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3527__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7302_ _7501_/CLK _7302_/D fanout579/X VGND VGND VPWR VPWR _7302_/Q sky130_fd_sc_hd__dfrtp_4
X_4514_ _4514_/A0 _5586_/A0 _4514_/S VGND VGND VPWR VPWR _4514_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7624__RESET_B fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold102 hold102/A VGND VGND VPWR VPWR hold102/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5494_ _4595_/Y _4601_/Y _4605_/Y _4834_/Y _4583_/B VGND VGND VPWR VPWR _5496_/C
+ sky130_fd_sc_hd__o32a_1
Xhold113 hold113/A VGND VGND VPWR VPWR _7469_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold124 hold124/A VGND VGND VPWR VPWR hold124/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold135 hold135/A VGND VGND VPWR VPWR hold135/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6677__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7233_ _7255_/CLK _7233_/D fanout565/X VGND VGND VPWR VPWR _7233_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_110_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4445_ _4445_/A0 _5979_/A0 _4448_/S VGND VGND VPWR VPWR _4445_/X sky130_fd_sc_hd__mux2_1
Xhold146 hold146/A VGND VGND VPWR VPWR _7563_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold157 hold157/A VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold168 hold168/A VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold179 hold179/A VGND VGND VPWR VPWR hold179/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7164_ _7189_/CLK _7164_/D fanout572/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout604 fanout605/X VGND VGND VPWR VPWR fanout604/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4376_ _4449_/B _5938_/C _4388_/B _4551_/D VGND VGND VPWR VPWR _4381_/S sky130_fd_sc_hd__and4_4
Xfanout615 input124/X VGND VGND VPWR VPWR _4888_/B sky130_fd_sc_hd__buf_12
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _7447_/Q _6144_/A _6120_/B _6379_/B1 _7519_/Q VGND VGND VPWR VPWR _6115_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4358__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7095_ _7096_/CLK _7095_/D fanout605/X VGND VGND VPWR VPWR _7095_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6046_ _7594_/Q _6051_/C _6929_/Q _6045_/Y VGND VGND VPWR VPWR _7594_/D sky130_fd_sc_hd__o31a_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6444__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4805__B _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6601__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _7278_/CLK _6948_/D fanout580/X VGND VGND VPWR VPWR _7653_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6879_ _7075_/CLK _6879_/D _6830_/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_0_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3718__B2 _7443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6380__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3437__A _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6668__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6132__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4143__A1 _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold680 hold680/A VGND VGND VPWR VPWR hold680/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6683__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold691 _4505_/X VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6467__B _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5891__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2070 _4189_/X VGND VGND VPWR VPWR hold167/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2081 _7658_/A VGND VGND VPWR VPWR hold714/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5798__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2092 _4211_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_188_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1380 hold1791/X VGND VGND VPWR VPWR hold1792/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1391 hold1/X VGND VGND VPWR VPWR _4197_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_87_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4715__B _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6199__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3957__B2 _7197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6371__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput207 _3441_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
Xoutput218 _7656_/X VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
XANTENNA__6659__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput229 _7666_/X VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
XANTENNA__6123__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ _4230_/A0 _4229_/X _4232_/S VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5882__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4161_ _6940_/Q _4161_/A1 _7260_/Q VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_1
X_4092_ _4563_/C _4563_/D _4562_/A _4562_/B VGND VGND VPWR VPWR _4095_/C sky130_fd_sc_hd__nor4_1
XANTENNA__4328__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4625__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6802_ _7111_/Q _6802_/A2 _6802_/B1 _7109_/Q VGND VGND VPWR VPWR _6802_/X sky130_fd_sc_hd__a22o_1
X_4994_ _5158_/A _5038_/B _5180_/A VGND VGND VPWR VPWR _5035_/B sky130_fd_sc_hd__and3_1
XANTENNA__3948__A1 _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6733_ _7180_/Q _6058_/X _6728_/X _6732_/X _6430_/X VGND VGND VPWR VPWR _6733_/Y
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_45_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3945_ _7335_/Q _3531_/X _3667_/X _7021_/Q _3944_/X VGND VGND VPWR VPWR _3961_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6664_ _7593_/Q _7117_/Q _6408_/C _6663_/X VGND VGND VPWR VPWR _6664_/X sky130_fd_sc_hd__a31o_1
X_3876_ _6989_/Q _4346_/C _5623_/B _3875_/X VGND VGND VPWR VPWR _3879_/C sky130_fd_sc_hd__a31o_4
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5615_ _5615_/A0 _5903_/A0 _5618_/S VGND VGND VPWR VPWR _5615_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6595_ _7396_/Q _6420_/C _6588_/X _6590_/X _6594_/X VGND VGND VPWR VPWR _6595_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_143_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5546_ _4741_/Y _4886_/Y _4891_/Y _4894_/Y VGND VGND VPWR VPWR _5546_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_143_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5477_ _5107_/A _5282_/B wire529/X _5105_/X _5395_/X VGND VGND VPWR VPWR _5559_/B
+ sky130_fd_sc_hd__a311o_1
XANTENNA__4125__A1 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7216_ _7075_/CLK _7216_/D _6868_/X VGND VGND VPWR VPWR _7216_/Q sky130_fd_sc_hd__dfrtn_1
X_4428_ _7107_/Q _4428_/B VGND VGND VPWR VPWR _4428_/Y sky130_fd_sc_hd__nand2b_4
XANTENNA__3479__A3 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout412 _3489_/Y VGND VGND VPWR VPWR _4491_/A sky130_fd_sc_hd__buf_12
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _4169_/B2
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5873__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout423 _6073_/X VGND VGND VPWR VPWR _6317_/C sky130_fd_sc_hd__buf_12
Xfanout434 _6404_/Y VGND VGND VPWR VPWR _6459_/B sky130_fd_sc_hd__buf_12
X_7147_ _7447_/CLK _7147_/D fanout598/X VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout445 _6023_/Y VGND VGND VPWR VPWR _6097_/B sky130_fd_sc_hd__buf_6
X_4359_ _4359_/A0 _5840_/A1 _4363_/S VGND VGND VPWR VPWR _4359_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout467 hold1476/X VGND VGND VPWR VPWR hold1477/A sky130_fd_sc_hd__buf_6
Xfanout478 hold2072/X VGND VGND VPWR VPWR _5979_/A0 sky130_fd_sc_hd__buf_12
X_7078_ _7096_/CLK _7078_/D fanout605/X VGND VGND VPWR VPWR _7658_/A sky130_fd_sc_hd__dfrtp_1
Xfanout489 hold43/X VGND VGND VPWR VPWR _5805_/A1 sky130_fd_sc_hd__buf_12
XANTENNA__5625__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6029_ _6027_/X _6028_/Y _6051_/C VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3636__B1 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4871__B_N _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6586__C1 _6585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A1 _7137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4551__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6353__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input67_A mgmt_gpio_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6105__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5616__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3890__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6041__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _7571_/Q _5983_/A _4491_/B _4422_/S input48/X VGND VGND VPWR VPWR _3730_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4461__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3661_ _4473_/A _4551_/C _4491_/C VGND VGND VPWR VPWR _3661_/X sky130_fd_sc_hd__and3_2
XANTENNA__4180__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6344__A2 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5001__C1 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4355__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5400_ _5397_/X _5482_/A _5481_/B VGND VGND VPWR VPWR _5400_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_0_153_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6380_ _7005_/Q _6097_/B _6120_/B _6379_/X VGND VGND VPWR VPWR _6380_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3508__C _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3592_ _7437_/Q _3525_/X _3590_/X _3591_/X _3589_/X VGND VGND VPWR VPWR _3592_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_141_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ _4605_/Y _4759_/Y _5007_/Y _4690_/Y _5184_/X VGND VGND VPWR VPWR _5331_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA_hold2436_A _7154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5262_ _5451_/A1 _4737_/Y _5255_/X _5077_/Y _4709_/Y VGND VGND VPWR VPWR _5564_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7001_ _7144_/CLK _7001_/D fanout572/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_4
X_4213_ _4213_/A0 _5948_/A1 _4214_/S VGND VGND VPWR VPWR _4213_/X sky130_fd_sc_hd__mux2_1
Xhold2806 hold2806/A VGND VGND VPWR VPWR hold2806/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2817 hold2817/A VGND VGND VPWR VPWR hold2817/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_167_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5193_ _5183_/A _5053_/C _5188_/X _5192_/X _5171_/X VGND VGND VPWR VPWR _5193_/X
+ sky130_fd_sc_hd__a311o_1
Xhold2828 hold2828/A VGND VGND VPWR VPWR hold2828/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2839 _7632_/Q VGND VGND VPWR VPWR _6786_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3866__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2603_A _7480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4144_ _4144_/A _4174_/B VGND VGND VPWR VPWR _4144_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_183_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6835__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5607__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3881__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4075_ hold41/A _4076_/B _4075_/S VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3618__B1 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_4_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__3633__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4977_ _5138_/A _5138_/B _5138_/D VGND VGND VPWR VPWR _4977_/X sky130_fd_sc_hd__and3_2
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6583__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6716_ _7053_/Q _6434_/B _6771_/A3 _6466_/X _7211_/Q VGND VGND VPWR VPWR _6716_/X
+ sky130_fd_sc_hd__a32o_1
X_3928_ _6897_/Q _6882_/Q _7248_/Q VGND VGND VPWR VPWR _3929_/A sky130_fd_sc_hd__nor3_2
XFILLER_0_117_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout519_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6647_ _6647_/A _6647_/B _6647_/C _6647_/D VGND VGND VPWR VPWR _6647_/Y sky130_fd_sc_hd__nor4_1
XANTENNA__6335__A2 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3859_ _3859_/A hold36/A _4551_/C _5992_/C VGND VGND VPWR VPWR _3859_/X sky130_fd_sc_hd__and4_2
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6578_ _7388_/Q _6413_/C _6426_/X _6577_/X VGND VGND VPWR VPWR _6578_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4897__A2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5529_ _5529_/A _5529_/B _5529_/C _5529_/D VGND VGND VPWR VPWR _5533_/A sky130_fd_sc_hd__and4_1
XANTENNA__6638__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5846__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7179__SET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4129__A_N _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input121_A wb_adr_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4265__B _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3624__A3 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_csclk_A _4169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5377__A3 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5782__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4281__A _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5096__B _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6326__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5129__A3 _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4337__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3560__A2 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3848__B1 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6262__B2 _7366_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4175__B input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4900_ _4601_/Y _4622_/Y _4726_/Y _4895_/Y _4896_/Y VGND VGND VPWR VPWR _4902_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_87_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5880_ _5880_/A0 _5997_/A1 _5883_/S VGND VGND VPWR VPWR _5880_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4831_ _4831_/A _4860_/A _4909_/D _4786_/C VGND VGND VPWR VPWR _5072_/C sky130_fd_sc_hd__nor4b_4
XFILLER_0_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6565__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6892__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7550_ _7555_/CLK _7550_/D fanout594/X VGND VGND VPWR VPWR _7550_/Q sky130_fd_sc_hd__dfrtp_2
X_4762_ _4772_/A _4801_/B _4803_/A _5404_/B VGND VGND VPWR VPWR _4763_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_6_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6501_ _7529_/Q _6058_/X _6422_/X _7289_/Q _6500_/X VGND VGND VPWR VPWR _6501_/X
+ sky130_fd_sc_hd__a221o_1
X_3713_ _7291_/Q _4212_/A _5731_/B input30/X _3503_/X VGND VGND VPWR VPWR _3713_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__3519__B _3519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7481_ _7560_/CLK _7481_/D fanout599/X VGND VGND VPWR VPWR _7481_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__7050__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4693_ _4733_/A _4733_/B _4801_/C VGND VGND VPWR VPWR _4794_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_172_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2553_A _7309_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6432_ _7527_/Q _6058_/X _6424_/X _7567_/Q VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__a22o_1
X_3644_ _7218_/Q _3643_/Y _3923_/S VGND VGND VPWR VPWR _3644_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_153_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6363_ _7054_/Q _6121_/A _6120_/B _6317_/C _7049_/Q VGND VGND VPWR VPWR _6363_/X
+ sky130_fd_sc_hd__a32o_1
X_3575_ input27/X _3488_/X _3490_/X input18/X _3574_/X VGND VGND VPWR VPWR _3575_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA_hold2720_A _7201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3535__A hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5314_ _5314_/A _5535_/A VGND VGND VPWR VPWR _5317_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5453__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3551__A2 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6294_ _7016_/Q _6086_/X _6121_/C _6988_/Q _6121_/X VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2603 _7480_/Q VGND VGND VPWR VPWR hold2603/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5245_ _4571_/Y _4843_/A _4879_/C _4960_/A VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__o22a_1
Xhold2614 hold872/X VGND VGND VPWR VPWR _5810_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__buf_8
Xhold2625 _7325_/Q VGND VGND VPWR VPWR hold841/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2636 hold862/X VGND VGND VPWR VPWR _5774_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2647 hold651/X VGND VGND VPWR VPWR _5997_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1902 hold292/X VGND VGND VPWR VPWR _5744_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2658 _7448_/Q VGND VGND VPWR VPWR hold2658/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1913 _5599_/X VGND VGND VPWR VPWR hold521/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5176_ _4605_/Y _4690_/Y _4971_/X _5014_/Y _5175_/X VGND VGND VPWR VPWR _5176_/X
+ sky130_fd_sc_hd__o311a_1
Xhold1924 hold524/X VGND VGND VPWR VPWR _4194_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2669 _7030_/Q VGND VGND VPWR VPWR hold765/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1935 _7247_/Q VGND VGND VPWR VPWR hold390/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4127_ input83/X _4127_/A1 _6896_/Q VGND VGND VPWR VPWR _4127_/X sky130_fd_sc_hd__mux2_1
Xhold1946 _6877_/Q VGND VGND VPWR VPWR hold466/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1957 _7165_/Q VGND VGND VPWR VPWR hold424/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1968 _7039_/Q VGND VGND VPWR VPWR hold422/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout469_A hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6253__B2 hold76/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1979 _7135_/Q VGND VGND VPWR VPWR hold452/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_127_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4058_ _7071_/Q _7074_/Q _7073_/Q VGND VGND VPWR VPWR _4058_/Y sky130_fd_sc_hd__nor3b_4
XANTENNA__5896__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_164_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6556__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5764__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6308__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3790__A2 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1820_A _7569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3445__A _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6459__C _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input169_A wb_stb_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3845__A3 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output290_A _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire462 _4430_/C VGND VGND VPWR VPWR wire462/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3781__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold509 hold509/A VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6180__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3533__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6483__A1 _7352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5286__A2 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5030_ _5038_/A _5038_/B _5030_/C VGND VGND VPWR VPWR _5031_/B sky130_fd_sc_hd__and3_1
XANTENNA__6483__B2 _7360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1209 hold2925/X VGND VGND VPWR VPWR hold1209/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_164_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2301_A _7510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3521__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6981_ _7633_/CLK _6981_/D VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfxtp_1
X_5932_ _5986_/A1 _5932_/A1 _5937_/S VGND VGND VPWR VPWR _5932_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5863_ _5863_/A0 _5863_/A1 _5865_/S VGND VGND VPWR VPWR _5863_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6538__A2 _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7602_ _7623_/CLK _7602_/D fanout575/X VGND VGND VPWR VPWR _7602_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4125__S _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4814_ _4909_/D _5260_/B _4814_/C VGND VGND VPWR VPWR _4814_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_173_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5794_ _5794_/A hold47/X VGND VGND VPWR VPWR _5802_/S sky130_fd_sc_hd__nand2_8
XANTENNA__4352__C _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7533_ _7578_/CLK _7533_/D fanout596/X VGND VGND VPWR VPWR _7533_/Q sky130_fd_sc_hd__dfrtp_4
X_4745_ _5100_/A _5079_/B _4755_/C VGND VGND VPWR VPWR _4746_/C sky130_fd_sc_hd__and3_1
XFILLER_0_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7464_ _7530_/CLK _7464_/D fanout600/X VGND VGND VPWR VPWR _7464_/Q sky130_fd_sc_hd__dfstp_4
X_4676_ _4675_/A _4675_/B _4675_/C _5071_/A VGND VGND VPWR VPWR _4679_/A sky130_fd_sc_hd__a31o_2
XFILLER_0_71_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6415_ _6427_/A _6467_/A _6747_/C VGND VGND VPWR VPWR _6419_/A sky130_fd_sc_hd__and3_4
XFILLER_0_114_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3627_ _7340_/Q _3531_/X _3532_/X input57/X _3626_/X VGND VGND VPWR VPWR _3632_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6171__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7395_ _7395_/CLK _7395_/D fanout598/X VGND VGND VPWR VPWR _7395_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6710__A2 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6346_ _7008_/Q _6082_/X _6097_/X _7184_/Q _6345_/X VGND VGND VPWR VPWR _6346_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5183__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3558_ _5590_/A _5640_/B _5640_/C VGND VGND VPWR VPWR _3558_/X sky130_fd_sc_hd__and3_4
Xhold3101 hold3101/A VGND VGND VPWR VPWR _4504_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3112 hold3112/A VGND VGND VPWR VPWR _4516_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3123 hold3123/A VGND VGND VPWR VPWR _4260_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3134 hold3134/A VGND VGND VPWR VPWR _4213_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6277_ _7422_/Q _6072_/X _6097_/X hold27/A _6276_/X VGND VGND VPWR VPWR _6280_/C
+ sky130_fd_sc_hd__a221o_1
Xhold2400 _4448_/X VGND VGND VPWR VPWR hold634/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout586_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3489_ _3507_/A _3576_/C VGND VGND VPWR VPWR _3489_/Y sky130_fd_sc_hd__nor2_2
Xhold3145 hold3145/A VGND VGND VPWR VPWR _5741_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__clkbuf_2
Xhold3156 hold3156/A VGND VGND VPWR VPWR _4304_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2411 _5967_/X VGND VGND VPWR VPWR hold619/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2422 _7348_/Q VGND VGND VPWR VPWR hold2422/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3167 hold3167/A VGND VGND VPWR VPWR _4192_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6474__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5228_ _5228_/A _5228_/B _5228_/C _5228_/D VGND VGND VPWR VPWR _5231_/A sky130_fd_sc_hd__nand4_1
XANTENNA__6474__B2 _7528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4564_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2433 _7232_/Q VGND VGND VPWR VPWR hold939/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3178 _7214_/Q VGND VGND VPWR VPWR _3997_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3189 _7108_/Q VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2444 hold732/X VGND VGND VPWR VPWR _5756_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2455 _7372_/Q VGND VGND VPWR VPWR hold977/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1710 _4512_/X VGND VGND VPWR VPWR hold333/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1721 _6883_/Q VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2466 _5625_/X VGND VGND VPWR VPWR hold2466/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3827__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2477 _7238_/Q VGND VGND VPWR VPWR hold2477/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1732 _5656_/X VGND VGND VPWR VPWR hold317/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1743 hold382/X VGND VGND VPWR VPWR _4392_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5159_ _5410_/A _4810_/C _5453_/B _5158_/X VGND VGND VPWR VPWR _5160_/D sky130_fd_sc_hd__a31o_1
Xhold2488 hold635/X VGND VGND VPWR VPWR _4481_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2499 _6960_/Q VGND VGND VPWR VPWR hold971/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4527__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1754 _5760_/X VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1765 hold284/X VGND VGND VPWR VPWR _5690_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1776 hold335/X VGND VGND VPWR VPWR _7394_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1787 _5977_/X VGND VGND VPWR VPWR hold309/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1798 hold330/X VGND VGND VPWR VPWR _5897_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6631__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6529__A2 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5201__A2 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3763__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6162__B1 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3249_A _7221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6465__A1 _7303_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5821__C hold48/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6768__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output303_A _3578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5976__A0 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4530_ _4530_/A0 _5815_/A1 _4532_/S VGND VGND VPWR VPWR _4530_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3754__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold306 hold306/A VGND VGND VPWR VPWR hold306/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6153__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4461_ _4473_/A _4551_/A _4551_/C _4551_/D VGND VGND VPWR VPWR _4466_/S sky130_fd_sc_hd__and4_4
Xhold317 hold317/A VGND VGND VPWR VPWR _7276_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold328 hold328/A VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_159_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6099__C _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold339 hold339/A VGND VGND VPWR VPWR _7460_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6200_ _7467_/Q _6121_/A _6120_/B _6317_/C _7515_/Q VGND VGND VPWR VPWR _6200_/X
+ sky130_fd_sc_hd__a32o_1
X_3412_ _7546_/Q VGND VGND VPWR VPWR _3412_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7180_ _7190_/CLK _7180_/D _6871_/A VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4392_ _5951_/A1 _4392_/A1 _4393_/S VGND VGND VPWR VPWR _4392_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6131_ _7408_/Q _6121_/C _6116_/C _6136_/C VGND VGND VPWR VPWR _6131_/X sky130_fd_sc_hd__o211a_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A2 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6456__A1 _7487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5731__C hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6062_ _6009_/Y _6019_/Y _6061_/X _6932_/Q VGND VGND VPWR VPWR _6062_/X sky130_fd_sc_hd__a22o_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4628__B _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _5607_/X VGND VGND VPWR VPWR _7238_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1017 hold2717/X VGND VGND VPWR VPWR hold2718/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3532__B _3537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5013_ _5158_/A _5183_/A _5013_/C VGND VGND VPWR VPWR _5013_/X sky130_fd_sc_hd__and3_2
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 hold2899/X VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1039 hold2889/X VGND VGND VPWR VPWR hold2890/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_23_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3690__A1 _7331_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6759__A2 _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6964_ _7189_/CLK _6964_/D fanout572/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5915_ _5915_/A0 _5996_/A1 _5919_/S VGND VGND VPWR VPWR _5915_/X sky130_fd_sc_hd__mux2_1
X_6895_ _7075_/CLK _6895_/D _6845_/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5719__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_192_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5846_ _5846_/A0 hold61/X _5847_/S VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3993__A2 _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6392__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5777_ _5993_/A1 _5777_/A1 hold49/X VGND VGND VPWR VPWR _5777_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_173_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4728_ _5260_/C _5387_/D _4790_/B VGND VGND VPWR VPWR _4763_/A sky130_fd_sc_hd__and3_1
XANTENNA_fanout501_A _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3745__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7516_ _7565_/CLK _7516_/D fanout603/X VGND VGND VPWR VPWR _7516_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_161_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7447_ _7447_/CLK _7447_/D fanout598/X VGND VGND VPWR VPWR _7447_/Q sky130_fd_sc_hd__dfstp_4
X_4659_ _5248_/A _5248_/B VGND VGND VPWR VPWR _4659_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_101_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6695__A1 _7138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold840 hold840/A VGND VGND VPWR VPWR _7285_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7378_ _7575_/CLK _7378_/D fanout595/X VGND VGND VPWR VPWR _7378_/Q sky130_fd_sc_hd__dfrtp_4
Xhold851 hold851/A VGND VGND VPWR VPWR _7429_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold862 hold862/A VGND VGND VPWR VPWR hold862/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold873 _5810_/X VGND VGND VPWR VPWR _7413_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6329_ _6958_/Q _6036_/Y _6775_/B1 VGND VGND VPWR VPWR _6329_/X sky130_fd_sc_hd__o21a_1
Xhold884 _5765_/X VGND VGND VPWR VPWR _7373_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold895 hold895/A VGND VGND VPWR VPWR hold895/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold281_A _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2230 _5712_/X VGND VGND VPWR VPWR hold571/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2241 _7502_/Q VGND VGND VPWR VPWR hold526/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2252 hold903/X VGND VGND VPWR VPWR _5800_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2263 hold598/X VGND VGND VPWR VPWR _5730_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2274 hold582/X VGND VGND VPWR VPWR _5784_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2285 _5829_/X VGND VGND VPWR VPWR hold581/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1540 hold200/X VGND VGND VPWR VPWR _7545_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2296 _7412_/Q VGND VGND VPWR VPWR hold909/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1551 hold272/X VGND VGND VPWR VPWR _7428_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1562 hold224/X VGND VGND VPWR VPWR _7258_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1573 _7353_/Q VGND VGND VPWR VPWR hold267/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1584 _3470_/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1595 _4397_/X VGND VGND VPWR VPWR hold299/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_67_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3984__A2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input97_A usr2_vcc_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_33_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3617__B _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6135__B1 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6150__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_csclk _7267_/CLK VGND VGND VPWR VPWR _7510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6438__A1 _7391_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7582_/CLK sky130_fd_sc_hd__clkbuf_16
X_3961_ _3961_/A _3961_/B _3961_/C _3961_/D VGND VGND VPWR VPWR _3995_/B sky130_fd_sc_hd__nor4_1
XANTENNA__5994__S hold37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5700_ _5700_/A0 hold84/X _5703_/S VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__mux2_1
X_6680_ _7052_/Q _6434_/B _6771_/A3 _6463_/X _7163_/Q VGND VGND VPWR VPWR _6680_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3892_ _7360_/Q _5803_/A hold12/A _3891_/X VGND VGND VPWR VPWR _3892_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_161_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5631_ _5640_/D _5631_/B VGND VGND VPWR VPWR _7256_/D sky130_fd_sc_hd__and2_1
XANTENNA__5177__A1 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4911__B _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5295__A _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3727__A2 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5562_ _5393_/X _5478_/B _5562_/C _5562_/D VGND VGND VPWR VPWR _5562_/Y sky130_fd_sc_hd__nand4bb_1
XFILLER_0_115_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7301_ _7412_/CLK _7301_/D fanout580/X VGND VGND VPWR VPWR _7301_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3527__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4513_ _4513_/A0 _5852_/A0 _4514_/S VGND VGND VPWR VPWR _4513_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6126__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold103 _5907_/X VGND VGND VPWR VPWR _7499_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5493_ _4595_/Y _4832_/Y _5528_/A3 _5492_/X VGND VGND VPWR VPWR _5493_/Y sky130_fd_sc_hd__o31ai_1
Xhold114 hold114/A VGND VGND VPWR VPWR hold114/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7232_ _7255_/CLK _7232_/D fanout565/X VGND VGND VPWR VPWR _7232_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6677__A1 _7178_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold125 hold125/A VGND VGND VPWR VPWR _6955_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold136 hold136/A VGND VGND VPWR VPWR _7099_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4444_ _4444_/A0 _5996_/A1 _4448_/S VGND VGND VPWR VPWR _4444_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold147 hold147/A VGND VGND VPWR VPWR hold147/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6838__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold158 hold158/A VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6141__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold169 hold169/A VGND VGND VPWR VPWR hold169/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7163_ _7213_/CLK _7163_/D fanout590/X VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_4
X_4375_ _5979_/A0 _4375_/A1 _4375_/S VGND VGND VPWR VPWR _4375_/X sky130_fd_sc_hd__mux2_1
Xfanout605 fanout606/X VGND VGND VPWR VPWR fanout605/X sky130_fd_sc_hd__buf_12
Xfanout616 input124/X VGND VGND VPWR VPWR _4887_/B sky130_fd_sc_hd__buf_12
XANTENNA__3543__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6114_ _7383_/Q _6109_/X _6110_/X _7431_/Q _6113_/X VGND VGND VPWR VPWR _6114_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7096_/CLK _7094_/D fanout605/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4358__B _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6434_/B _6574_/B _6051_/C VGND VGND VPWR VPWR _6045_/Y sky130_fd_sc_hd__o21ai_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5101__A1 _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6854__A _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6601__A1 _7517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4093__B _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6947_ _7278_/CLK _6947_/D fanout580/X VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4612__B1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3966__A2 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6878_ _7201_/CLK _6878_/D _6833_/A VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5829_ _5829_/A0 _5991_/A1 _5829_/S VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4821__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1566_A _7452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3718__A2 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6380__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6117__B1 _6116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1733_A _7533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4143__A2 _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold670 hold670/A VGND VGND VPWR VPWR hold670/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold681 hold681/A VGND VGND VPWR VPWR _7547_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6467__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold692 hold692/A VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input151_A wb_dat_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2060 hold622/X VGND VGND VPWR VPWR _5849_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2071 hold167/X VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2082 hold714/X VGND VGND VPWR VPWR _4413_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2093 _7659_/A VGND VGND VPWR VPWR hold775/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1370 _7577_/Q VGND VGND VPWR VPWR _5995_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1381 hold2281/X VGND VGND VPWR VPWR hold2282/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input12_A mask_rev_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1392 _4197_/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_59_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4715__C _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6356__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4223__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6371__A3 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6108__B1 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput208 _3440_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XFILLER_0_11_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6659__B2 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput219 _7657_/X VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5331__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5331__B2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ _7282_/Q input1/X _4159_/Y VGND VGND VPWR VPWR _4160_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__6081__B_N _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4178__B _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3893__B2 _7464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4091_ _4562_/C _4562_/D _4091_/C input116/X VGND VGND VPWR VPWR _4093_/D sky130_fd_sc_hd__nor4b_1
XFILLER_0_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4625__C _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6801_ _6800_/X hold462/A _6822_/S VGND VGND VPWR VPWR _7637_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_175_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5398__A1 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4993_ _5295_/C _5038_/B _5180_/A VGND VGND VPWR VPWR _5035_/A sky130_fd_sc_hd__and3_1
XFILLER_0_93_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3944_ _6897_/Q _6882_/Q _7248_/Q _5587_/C _5619_/B VGND VGND VPWR VPWR _3944_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA__3948__A2 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6732_ _7130_/Q _6424_/X _6730_/X _6731_/X VGND VGND VPWR VPWR _6732_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_129_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6663_ _7172_/Q _6747_/B _6747_/C _6408_/A _7147_/Q VGND VGND VPWR VPWR _6663_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3875_ _6928_/Q _4212_/A _5659_/B _3861_/X VGND VGND VPWR VPWR _3875_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_73_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3538__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4133__S _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5614_ _5947_/A _5614_/B hold47/X VGND VGND VPWR VPWR _5614_/X sky130_fd_sc_hd__and3_2
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6594_ _7516_/Q _6435_/X _6591_/X _6593_/X VGND VGND VPWR VPWR _6594_/X sky130_fd_sc_hd__a211o_4
XFILLER_0_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_777 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5545_ _5545_/A _5545_/B _5545_/C _5545_/D VGND VGND VPWR VPWR _5548_/B sky130_fd_sc_hd__nor4_1
XFILLER_0_170_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3581__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_5476_ _5476_/A _5476_/B _5476_/C VGND VGND VPWR VPWR _5478_/B sky130_fd_sc_hd__nand3_1
X_4427_ _4427_/A _7109_/Q _7110_/Q _7111_/Q VGND VGND VPWR VPWR _4430_/C sky130_fd_sc_hd__nor4_4
X_7215_ _4150_/A1 _7215_/D _6867_/X VGND VGND VPWR VPWR _7215_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_0_111_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout499_A hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout413 hold71/X VGND VGND VPWR VPWR _4449_/B sky130_fd_sc_hd__buf_12
X_7146_ _7266_/CLK _7146_/D fanout567/X VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_4
X_4358_ _4473_/A _4551_/C _4491_/C _4551_/D VGND VGND VPWR VPWR _4363_/S sky130_fd_sc_hd__and4_4
Xfanout435 _6645_/C VGND VGND VPWR VPWR _6747_/C sky130_fd_sc_hd__buf_12
XANTENNA__3884__A1 _7528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout446 _6022_/X VGND VGND VPWR VPWR _6136_/B sky130_fd_sc_hd__buf_12
XANTENNA__5899__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout457 _5451_/A1 VGND VGND VPWR VPWR _5563_/A1 sky130_fd_sc_hd__buf_8
XANTENNA_input4_A mask_rev_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout468 hold61/X VGND VGND VPWR VPWR _5954_/A1 sky130_fd_sc_hd__clkbuf_16
X_7077_ _7096_/CLK _7077_/D fanout605/X VGND VGND VPWR VPWR _7657_/A sky130_fd_sc_hd__dfrtp_1
Xfanout479 _5951_/A1 VGND VGND VPWR VPWR _5647_/A0 sky130_fd_sc_hd__buf_12
X_4289_ _3570_/Y _4289_/A1 _4289_/S VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__mux2_1
X_6028_ _7589_/Q _7588_/Q _6106_/B VGND VGND VPWR VPWR _6028_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__3636__A1 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3636__B2 _7532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5389__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A2 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4551__B _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6105__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3627__B2 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6577__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6329__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4461__B _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3660_ _5830_/C _4491_/A _4491_/B VGND VGND VPWR VPWR _4467_/A sky130_fd_sc_hd__and3_4
XANTENNA__4180__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6344__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5552__A1 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3591_ input59/X _3933_/A _3519_/B _5704_/A _7325_/Q VGND VGND VPWR VPWR _3591_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_141_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5330_ _4605_/Y _4759_/Y _5007_/Y _4690_/Y _5173_/X VGND VGND VPWR VPWR _5554_/A
+ sky130_fd_sc_hd__o221a_1
X_5261_ _4709_/Y _4727_/Y _4946_/Y _5077_/Y _5260_/Y VGND VGND VPWR VPWR _5265_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5304__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6501__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2331_A _7323_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7000_ _7633_/CLK _7000_/D VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfxtp_1
X_4212_ _4212_/A _5640_/C _5640_/D VGND VGND VPWR VPWR _4214_/S sky130_fd_sc_hd__and3_1
Xhold2807 hold2807/A VGND VGND VPWR VPWR hold2807/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5192_ _5034_/C _5188_/X _5190_/X _5191_/X VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__a211o_1
Xhold2818 _6993_/Q VGND VGND VPWR VPWR _4310_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2829 _7439_/Q VGND VGND VPWR VPWR hold2829/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4143_ _7570_/Q _4142_/A _4142_/Y VGND VGND VPWR VPWR _4143_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA_clkbuf_leaf_2_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4074_ hold7/A hold41/A _4075_/S VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3618__B2 _7316_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5083__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2798_A _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6568__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4976_ _4956_/A _4956_/B _4975_/X _4826_/Y VGND VGND VPWR VPWR _5438_/B sky130_fd_sc_hd__a211o_1
XANTENNA__5240__B1 wire533/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6583__A3 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6715_ _6969_/Q _6420_/A _6704_/X _6714_/X VGND VGND VPWR VPWR _6715_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_135_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3927_ _7263_/Q _5722_/A _5640_/B _5640_/C VGND VGND VPWR VPWR _3927_/X sky130_fd_sc_hd__and4_2
XANTENNA__5791__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3858_ _3858_/A1 _3996_/A _3856_/Y _3857_/X VGND VGND VPWR VPWR _7216_/D sky130_fd_sc_hd__a22o_1
X_6646_ _7462_/Q _6455_/X _6645_/X _6644_/X _6643_/X VGND VGND VPWR VPWR _6647_/D
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6335__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6577_ _7484_/Q _6447_/C _6459_/C _6421_/X _7324_/Q VGND VGND VPWR VPWR _6577_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6740__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3789_ _7346_/Q _3590_/C _3669_/C _3525_/X _7434_/Q VGND VGND VPWR VPWR _3789_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_116_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3554__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4897__A3 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5528_ _4595_/Y _4832_/Y _5528_/A3 _5422_/D _5294_/A VGND VGND VPWR VPWR _5529_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5459_ _5222_/A _5107_/A _5248_/A _5458_/X VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_2_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1529_A _7532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7129_ _7415_/CLK _7129_/D fanout593/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4827__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_wb_clk_i clkbuf_3_7_0_wb_clk_i/X VGND VGND VPWR VPWR _7644_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6271__A2 _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4265__C _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4282__A1 _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input114_A wb_adr_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold3279_A _6879_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6731__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3848__A1 _7226_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4737__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6262__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4273__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4830_ _4830_/A _4830_/B _4830_/C VGND VGND VPWR VPWR _4837_/A sky130_fd_sc_hd__nor3_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4903__C _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _4772_/A _4801_/B _5404_/B VGND VGND VPWR VPWR _4761_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__4191__B _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5773__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2281_A _7291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6500_ _7369_/Q _6651_/B _6651_/C _6457_/X _7473_/Q VGND VGND VPWR VPWR _6500_/X
+ sky130_fd_sc_hd__a32o_1
X_3712_ _7515_/Q _5920_/A _3704_/X _3706_/X _3711_/X VGND VGND VPWR VPWR _3732_/B
+ sky130_fd_sc_hd__a2111o_2
X_7480_ _7565_/CLK _7480_/D fanout600/X VGND VGND VPWR VPWR _7480_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3519__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4692_ _5038_/A _4758_/B _5328_/B VGND VGND VPWR VPWR _4692_/Y sky130_fd_sc_hd__nand3_4
XANTENNA_clkbuf_3_6_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6431_ _6431_/A _6431_/B _6431_/C VGND VGND VPWR VPWR _6431_/Y sky130_fd_sc_hd__nand3_4
X_3643_ _3643_/A _3643_/B _3643_/C VGND VGND VPWR VPWR _3643_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__6722__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4411__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6362_ _6357_/X _6362_/B _6362_/C VGND VGND VPWR VPWR _6362_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_113_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7090__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3574_ _7573_/Q _5911_/A _5965_/A hold72/A _7565_/Q VGND VGND VPWR VPWR _3574_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3535__B _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5313_ _4723_/Y _4796_/Y _4978_/Y _4793_/Y _5312_/X VGND VGND VPWR VPWR _5535_/A
+ sky130_fd_sc_hd__o221a_1
X_6293_ _7021_/Q _6070_/X _6087_/X _7051_/Q _6292_/X VGND VGND VPWR VPWR _6293_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3551__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5244_ _5367_/B _5545_/A _5244_/C VGND VGND VPWR VPWR _5247_/B sky130_fd_sc_hd__nor3_1
Xhold2604 hold2604/A VGND VGND VPWR VPWR _5886_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3839__A1 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2615 _7357_/Q VGND VGND VPWR VPWR hold854/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3839__B2 _7199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2626 hold841/X VGND VGND VPWR VPWR _5711_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5175_ _4956_/B _5174_/Y _5012_/Y VGND VGND VPWR VPWR _5175_/X sky130_fd_sc_hd__a21o_1
Xhold2637 _7571_/Q VGND VGND VPWR VPWR hold639/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2648 _7555_/Q VGND VGND VPWR VPWR hold688/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1903 _5744_/X VGND VGND VPWR VPWR hold293/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2659 hold2659/A VGND VGND VPWR VPWR _5850_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1914 _7573_/Q VGND VGND VPWR VPWR hold114/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1925 _4194_/X VGND VGND VPWR VPWR hold525/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4126_ _6897_/Q _4128_/B VGND VGND VPWR VPWR _4126_/Y sky130_fd_sc_hd__nor2_1
Xhold1936 hold390/X VGND VGND VPWR VPWR _5618_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1947 hold466/X VGND VGND VPWR VPWR _4188_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1958 hold424/X VGND VGND VPWR VPWR _4513_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1969 hold422/X VGND VGND VPWR VPWR _4368_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4057_ _4057_/A0 _4076_/B _4057_/S VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4264__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout531_A _4940_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4382__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6556__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4813__C _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_163_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4959_ _5248_/A _5248_/B _5453_/C _4953_/X _5113_/A VGND VGND VPWR VPWR _4959_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_164_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3775__B1 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7178__RESET_B fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6308__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6629_ _7542_/Q _6408_/D _6435_/X _7518_/Q VGND VGND VPWR VPWR _6629_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3790__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5516__B2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4321__S _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6492__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4255__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5755__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3766__B1 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3781__A3 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire452 _4825_/Y VGND VGND VPWR VPWR _5113_/B sky130_fd_sc_hd__buf_2
Xwire463 wire463/A VGND VGND VPWR VPWR _4428_/B sky130_fd_sc_hd__buf_4
XANTENNA__4231__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6180__A1 _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6180__B2 _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3533__A3 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6483__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5286__A3 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4494__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5691__A0 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5997__S hold37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6235__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4246__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6980_ _7633_/CLK _6980_/D VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5931_ _5985_/A1 _5931_/A1 _5937_/S VGND VGND VPWR VPWR _5931_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4914__B _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5994__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5862_ _5997_/A1 _5862_/A1 _5865_/S VGND VGND VPWR VPWR _5862_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6538__A3 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7601_ _7601_/CLK _7601_/D fanout569/X VGND VGND VPWR VPWR _7601_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5746__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4813_ _4984_/B _5260_/B _4814_/C VGND VGND VPWR VPWR _5399_/C sky130_fd_sc_hd__and3_4
XFILLER_0_145_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5793_ _5793_/A0 _5991_/A1 _5793_/S VGND VGND VPWR VPWR _5793_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5210__A3 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3757__B1 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7532_ _7566_/CLK _7532_/D fanout596/X VGND VGND VPWR VPWR _7532_/Q sky130_fd_sc_hd__dfrtp_4
X_4744_ _4879_/C _5282_/B VGND VGND VPWR VPWR _4744_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_44_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4675_ _4675_/A _4675_/B _4675_/C VGND VGND VPWR VPWR _4675_/Y sky130_fd_sc_hd__nand3_2
X_7463_ _7565_/CLK _7463_/D fanout599/X VGND VGND VPWR VPWR _7463_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_71_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3509__B1 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6414_ _6462_/D _6435_/B _6463_/A _6651_/B VGND VGND VPWR VPWR _6420_/C sky130_fd_sc_hd__and4_4
X_3626_ _7428_/Q _5875_/A hold12/A _5704_/A _7324_/Q VGND VGND VPWR VPWR _3626_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6171__A1 _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6171__B2 _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7394_ _7578_/CLK _7394_/D fanout604/X VGND VGND VPWR VPWR _7394_/Q sky130_fd_sc_hd__dfrtp_4
X_6345_ _7048_/Q _6332_/B _6317_/C _6110_/X _7174_/Q VGND VGND VPWR VPWR _6345_/X
+ sky130_fd_sc_hd__a32o_1
X_3557_ _3511_/C _3557_/B _3557_/C VGND VGND VPWR VPWR _3557_/X sky130_fd_sc_hd__and3b_2
Xhold3102 _7036_/Q VGND VGND VPWR VPWR hold3102/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3113 _6962_/Q VGND VGND VPWR VPWR hold3113/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3124 _4260_/X VGND VGND VPWR VPWR hold3124/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6276_ _7494_/Q _6094_/A _6093_/X _6119_/X _7406_/Q VGND VGND VPWR VPWR _6276_/X
+ sky130_fd_sc_hd__a32o_1
X_3488_ _5722_/A _4449_/B _5612_/B VGND VGND VPWR VPWR _3488_/X sky130_fd_sc_hd__and3_4
Xhold3135 _4213_/X VGND VGND VPWR VPWR hold3135/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2401 _7411_/Q VGND VGND VPWR VPWR hold104/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3146 _7011_/Q VGND VGND VPWR VPWR hold3146/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4562_/D sky130_fd_sc_hd__clkbuf_2
Xhold3157 _7243_/Q VGND VGND VPWR VPWR hold3157/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2412 _7124_/Q VGND VGND VPWR VPWR hold975/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5227_ _4775_/C _4885_/X _4907_/X VGND VGND VPWR VPWR _5228_/D sky130_fd_sc_hd__a21oi_2
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2423 hold2423/A VGND VGND VPWR VPWR _5737_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3168 _7235_/Q VGND VGND VPWR VPWR hold3168/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout481_A _5735_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2434 hold939/X VGND VGND VPWR VPWR _5600_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3179 _7217_/Q VGND VGND VPWR VPWR _3797_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1700 hold1700/A VGND VGND VPWR VPWR _5927_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2445 _5756_/X VGND VGND VPWR VPWR hold733/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1711 _7253_/Q VGND VGND VPWR VPWR hold336/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2456 hold977/X VGND VGND VPWR VPWR _5764_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1722 hold41/X VGND VGND VPWR VPWR _4183_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2467 _6989_/Q VGND VGND VPWR VPWR hold662/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5158_ _5158_/A _5295_/B _5410_/A VGND VGND VPWR VPWR _5158_/X sky130_fd_sc_hd__and3_1
Xhold2478 hold2478/A VGND VGND VPWR VPWR _5607_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1733 _7533_/Q VGND VGND VPWR VPWR hold118/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1744 _7384_/Q VGND VGND VPWR VPWR hold1744/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2489 _6876_/Q VGND VGND VPWR VPWR hold963/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1755 _7469_/Q VGND VGND VPWR VPWR hold112/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1766 _5690_/X VGND VGND VPWR VPWR hold285/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6226__A2 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4109_ _7109_/Q _4084_/X _4425_/A VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__a21o_1
X_5089_ _5091_/C _5089_/B _5089_/C _5094_/A VGND VGND VPWR VPWR _5089_/Y sky130_fd_sc_hd__nand4_4
Xhold1777 _7570_/Q VGND VGND VPWR VPWR hold386/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1788 _7401_/Q VGND VGND VPWR VPWR hold402/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_168_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1799 _7314_/Q VGND VGND VPWR VPWR hold344/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5985__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3748__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_70 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6162__A1 _7521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input42_A mgmt_gpio_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6465__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5673__A0 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4476__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2990 hold722/X VGND VGND VPWR VPWR _4327_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_187_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5425__B1 _4758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5728__A1 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7215__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4460_ _4460_/A0 _5979_/A0 _4460_/S VGND VGND VPWR VPWR _4460_/X sky130_fd_sc_hd__mux2_1
Xhold307 hold307/A VGND VGND VPWR VPWR _7298_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold318 _7169_/Q VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3411_ _7554_/Q VGND VGND VPWR VPWR _3411_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6099__D _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold329 hold329/A VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_151_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4391_ _5815_/A1 hold356/X _4393_/S VGND VGND VPWR VPWR _4391_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6130_ _7472_/Q _6032_/Y _6332_/C _7488_/Q _6129_/X VGND VGND VPWR VPWR _6130_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4909__B _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A3 _4744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6061_ _7585_/Q _7584_/Q _7586_/Q _7587_/Q VGND VGND VPWR VPWR _6061_/X sky130_fd_sc_hd__a211o_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6456__A2 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 hold2598/X VGND VGND VPWR VPWR hold2599/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5328_/A _5328_/B _5013_/C VGND VGND VPWR VPWR _5012_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1018 hold2719/X VGND VGND VPWR VPWR _7335_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3532__C _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1029 hold2741/X VGND VGND VPWR VPWR hold2742/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4219__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3690__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6759__A3 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5967__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6963_ _7070_/CLK _6963_/D fanout590/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_177_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5914_ _5914_/A0 _5914_/A1 _5919_/S VGND VGND VPWR VPWR _5914_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6894_ _4127_/A1 _6894_/D _6844_/X VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfrtp_1
X_5845_ _5845_/A0 _5998_/A1 _5847_/S VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3993__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5776_ _5776_/A hold48/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7515_ _7530_/CLK _7515_/D fanout600/X VGND VGND VPWR VPWR _7515_/Q sky130_fd_sc_hd__dfrtp_4
X_4727_ _5260_/C _5387_/D VGND VGND VPWR VPWR _4727_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_133_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7446_ _7510_/CLK _7446_/D fanout603/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfrtp_4
X_4658_ _4954_/A _5248_/A _5213_/A VGND VGND VPWR VPWR _4952_/B sky130_fd_sc_hd__and3_2
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR _4142_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3609_ _3608_/X _3609_/A1 _3996_/A VGND VGND VPWR VPWR _3609_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold830 _4520_/X VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6695__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold841 hold841/A VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7377_ _7487_/CLK _7377_/D fanout593/X VGND VGND VPWR VPWR _7377_/Q sky130_fd_sc_hd__dfrtp_4
X_4589_ _4825_/A _5071_/A VGND VGND VPWR VPWR _5115_/B sky130_fd_sc_hd__and2b_4
Xhold852 hold852/A VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold863 _5774_/X VGND VGND VPWR VPWR _7381_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold874 hold874/A VGND VGND VPWR VPWR hold874/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6328_ _6312_/X _6314_/X _6327_/Y VGND VGND VPWR VPWR _6328_/X sky130_fd_sc_hd__a21bo_4
Xhold885 hold885/A VGND VGND VPWR VPWR hold885/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4819__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold896 _4274_/X VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6259_ _7285_/Q _6036_/Y _6067_/A VGND VGND VPWR VPWR _6259_/X sky130_fd_sc_hd__o21a_1
Xhold2220 _5667_/X VGND VGND VPWR VPWR hold523/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4458__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5655__A0 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2231 _7462_/Q VGND VGND VPWR VPWR hold502/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2242 hold526/X VGND VGND VPWR VPWR _5910_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2253 _5800_/X VGND VGND VPWR VPWR hold904/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2264 _5730_/X VGND VGND VPWR VPWR hold599/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1530 hold211/X VGND VGND VPWR VPWR _5944_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2275 _5784_/X VGND VGND VPWR VPWR hold583/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1541 _7514_/Q VGND VGND VPWR VPWR hold229/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2286 _7347_/Q VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2297 hold909/X VGND VGND VPWR VPWR _5809_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1552 _7508_/Q VGND VGND VPWR VPWR hold205/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1563 _7524_/Q VGND VGND VPWR VPWR hold215/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1574 hold267/X VGND VGND VPWR VPWR _5743_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3681__A2 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1585 hold20/X VGND VGND VPWR VPWR _3576_/C sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5407__B1 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1596 _7313_/Q VGND VGND VPWR VPWR hold265/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5958__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4630__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4570__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5186__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3617__C _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6686__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5894__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6438__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5646__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4745__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5949__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6610__A2 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3960_ _7122_/Q _3665_/X _3952_/X _3954_/X _3959_/X VGND VGND VPWR VPWR _3961_/D
+ sky130_fd_sc_hd__a2111o_4
XFILLER_0_57_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3891_ _7193_/Q _4545_/A _3669_/X _6968_/Q _3890_/X VGND VGND VPWR VPWR _3891_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5630_ _5630_/A0 _5948_/A1 _5630_/S VGND VGND VPWR VPWR _5630_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5177__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4911__C _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4385__A0 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5561_ _5563_/A1 _4814_/Y _5471_/X _5278_/B VGND VGND VPWR VPWR _5562_/D sky130_fd_sc_hd__o31a_1
XFILLER_0_170_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7300_ _7501_/CLK _7300_/D fanout582/X VGND VGND VPWR VPWR _7300_/Q sky130_fd_sc_hd__dfrtp_4
X_4512_ _4512_/A0 _5815_/A1 _4514_/S VGND VGND VPWR VPWR _4512_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6126__A1 _7528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3527__C _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5492_ _5486_/Y _5488_/Y _5532_/B _5492_/D VGND VGND VPWR VPWR _5492_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6126__B2 _7480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold104 hold104/A VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_80_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold115 hold115/A VGND VGND VPWR VPWR _7573_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7231_ _7231_/CLK _7231_/D _4128_/B VGND VGND VPWR VPWR _7231_/Q sky130_fd_sc_hd__dfrtp_4
Xhold126 hold126/A VGND VGND VPWR VPWR hold126/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6677__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4443_ _4443_/A0 _5986_/A1 _4448_/S VGND VGND VPWR VPWR _4443_/X sky130_fd_sc_hd__mux2_1
Xhold137 hold137/A VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold148 hold148/A VGND VGND VPWR VPWR _7443_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold159 hold159/A VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4374_ _5852_/A0 _4374_/A1 _4375_/S VGND VGND VPWR VPWR _4374_/X sky130_fd_sc_hd__mux2_1
X_7162_ _7212_/CLK _7162_/D fanout573/X VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout606 input75/X VGND VGND VPWR VPWR fanout606/X sky130_fd_sc_hd__buf_12
XANTENNA__3543__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout617 _4879_/C VGND VGND VPWR VPWR _5282_/A sky130_fd_sc_hd__buf_12
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6113_ _7367_/Q _6144_/C _6084_/X _6112_/X _7479_/Q VGND VGND VPWR VPWR _6113_/X
+ sky130_fd_sc_hd__a32o_1
X_7093_ _7096_/CLK _7093_/D fanout604/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__A0 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4358__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _7594_/Q _7593_/Q VGND VGND VPWR VPWR _6467_/A sky130_fd_sc_hd__and2b_4
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6601__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6946_ _7577_/CLK _6946_/D fanout583/X VGND VGND VPWR VPWR _7652_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__6870__A _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4612__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3966__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6877_ _7201_/CLK _6877_/D _6833_/A VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5828_ _5828_/A0 _5999_/A1 _5829_/S VGND VGND VPWR VPWR _5828_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout611_A _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4821__C _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3718__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5759_ _5993_/A1 _5759_/A1 _5766_/S VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_134_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6117__A1 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6117__B2 _7311_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6668__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7429_ _7429_/CLK _7429_/D fanout583/X VGND VGND VPWR VPWR _7429_/Q sky130_fd_sc_hd__dfrtp_4
Xhold660 hold660/A VGND VGND VPWR VPWR hold660/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold671 _4493_/X VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold682 hold682/A VGND VGND VPWR VPWR hold682/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold693 _5862_/X VGND VGND VPWR VPWR _7459_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input144_A wb_dat_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2050 _4483_/X VGND VGND VPWR VPWR hold491/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4300__A0 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2061 _5849_/X VGND VGND VPWR VPWR _7447_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2072 hold83/X VGND VGND VPWR VPWR hold2072/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2083 _4413_/X VGND VGND VPWR VPWR hold715/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2094 hold775/X VGND VGND VPWR VPWR _4415_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1360 _6786_/B VGND VGND VPWR VPWR hold2840/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1371 hold1410/X VGND VGND VPWR VPWR hold1411/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1382 _7346_/Q VGND VGND VPWR VPWR _5735_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1393 hold2/X VGND VGND VPWR VPWR _4256_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5800__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput209 _3439_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XANTENNA__6659__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5331__A2 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3893__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4090_ _4564_/C _4564_/D _4563_/A _4563_/B VGND VGND VPWR VPWR _4095_/B sky130_fd_sc_hd__nor4_1
XANTENNA__5095__A1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6292__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4906__C _5185_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6800_ _7109_/Q _6800_/A2 _6800_/B1 _4426_/Y _6799_/X VGND VGND VPWR VPWR _6800_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5398__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4992_ _5038_/A _5183_/A _5038_/B _5053_/C VGND VGND VPWR VPWR _4992_/Y sky130_fd_sc_hd__nand4_1
X_6731_ _7004_/Q _6419_/D _6446_/X _7190_/Q VGND VGND VPWR VPWR _6731_/X sky130_fd_sc_hd__a22o_1
X_3943_ input71/X _4231_/S _3934_/X _3935_/X _3942_/X VGND VGND VPWR VPWR _3961_/A
+ sky130_fd_sc_hd__a2111o_4
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4414__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6662_ _6874_/Q _6447_/C _6459_/C _6661_/X VGND VGND VPWR VPWR _6662_/X sky130_fd_sc_hd__a31o_1
X_3874_ _7280_/Q _5947_/A _5659_/B _3598_/X VGND VGND VPWR VPWR _3879_/B sky130_fd_sc_hd__a31o_2
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5613_ _5613_/A0 _5948_/A1 _5613_/S VGND VGND VPWR VPWR _5613_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3538__B _3569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6593_ _7548_/Q _6419_/A _6419_/C _7564_/Q _6592_/X VGND VGND VPWR VPWR _6593_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_171_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5544_ _5453_/C _5180_/B _5248_/B _5453_/A VGND VGND VPWR VPWR _5545_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3581__B2 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ _4722_/Y _4748_/Y _4806_/Y _5563_/A1 VGND VGND VPWR VPWR _5476_/C sky130_fd_sc_hd__a211o_1
XANTENNA__5858__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7214_ _4150_/A1 _7214_/D _6866_/X VGND VGND VPWR VPWR _7214_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4426_ _7109_/Q _7110_/Q _7111_/Q VGND VGND VPWR VPWR _4426_/Y sky130_fd_sc_hd__nor3_2
Xfanout403 wire406/X VGND VGND VPWR VPWR _4212_/A sky130_fd_sc_hd__buf_12
X_7145_ _7266_/CLK _7145_/D fanout567/X VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout414 hold71/X VGND VGND VPWR VPWR _5830_/C sky130_fd_sc_hd__buf_8
Xfanout425 _4861_/X VGND VGND VPWR VPWR _5038_/B sky130_fd_sc_hd__buf_6
X_4357_ _4357_/A0 _5586_/A0 _4357_/S VGND VGND VPWR VPWR _4357_/X sky130_fd_sc_hd__mux2_1
Xfanout436 _6093_/X VGND VGND VPWR VPWR _6332_/C sky130_fd_sc_hd__buf_12
XANTENNA__3884__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout447 _6072_/B VGND VGND VPWR VPWR _6144_/A sky130_fd_sc_hd__buf_12
Xfanout458 _4705_/Y VGND VGND VPWR VPWR _5451_/A1 sky130_fd_sc_hd__buf_8
X_7076_ _7096_/CLK _7076_/D fanout605/X VGND VGND VPWR VPWR _7656_/A sky130_fd_sc_hd__dfrtp_1
Xfanout469 hold61/X VGND VGND VPWR VPWR _5999_/A1 sky130_fd_sc_hd__buf_4
X_4288_ _3607_/Y _4288_/A1 _4289_/S VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_4_14__f_wb_clk_i clkbuf_3_7_0_wb_clk_i/X VGND VGND VPWR VPWR _7646_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6283__B1 _6281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6027_ _7589_/Q _7588_/Q _6106_/B VGND VGND VPWR VPWR _6027_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout561_A _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4816__C _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _7601_/CLK _6929_/D _6865_/A VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfstp_4
Xclkbuf_leaf_31_csclk _7267_/CLK VGND VGND VPWR VPWR _7565_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3939__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4551__C _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_csclk _7496_/CLK VGND VGND VPWR VPWR _7581_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_161_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3572__A1 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5849__A0 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold490 hold490/A VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3875__A2 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6274__B1 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3627__A2 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1190 hold1190/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
XFILLER_0_150_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6577__A1 _7484_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6577__B2 _7324_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4742__B _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4234__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4461__C _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4180__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3590_ _7477_/Q _5875_/A _3590_/C VGND VGND VPWR VPWR _3590_/X sky130_fd_sc_hd__and3_1
XANTENNA__5552__A2 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5260_ _5260_/A _5260_/B _5260_/C _5260_/D VGND VGND VPWR VPWR _5260_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__6501__A1 _7529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6501__B2 _7289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4211_ _4211_/A0 _5955_/A1 _4211_/S VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
X_5191_ _4929_/A _5180_/A _5180_/B _5035_/C VGND VGND VPWR VPWR _5191_/X sky130_fd_sc_hd__a31o_1
Xhold2808 _6979_/Q VGND VGND VPWR VPWR _4289_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2819 hold2819/A VGND VGND VPWR VPWR hold2819/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3866__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4142_ _4142_/A _4142_/B VGND VGND VPWR VPWR _4142_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__6265__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4073_ hold4/A hold7/A _4075_/S VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4409__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3618__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6568__B2 _7515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4975_ _4984_/B _4984_/A _4660_/Y _4672_/X VGND VGND VPWR VPWR _4975_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5240__B2 _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3549__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6714_ _6990_/Q _6420_/B _6706_/X _6710_/X _6713_/X VGND VGND VPWR VPWR _6714_/X
+ sky130_fd_sc_hd__a2111o_1
X_3926_ _6874_/Q _5875_/A _5632_/B _3494_/X _7471_/Q VGND VGND VPWR VPWR _3926_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6645_ _7438_/Q _6747_/B _6645_/C VGND VGND VPWR VPWR _6645_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3857_ _3924_/A1 _3856_/A _7073_/Q _6893_/Q VGND VGND VPWR VPWR _3857_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_15_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6576_ _7380_/Q _6408_/B _6423_/X _7332_/Q _6575_/X VGND VGND VPWR VPWR _6576_/X
+ sky130_fd_sc_hd__a221o_1
X_3788_ _7170_/Q _3647_/X _4340_/A _7019_/Q _3787_/X VGND VGND VPWR VPWR _3788_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3554__A1 _4176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3554__B2 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5527_ hold130/A _5580_/A2 _5560_/B _5526_/X _5515_/X VGND VGND VPWR VPWR _7206_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5458_ _5107_/A _5248_/A _5094_/A _5252_/B VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__a31o_1
X_4409_ _4409_/A0 _4408_/X _4423_/S VGND VGND VPWR VPWR _4409_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5389_ _4601_/Y _4700_/Y _4844_/Y _4789_/Y VGND VGND VPWR VPWR _5518_/C sky130_fd_sc_hd__a31o_1
X_7128_ _7395_/CLK _7128_/D fanout598/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold187_A _7492_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4319__S _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7496__SET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7059_ _7190_/CLK _7059_/D fanout573/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4795__A_N _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6271__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4282__A2 _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__A1 _7323_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__B2 _7363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A wb_adr_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input72_A mgmt_gpio_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5298__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3848__A2 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6247__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4229__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5470__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4760_ _5139_/D _4760_/B _4760_/C _4760_/D VGND VGND VPWR VPWR _4763_/C sky130_fd_sc_hd__nand4_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4191__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3784__A1 _7538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3711_ input24/X _3488_/X _3707_/X _3708_/X _3710_/X VGND VGND VPWR VPWR _3711_/X
+ sky130_fd_sc_hd__a2111o_2
XANTENNA__3784__B2 _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4691_ _5038_/A _4758_/B _5328_/B VGND VGND VPWR VPWR _5297_/A sky130_fd_sc_hd__and3_2
XANTENNA_clkbuf_leaf_24_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6430_ _6431_/A _6431_/B _6431_/C VGND VGND VPWR VPWR _6430_/X sky130_fd_sc_hd__and3_4
X_3642_ _3642_/A _3642_/B _3642_/C _3642_/D VGND VGND VPWR VPWR _3643_/C sky130_fd_sc_hd__nor4_2
XFILLER_0_102_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6722__A1 _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5525__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6722__B2 _7154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6361_ _7039_/Q _6111_/X _6121_/X _6991_/Q _6360_/X VGND VGND VPWR VPWR _6362_/C
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3573_ _3572_/X _3573_/A1 _3996_/A VGND VGND VPWR VPWR _7221_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_113_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2441_A _7316_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2539_A _7178_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5312_ _4667_/A _4692_/Y _4768_/Y _4796_/Y _4755_/Y VGND VGND VPWR VPWR _5312_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3535__C _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6292_ _7197_/Q _6332_/B _6079_/X _6094_/X _7209_/Q VGND VGND VPWR VPWR _6292_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6486__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5243_ _5248_/B _5453_/A _5243_/C VGND VGND VPWR VPWR _5367_/B sky130_fd_sc_hd__and3_1
Xhold2605 _7429_/Q VGND VGND VPWR VPWR hold850/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2616 hold854/X VGND VGND VPWR VPWR _5747_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2627 _6953_/Q VGND VGND VPWR VPWR hold647/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5174_ _5282_/A _5011_/B _5183_/C VGND VGND VPWR VPWR _5174_/Y sky130_fd_sc_hd__a21oi_4
Xhold2638 hold639/X VGND VGND VPWR VPWR _5988_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2649 hold688/X VGND VGND VPWR VPWR _5970_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1904 hold293/X VGND VGND VPWR VPWR _7354_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1915 hold114/X VGND VGND VPWR VPWR _5990_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4139__S _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1926 _7474_/Q VGND VGND VPWR VPWR hold1926/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4125_ input84/X _4168_/D _6897_/Q VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_2
Xhold1937 _5618_/X VGND VGND VPWR VPWR hold391/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1948 _4188_/X VGND VGND VPWR VPWR hold467/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1959 _4513_/X VGND VGND VPWR VPWR hold425/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6253__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4056_ _6910_/Q _6909_/Q _6908_/Q _7071_/Q VGND VGND VPWR VPWR _4057_/S sky130_fd_sc_hd__and4bb_1
XFILLER_0_78_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout357_A _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4382__B _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4958_ _4958_/A _4958_/B _4958_/C VGND VGND VPWR VPWR _4962_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_148_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3775__A1 _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3775__B2 _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3909_ _6963_/Q _5632_/B _5659_/B _5794_/A _7400_/Q VGND VGND VPWR VPWR _3909_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4972__B1 _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4889_ _4889_/A _4889_/B VGND VGND VPWR VPWR _4891_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6628_ _7310_/Q _6420_/B _6463_/X _7430_/Q _6627_/X VGND VGND VPWR VPWR _6628_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_172_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6559_ _7323_/Q _6421_/X _6462_/X _7363_/Q _6558_/X VGND VGND VPWR VPWR _6559_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_hold1541_A _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6477__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4557__B _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6229__B1 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6099__A_N _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_179_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3766__A1 _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6704__A1 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire453 _4743_/Y VGND VGND VPWR VPWR _4755_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6180__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4748__A _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__A _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6483__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4467__B _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5443__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6640__B1 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5930_ hold464/X _5930_/A1 _5937_/S VGND VGND VPWR VPWR _5930_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4914__C _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5861_ _5987_/A1 _5861_/A1 _5865_/S VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7600_ _7601_/CLK _7600_/D fanout567/X VGND VGND VPWR VPWR _7600_/Q sky130_fd_sc_hd__dfrtp_1
X_4812_ _4812_/A _4812_/B _4812_/C VGND VGND VPWR VPWR _4818_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_185_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2489_A _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5792_ _5792_/A0 _5999_/A1 _5793_/S VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7531_ _7560_/CLK _7531_/D fanout599/X VGND VGND VPWR VPWR _7531_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3757__B2 _7578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4743_ _4743_/A _4856_/A _5073_/B VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4422__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7462_ _7580_/CLK _7462_/D fanout594/X VGND VGND VPWR VPWR _7462_/Q sky130_fd_sc_hd__dfrtp_2
X_4674_ _5071_/A _4675_/A _4675_/B _4675_/C VGND VGND VPWR VPWR _4679_/C sky130_fd_sc_hd__nand4_4
XFILLER_0_114_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6413_ _6434_/B _6747_/C _6413_/C VGND VGND VPWR VPWR _6420_/B sky130_fd_sc_hd__and3_4
XFILLER_0_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3625_ _7460_/Q _5857_/A _5929_/A _7524_/Q _3624_/X VGND VGND VPWR VPWR _3632_/A
+ sky130_fd_sc_hd__a221o_1
X_7393_ _7471_/CLK _7393_/D fanout593/X VGND VGND VPWR VPWR _7393_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6171__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4182__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6344_ _7038_/Q _6121_/C _6084_/X _6112_/X _6876_/Q VGND VGND VPWR VPWR _6344_/X
+ sky130_fd_sc_hd__a32o_1
X_3556_ hold36/X _5722_/A _5731_/B VGND VGND VPWR VPWR _5704_/A sky130_fd_sc_hd__and3_4
Xhold3103 hold3103/A VGND VGND VPWR VPWR _4365_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3114 hold3114/A VGND VGND VPWR VPWR _4266_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6275_ _7470_/Q _6087_/X _6094_/X _7510_/Q _6274_/X VGND VGND VPWR VPWR _6280_/B
+ sky130_fd_sc_hd__a221o_1
X_3487_ _7406_/Q _5794_/A _3486_/X input10/X _3479_/X VGND VGND VPWR VPWR _3487_/X
+ sky130_fd_sc_hd__a221o_2
Xhold3125 _7222_/Q VGND VGND VPWR VPWR hold3125/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3136 _7061_/Q VGND VGND VPWR VPWR hold3136/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3562__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2402 hold104/X VGND VGND VPWR VPWR _5808_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3147 hold3147/A VGND VGND VPWR VPWR _4335_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4562_/C sky130_fd_sc_hd__clkbuf_2
Xhold3158 hold3158/A VGND VGND VPWR VPWR _5613_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2413 hold975/X VGND VGND VPWR VPWR _4464_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5226_ _4933_/B _5213_/C _5342_/B _5102_/B _5357_/B2 VGND VGND VPWR VPWR _5226_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5131__B1 _5028_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6474__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2424 _7293_/Q VGND VGND VPWR VPWR hold718/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3169 hold3169/A VGND VGND VPWR VPWR _5604_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5682__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2435 _5600_/X VGND VGND VPWR VPWR hold940/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1701 _5927_/X VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2446 _7393_/Q VGND VGND VPWR VPWR hold933/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2457 _6991_/Q VGND VGND VPWR VPWR hold973/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1712 hold336/X VGND VGND VPWR VPWR _5627_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1723 _4183_/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2468 hold662/X VGND VGND VPWR VPWR _4305_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5157_ _5387_/C _4815_/B _5453_/B _4977_/X _4823_/B VGND VGND VPWR VPWR _5160_/C
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout474_A hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1734 hold118/X VGND VGND VPWR VPWR _5945_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2479 _6958_/Q VGND VGND VPWR VPWR hold658/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1745 hold1745/A VGND VGND VPWR VPWR _5778_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4108_ _6751_/S _6427_/A _4105_/B _4107_/Y _4100_/X VGND VGND VPWR VPWR _6932_/D
+ sky130_fd_sc_hd__a41o_1
Xhold1756 hold112/X VGND VGND VPWR VPWR _5873_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1767 hold285/X VGND VGND VPWR VPWR _7306_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5088_ _5222_/A _5086_/B _5087_/Y VGND VGND VPWR VPWR _5088_/Y sky130_fd_sc_hd__a21oi_1
Xhold1778 hold386/X VGND VGND VPWR VPWR _5987_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1789 hold402/X VGND VGND VPWR VPWR _5797_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4039_ _4039_/A0 _4038_/X _4040_/A VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_177_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1589_A _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4840__B _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3737__A _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_60 _6212_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4568__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3920__B2 _7260_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3472__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input35_A mask_rev_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3684__B1 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2980 _4535_/X VGND VGND VPWR VPWR hold2980/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2991 _7352_/Q VGND VGND VPWR VPWR hold2991/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_89_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5425__A1 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5399__A _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3987__A1 _7287_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3739__A1 _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3647__A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4242__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7069__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6689__B1 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold308 hold308/A VGND VGND VPWR VPWR hold308/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold319 hold319/A VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4164__A1 _4164_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4390_ _5583_/A0 _4390_/A1 _4393_/S VGND VGND VPWR VPWR _4390_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5581__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _6060_/A1 _6019_/Y _6059_/X _6051_/C VGND VGND VPWR VPWR _7598_/D sky130_fd_sc_hd__a22o_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5664__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1008 hold2825/X VGND VGND VPWR VPWR hold2826/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_84_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5011_ _5011_/A _5011_/B _5328_/B _5328_/A VGND VGND VPWR VPWR _5011_/Y sky130_fd_sc_hd__nand4_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 hold2779/X VGND VGND VPWR VPWR hold2780/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5801__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6208__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6613__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3690__A3 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4417__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6962_ _7268_/CLK _6962_/D fanout572/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5913_ _5913_/A0 _5985_/A1 _5919_/S VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__mux2_1
X_6893_ _4127_/A1 _6893_/D _6843_/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5844_ _5844_/A0 _5979_/A0 _5847_/S VGND VGND VPWR VPWR _5844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5775_ _5775_/A0 hold17/X _5775_/S VGND VGND VPWR VPWR _5775_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6392__A2 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7514_ _7565_/CLK _7514_/D fanout602/X VGND VGND VPWR VPWR _7514_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_161_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4726_ _5222_/B _4726_/B _4726_/C _5005_/A VGND VGND VPWR VPWR _4726_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_44_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7445_ _7522_/CLK _7445_/D fanout605/X VGND VGND VPWR VPWR _7445_/Q sky130_fd_sc_hd__dfrtp_4
X_4657_ _4657_/A _4657_/B _4657_/C _4657_/D VGND VGND VPWR VPWR _5248_/B sky130_fd_sc_hd__and4_4
XFILLER_0_140_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4155__A1 _4135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_2
X_3608_ _7219_/Q _3607_/Y _3923_/S VGND VGND VPWR VPWR _3608_/X sky130_fd_sc_hd__mux2_1
Xhold820 _5586_/X VGND VGND VPWR VPWR _7213_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_4
X_7376_ _7563_/CLK _7376_/D fanout599/X VGND VGND VPWR VPWR _7376_/Q sky130_fd_sc_hd__dfstp_4
X_4588_ _4562_/Y _4585_/Y _4593_/A _5071_/A VGND VGND VPWR VPWR _5295_/A sky130_fd_sc_hd__a2bb2o_4
Xhold831 hold831/A VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap550 _4608_/Y VGND VGND VPWR VPWR _4869_/A2 sky130_fd_sc_hd__buf_6
Xhold842 _5711_/X VGND VGND VPWR VPWR _7325_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3902__A1 _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold853 _4454_/X VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold864 hold864/A VGND VGND VPWR VPWR hold864/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6327_ _6327_/A _6327_/B _6327_/C _6327_/D VGND VGND VPWR VPWR _6327_/Y sky130_fd_sc_hd__nor4_1
Xhold875 hold875/A VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3539_ _7430_/Q _3537_/X _5929_/A _7526_/Q _3536_/X VGND VGND VPWR VPWR _3539_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout591_A fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmgmt_gpio_15_buff_inst _4161_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_8
Xhold886 _5646_/X VGND VGND VPWR VPWR _7267_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold897 hold897/A VGND VGND VPWR VPWR hold897/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6258_ _6243_/X _6245_/X _6257_/Y VGND VGND VPWR VPWR _6258_/X sky130_fd_sc_hd__a21bo_2
XFILLER_0_110_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2210 _5694_/X VGND VGND VPWR VPWR hold515/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2221 hold523/X VGND VGND VPWR VPWR _7286_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2232 hold502/X VGND VGND VPWR VPWR _5865_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5209_ _4943_/B _4915_/C _4946_/Y _4774_/Y VGND VGND VPWR VPWR _5228_/A sky130_fd_sc_hd__o2bb2a_1
Xhold2243 _5910_/X VGND VGND VPWR VPWR hold527/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2254 _7312_/Q VGND VGND VPWR VPWR hold604/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6189_ _6181_/X _6094_/A _6186_/X _6184_/X _6188_/X VGND VGND VPWR VPWR _6189_/X
+ sky130_fd_sc_hd__a2111o_4
Xhold1520 hold217/X VGND VGND VPWR VPWR _4443_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2265 hold599/X VGND VGND VPWR VPWR _7342_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2276 _7574_/Q VGND VGND VPWR VPWR hold516/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1531 _5944_/X VGND VGND VPWR VPWR hold212/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1542 hold229/X VGND VGND VPWR VPWR _5924_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2287 hold86/X VGND VGND VPWR VPWR _5736_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1553 hold205/X VGND VGND VPWR VPWR _5917_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2298 _7324_/Q VGND VGND VPWR VPWR hold901/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1564 hold215/X VGND VGND VPWR VPWR _5935_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5407__A1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1575 _5743_/X VGND VGND VPWR VPWR hold268/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1586 _3502_/X VGND VGND VPWR VPWR _4455_/C sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1597 hold265/X VGND VGND VPWR VPWR _5698_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_156_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_168_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5947__A _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7509__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6383__A2 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6135__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6686__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4298__A _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4879__A_N _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4237__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3890_ _7178_/Q _5938_/C _5619_/B _3525_/X _7432_/Q VGND VGND VPWR VPWR _3890_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_156_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6374__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5582__A0 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5295__C _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5560_ _5560_/A _5560_/B _5560_/C VGND VGND VPWR VPWR _5560_/X sky130_fd_sc_hd__and3_1
XFILLER_0_170_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4511_ _4511_/A0 _5583_/A0 _4514_/S VGND VGND VPWR VPWR _4511_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6126__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5491_ _5491_/A _5531_/B _5491_/C _5531_/C VGND VGND VPWR VPWR _5492_/D sky130_fd_sc_hd__and4_1
XFILLER_0_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold105 _5808_/X VGND VGND VPWR VPWR _7411_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7230_ _7255_/CLK _7230_/D _4128_/B VGND VGND VPWR VPWR _7230_/Q sky130_fd_sc_hd__dfstp_4
X_4442_ _4442_/A0 _5985_/A1 _4448_/S VGND VGND VPWR VPWR _4442_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold116 hold116/A VGND VGND VPWR VPWR hold116/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold127 _4532_/X VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold138 _5700_/X VGND VGND VPWR VPWR _7315_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5885__A1 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold149 hold149/A VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_186_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7161_ _7191_/CLK _7161_/D _6871_/A VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_4
X_4373_ _5914_/A1 _4373_/A1 _4375_/S VGND VGND VPWR VPWR _4373_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3896__B1 _3862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2521_A _7360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6119_/B _6144_/A _6112_/C _6112_/D VGND VGND VPWR VPWR _6112_/X sky130_fd_sc_hd__and4b_4
Xfanout607 _6780_/B VGND VGND VPWR VPWR _4309_/B sky130_fd_sc_hd__buf_12
Xfanout618 _4945_/A VGND VGND VPWR VPWR _4879_/C sky130_fd_sc_hd__buf_12
XANTENNA__3543__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7092_ _7510_/CLK _7092_/D fanout603/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4358__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13__f_wb_clk_i clkbuf_3_6_0_wb_clk_i/X VGND VGND VPWR VPWR _4164_/A1 sky130_fd_sc_hd__clkbuf_16
X_6043_ _7594_/Q _7593_/Q VGND VGND VPWR VPWR _6424_/C sky130_fd_sc_hd__nor2_8
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _7429_/CLK _6945_/D fanout583/X VGND VGND VPWR VPWR _7651_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5767__A _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6876_ _7201_/CLK _6876_/D _6833_/A VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__3820__B1 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5827_ _5827_/A0 _5863_/A0 _5829_/S VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_162_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6365__A2 _6072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5758_ _5758_/A hold48/X VGND VGND VPWR VPWR _5766_/S sky130_fd_sc_hd__nand2_8
XANTENNA_fanout604_A fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4709_ _4887_/B _4879_/C _5387_/B VGND VGND VPWR VPWR _4709_/Y sky130_fd_sc_hd__nand3_4
XANTENNA_clkbuf_leaf_72_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6117__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5689_ _5896_/A0 _5689_/A1 _5694_/S VGND VGND VPWR VPWR _5689_/X sky130_fd_sc_hd__mux2_1
X_7428_ _7582_/CLK _7428_/D fanout584/X VGND VGND VPWR VPWR _7428_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5325__B1 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6668__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5876__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7359_ _7359_/CLK _7359_/D fanout575/X VGND VGND VPWR VPWR _7359_/Q sky130_fd_sc_hd__dfstp_2
Xhold650 hold650/A VGND VGND VPWR VPWR _7255_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold661 _4193_/X VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6110__B _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold672 hold672/A VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1621_A _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold683 hold683/A VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5007__A _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold694 hold694/A VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5628__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4846__A _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2040 hold2040/A VGND VGND VPWR VPWR hold464/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2051 _7069_/Q VGND VGND VPWR VPWR hold384/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2062 _7649_/A VGND VGND VPWR VPWR hold682/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2073 _5898_/X VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input137_A wb_dat_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2084 _7668_/A VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2095 _4415_/X VGND VGND VPWR VPWR hold776/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1350 _4321_/A1 VGND VGND VPWR VPWR hold2863/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1361 _6783_/A1 VGND VGND VPWR VPWR hold2896/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1372 hold1577/X VGND VGND VPWR VPWR hold1578/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 hold1404/X VGND VGND VPWR VPWR hold1405/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1394 _4256_/X VGND VGND VPWR VPWR hold1394/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6780__B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5677__A hold12/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4581__A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4367__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3575__C1 _3574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4119__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5867__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3893__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4756__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3660__A _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6292__A1 _7197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2102_A _7443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4991_ _5183_/A _5203_/B _5038_/B _5158_/A VGND VGND VPWR VPWR _5037_/B sky130_fd_sc_hd__nand4_1
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6595__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5398__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5587__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6730_ _7150_/Q _6408_/A _6420_/A _6970_/Q _6729_/X VGND VGND VPWR VPWR _6730_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4491__A _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3942_ input61/X _5643_/A _3938_/X _3939_/X _3941_/X VGND VGND VPWR VPWR _3942_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3802__B1 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6661_ _6967_/Q _6420_/A _6421_/X _7006_/Q _6660_/X VGND VGND VPWR VPWR _6661_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6347__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3873_ _7544_/Q _3519_/X _3866_/X _3868_/X _3872_/X VGND VGND VPWR VPWR _3879_/A
+ sky130_fd_sc_hd__a2111o_4
XFILLER_0_190_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5612_ hold36/X _5612_/B _5612_/C _5640_/D VGND VGND VPWR VPWR _5613_/S sky130_fd_sc_hd__and4_1
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3538__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6592_ _7468_/Q _6434_/B _6574_/C _6466_/X _7508_/Q VGND VGND VPWR VPWR _6592_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_144_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5543_ _5543_/A _5543_/B _5543_/C VGND VGND VPWR VPWR _5543_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3581__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5474_ _5521_/B _5564_/B _5474_/C _5518_/A VGND VGND VPWR VPWR _5478_/A sky130_fd_sc_hd__nand4_1
X_7213_ _7213_/CLK _7213_/D fanout590/X VGND VGND VPWR VPWR _7213_/Q sky130_fd_sc_hd__dfrtp_4
X_4425_ _4425_/A _4425_/B _4425_/C _4424_/Y VGND VGND VPWR VPWR _4430_/B sky130_fd_sc_hd__nor4b_2
X_7144_ _7144_/CLK _7144_/D fanout567/X VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4530__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4356_ _4356_/A0 _5852_/A0 _4357_/S VGND VGND VPWR VPWR _4356_/X sky130_fd_sc_hd__mux2_1
Xfanout415 _5938_/B VGND VGND VPWR VPWR _5640_/B sky130_fd_sc_hd__buf_12
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout437 _6078_/X VGND VGND VPWR VPWR _6120_/B sky130_fd_sc_hd__buf_12
Xfanout448 _4859_/C VGND VGND VPWR VPWR _5183_/C sky130_fd_sc_hd__buf_12
X_7075_ _7075_/CLK _7075_/D _6865_/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_2
X_4287_ _3643_/Y _4287_/A1 _4289_/S VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout387_A _5911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6026_ _6051_/C _6929_/Q _7589_/Q _6025_/Y VGND VGND VPWR VPWR _7589_/D sky130_fd_sc_hd__o31a_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6586__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__A3 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6440__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6928_ _7363_/CLK _6928_/D fanout575/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold132_A _3519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6859_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6859_/X sky130_fd_sc_hd__and2_1
XANTENNA__6338__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4551__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4349__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1669_A _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6121__A _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6510__A2 _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold480 hold480/A VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold491 hold491/A VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3875__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4576__A _4615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6274__A1 _7518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1180 hold1180/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1191 hold2824/X VGND VGND VPWR VPWR hold1191/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6577__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6329__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4461__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3655__A _7672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6031__A _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6501__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4210_ _4210_/A0 _5954_/A1 _4211_/S VGND VGND VPWR VPWR _4210_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4512__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5190_ _5030_/C _5188_/X _5189_/X _5187_/X VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__a211o_1
Xhold2809 hold2809/A VGND VGND VPWR VPWR hold2809/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4141_ _7578_/Q _4142_/A _4140_/Y VGND VGND VPWR VPWR _4141_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__4917__C _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6265__B2 _7334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4072_ hold82/A hold4/A _4075_/S VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_20_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3618__A3 _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4597__A_N _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6568__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4974_ _4996_/A _4974_/B _4974_/C _4974_/D VGND VGND VPWR VPWR _5342_/C sky130_fd_sc_hd__and4_1
XFILLER_0_176_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7073__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5240__A2 _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6713_ _7003_/Q _6455_/B _6574_/B _6651_/B _6712_/X VGND VGND VPWR VPWR _6713_/X
+ sky130_fd_sc_hd__a41o_1
X_3925_ _7046_/Q _5830_/C _5947_/B _4388_/B VGND VGND VPWR VPWR _3925_/X sky130_fd_sc_hd__and4_1
XFILLER_0_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6644_ _7502_/Q _6447_/C _6429_/X _6420_/C _7398_/Q VGND VGND VPWR VPWR _6644_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_128_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3856_ _3856_/A _3856_/B VGND VGND VPWR VPWR _3856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6575_ _7356_/Q _6413_/C _6459_/C _6462_/X _7364_/Q VGND VGND VPWR VPWR _6575_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3787_ _7247_/Q _5947_/A _3519_/B _3515_/X _7238_/Q VGND VGND VPWR VPWR _3787_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3565__A hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6740__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3554__A2 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5526_ _5038_/A _4846_/B _5118_/C _5525_/X VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_112_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5457_ _5457_/A _5457_/B VGND VGND VPWR VPWR _5457_/Y sky130_fd_sc_hd__nand2_1
X_4408_ _4441_/A0 _5993_/A1 _4422_/S VGND VGND VPWR VPWR _4408_/X sky130_fd_sc_hd__mux2_1
X_5388_ _5091_/A _5260_/C _5387_/D _5081_/A _5387_/X VGND VGND VPWR VPWR _5521_/A
+ sky130_fd_sc_hd__a41oi_4
XANTENNA_clkbuf_0__1111__A _3733_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7127_ _7395_/CLK _7127_/D fanout598/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_4
X_4339_ _4339_/A0 _5586_/A0 _4339_/S VGND VGND VPWR VPWR _4339_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6256__A1 _7533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4827__C _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7058_ _7189_/CLK _7058_/D fanout572/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfstp_1
X_6009_ _6932_/Q _6751_/S VGND VGND VPWR VPWR _6009_/Y sky130_fd_sc_hd__nor2_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__A2 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6116__A _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1953_A _7034_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6731__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_190_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input65_A mgmt_gpio_in[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6786__A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5298__A2 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3848__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6247__B2 _7309_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4245__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _7579_/Q _3501_/X _4248_/S _4150_/A1 _3709_/X VGND VGND VPWR VPWR _3710_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_28_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3784__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4690_ _5328_/A _5328_/B VGND VGND VPWR VPWR _4690_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3641_ _7372_/Q _5758_/A _3527_/X _6916_/Q _3640_/X VGND VGND VPWR VPWR _3642_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6183__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6722__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6360_ _7009_/Q _6144_/C _6081_/X _6097_/X _7185_/Q VGND VGND VPWR VPWR _6360_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3536__A2 _3496_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5930__A0 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3572_ _3609_/A1 _3570_/Y _3923_/S VGND VGND VPWR VPWR _3572_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5311_ _5311_/A _5311_/B _5488_/A VGND VGND VPWR VPWR _5314_/A sky130_fd_sc_hd__and3_1
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6291_ _7061_/Q _6032_/Y _6081_/X _7192_/Q _6290_/X VGND VGND VPWR VPWR _6291_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5804__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5289__A2 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6486__B2 _7288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5242_ _5222_/A _5248_/B _5453_/A _4941_/B VGND VGND VPWR VPWR _5545_/A sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_30_csclk _7267_/CLK VGND VGND VPWR VPWR _7530_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2606 hold850/X VGND VGND VPWR VPWR _5828_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2617 _7477_/Q VGND VGND VPWR VPWR hold870/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5173_ _4605_/Y _5528_/A3 _5046_/A _5046_/B _4690_/Y VGND VGND VPWR VPWR _5173_/X
+ sky130_fd_sc_hd__o32a_1
Xhold2628 hold647/X VGND VGND VPWR VPWR _4255_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2639 _7387_/Q VGND VGND VPWR VPWR hold637/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1905 _7549_/Q VGND VGND VPWR VPWR hold1905/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5105__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4124_ _4005_/C _4123_/B _4123_/Y _4124_/B2 VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__a22o_1
Xhold1916 _5990_/X VGND VGND VPWR VPWR hold115/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1927 hold1927/A VGND VGND VPWR VPWR _5879_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1938 _7402_/Q VGND VGND VPWR VPWR hold360/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1949 _7125_/Q VGND VGND VPWR VPWR hold476/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_8
X_4055_ _4076_/B _7071_/Q _3856_/A _4054_/X VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_45_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7432_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4155__S _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4382__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4957_ _4953_/X _4956_/Y _4955_/X VGND VGND VPWR VPWR _4958_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3908_ _7230_/Q _3617_/X _3682_/X _7225_/Q _3907_/X VGND VGND VPWR VPWR _3913_/B
+ sky130_fd_sc_hd__a221o_4
XANTENNA__3775__A2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4972__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout517_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4888_ _4856_/A _4888_/B _5282_/A _5058_/D VGND VGND VPWR VPWR _4888_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_0_74_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6627_ _7358_/Q _6459_/B _6459_/C _6408_/B _7382_/Q VGND VGND VPWR VPWR _6627_/X
+ sky130_fd_sc_hd__a32o_1
X_3839_ _7043_/Q _4370_/A _3673_/X _7199_/Q VGND VGND VPWR VPWR _3839_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_62_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5516__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_171_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5921__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6558_ _7443_/Q _6424_/C _6771_/A3 _6466_/X _7507_/Q VGND VGND VPWR VPWR _6558_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5509_ _4726_/Y _4796_/Y _4844_/Y _4930_/B _5237_/C VGND VGND VPWR VPWR _5510_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6489_ _7552_/Q _6408_/A _6408_/D _7536_/Q _6488_/X VGND VGND VPWR VPWR _6494_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6477__A1 _7512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6477__B2 _7504_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4488__A0 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4838__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7187__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6229__A1 _7524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6244__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4573__B _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A2 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3766__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4963__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6165__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6704__A2 _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7512__SET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6180__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3933__A _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4748__B _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__B _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5140__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5979__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6640__B2 _7470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3454__A1 _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5860_ _5896_/A0 _5860_/A1 _5865_/S VGND VGND VPWR VPWR _5860_/X sky130_fd_sc_hd__mux2_1
X_4811_ _4811_/A _5138_/A _5138_/B _5113_/A VGND VGND VPWR VPWR _4812_/C sky130_fd_sc_hd__nand4_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5791_ _5791_/A0 _5953_/A1 _5793_/S VGND VGND VPWR VPWR _5791_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7530_ _7530_/CLK _7530_/D fanout600/X VGND VGND VPWR VPWR _7530_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3757__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4742_ _4888_/B _5282_/A VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__nand2b_4
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7461_ _7478_/CLK _7461_/D fanout585/X VGND VGND VPWR VPWR _7461_/Q sky130_fd_sc_hd__dfrtp_4
X_4673_ _5071_/A _4675_/B _4675_/C VGND VGND VPWR VPWR _4673_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__6156__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6412_ _6463_/A _6747_/C _6651_/B VGND VGND VPWR VPWR _6420_/A sky130_fd_sc_hd__and3_4
XFILLER_0_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5903__A0 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3624_ _7300_/Q hold12/A _4346_/C _5776_/A _7388_/Q VGND VGND VPWR VPWR _3624_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3509__A2 _3564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7392_ _7566_/CLK _7392_/D fanout599/X VGND VGND VPWR VPWR _7392_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6171__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6343_ _7018_/Q _6121_/C _6086_/X _6342_/X VGND VGND VPWR VPWR _6343_/X sky130_fd_sc_hd__a31o_1
X_3555_ _5785_/A _4551_/A hold22/A VGND VGND VPWR VPWR _5776_/A sky130_fd_sc_hd__and3_4
Xhold3104 _7209_/Q VGND VGND VPWR VPWR hold3104/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6274_ _7518_/Q _6094_/A _6317_/C _6085_/X _7502_/Q VGND VGND VPWR VPWR _6274_/X
+ sky130_fd_sc_hd__a32o_1
X_3486_ _5590_/A _4449_/B _5612_/B VGND VGND VPWR VPWR _3486_/X sky130_fd_sc_hd__and3_4
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3115 _4266_/X VGND VGND VPWR VPWR hold3115/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3126 hold3126/A VGND VGND VPWR VPWR _5588_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_110_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3562__B _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3137 hold3137/A VGND VGND VPWR VPWR _4395_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5225_ _4933_/B _5213_/C _5342_/B _5102_/B _5357_/B2 VGND VGND VPWR VPWR _5228_/C
+ sky130_fd_sc_hd__a32oi_2
XANTENNA__5131__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2403 _6965_/Q VGND VGND VPWR VPWR hold999/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3148 _7559_/Q VGND VGND VPWR VPWR hold3148/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3159 _5613_/X VGND VGND VPWR VPWR _7243_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2414 _7149_/Q VGND VGND VPWR VPWR hold957/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2425 hold718/X VGND VGND VPWR VPWR _5675_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2436 _7154_/Q VGND VGND VPWR VPWR hold987/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1702 _7529_/Q VGND VGND VPWR VPWR hold312/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2447 hold933/X VGND VGND VPWR VPWR _5788_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5156_ _5156_/A _5156_/B _5156_/C VGND VGND VPWR VPWR _5160_/B sky130_fd_sc_hd__nand3_1
Xhold2458 hold973/X VGND VGND VPWR VPWR _4307_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1713 _5627_/X VGND VGND VPWR VPWR hold337/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1724 hold42/X VGND VGND VPWR VPWR hold1724/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2469 _7288_/Q VGND VGND VPWR VPWR hold631/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3693__A1 _7347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1735 _5945_/X VGND VGND VPWR VPWR hold119/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4107_ _4107_/A _4117_/B VGND VGND VPWR VPWR _4107_/Y sky130_fd_sc_hd__nor2_1
Xhold1746 _5778_/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1757 _5873_/X VGND VGND VPWR VPWR hold113/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5087_ _4717_/Y _4960_/A _5086_/Y _5085_/Y VGND VGND VPWR VPWR _5087_/Y sky130_fd_sc_hd__o211ai_1
Xhold1768 _7062_/Q VGND VGND VPWR VPWR hold1768/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1779 _5987_/X VGND VGND VPWR VPWR hold387/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4038_ _4037_/Y _4029_/X _4025_/A _6901_/Q VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_154_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6395__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A0 _5998_/A1 _5991_/S VGND VGND VPWR VPWR _5989_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_176_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3748__A2 _3506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3737__B _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_50 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7659_ _7659_/A VGND VGND VPWR VPWR _7659_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_61 _6212_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_72 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4849__A _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3920__A2 _5929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input167_A wb_sel_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput190 _3422_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_0_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3684__A1 _7283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3684__B2 _7451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2970 _6963_/Q VGND VGND VPWR VPWR hold2970/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input28_A mask_rev_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2981 _7163_/Q VGND VGND VPWR VPWR hold2981/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2992 hold2992/A VGND VGND VPWR VPWR _5742_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_leaf_67_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5399__B _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3987__A2 _3543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5189__A1 _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6386__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3928__A _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3739__A2 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4750__C _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3647__B _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6689__A1 _7198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6153__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold309 hold309/A VGND VGND VPWR VPWR _7561_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4759__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3663__A _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3911__A2 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4909__D _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_12__f_wb_clk_i clkbuf_3_6_0_wb_clk_i/X VGND VGND VPWR VPWR _7207_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_175_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _4996_/A _5339_/C _5553_/A1 VGND VGND VPWR VPWR _5011_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1009 _4433_/X VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_30_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6961_ _7024_/CLK _6961_/D fanout566/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_108_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5102__B _5102_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5912_ _5912_/A0 hold464/X _5919_/S VGND VGND VPWR VPWR _5912_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3978__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6892_ _4127_/A1 _6892_/D _6842_/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5843_ _5843_/A0 _5996_/A1 _5847_/S VGND VGND VPWR VPWR _5843_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6377__B1 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_192_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5774_ _5774_/A0 _5999_/A1 _5775_/S VGND VGND VPWR VPWR _5774_/X sky130_fd_sc_hd__mux2_1
X_7513_ _7513_/CLK _7513_/D fanout602/X VGND VGND VPWR VPWR _7513_/Q sky130_fd_sc_hd__dfrtp_4
X_4725_ _5222_/B _4726_/B _4726_/C _5005_/A VGND VGND VPWR VPWR _4725_/X sky130_fd_sc_hd__and4_1
XFILLER_0_90_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6129__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2933_A _7027_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4656_ _4667_/A _4608_/Y _4657_/C _4657_/B VGND VGND VPWR VPWR _4889_/A sky130_fd_sc_hd__o211ai_4
X_7444_ _7565_/CLK _7444_/D fanout599/X VGND VGND VPWR VPWR _7444_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3607_ _3575_/X _3607_/B _3607_/C VGND VGND VPWR VPWR _3607_/Y sky130_fd_sc_hd__nand3b_4
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _4176_/B sky130_fd_sc_hd__buf_4
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_2
Xhold810 hold810/A VGND VGND VPWR VPWR _7421_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4587_ _5071_/A _4593_/A _4687_/B VGND VGND VPWR VPWR _4755_/A sky130_fd_sc_hd__a21boi_4
Xhold821 hold821/A VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7375_ _7471_/CLK _7375_/D fanout593/X VGND VGND VPWR VPWR _7375_/Q sky130_fd_sc_hd__dfstp_2
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR _4140_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold832 _5954_/X VGND VGND VPWR VPWR _7541_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap551 _5387_/B VGND VGND VPWR VPWR _5399_/B sky130_fd_sc_hd__buf_12
Xhold843 hold843/A VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold854 hold854/A VGND VGND VPWR VPWR hold854/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6326_ _7052_/Q _6087_/X _6120_/X _7017_/Q _6325_/X VGND VGND VPWR VPWR _6327_/D
+ sky130_fd_sc_hd__a221o_1
X_3538_ _4551_/A _3569_/A _5938_/C VGND VGND VPWR VPWR _5929_/A sky130_fd_sc_hd__and3_4
Xhold865 _5702_/X VGND VGND VPWR VPWR _7317_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4388__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold876 hold876/A VGND VGND VPWR VPWR hold876/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold887 hold887/A VGND VGND VPWR VPWR hold887/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold898 _5755_/X VGND VGND VPWR VPWR _7364_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5104__A1 _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6257_ _6257_/A _6257_/B _6257_/C _6257_/D VGND VGND VPWR VPWR _6257_/Y sky130_fd_sc_hd__nor4_1
XANTENNA__6301__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3469_ _6901_/Q _6900_/Q _4025_/A VGND VGND VPWR VPWR _3469_/X sky130_fd_sc_hd__mux2_1
Xhold2200 _7494_/Q VGND VGND VPWR VPWR hold492/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2211 _7470_/Q VGND VGND VPWR VPWR hold543/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2222 _6907_/Q VGND VGND VPWR VPWR _3450_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_5208_ _5451_/A1 _4796_/Y _4946_/Y _4930_/C VGND VGND VPWR VPWR _5208_/Y sky130_fd_sc_hd__o31ai_1
Xhold2233 _5865_/X VGND VGND VPWR VPWR hold503/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2244 _7296_/Q VGND VGND VPWR VPWR hold536/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6188_ _7442_/Q _6097_/X _6121_/X _7306_/Q _6187_/X VGND VGND VPWR VPWR _6188_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2255 hold604/X VGND VGND VPWR VPWR _5697_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1510 hold25/X VGND VGND VPWR VPWR _5937_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1521 _4443_/X VGND VGND VPWR VPWR hold218/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2266 _7486_/Q VGND VGND VPWR VPWR hold555/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5139_ _5013_/X _5139_/B _5139_/C _5139_/D VGND VGND VPWR VPWR _5139_/X sky130_fd_sc_hd__and4b_1
Xhold2277 hold516/X VGND VGND VPWR VPWR _5991_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1532 hold212/X VGND VGND VPWR VPWR _7532_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1543 _5924_/X VGND VGND VPWR VPWR hold230/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2288 _7422_/Q VGND VGND VPWR VPWR hold600/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2299 hold901/X VGND VGND VPWR VPWR _5710_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1554 _5917_/X VGND VGND VPWR VPWR hold206/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1565 _5935_/X VGND VGND VPWR VPWR hold216/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1576 hold268/X VGND VGND VPWR VPWR _7353_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5407__A2 _4945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1587 _4391_/X VGND VGND VPWR VPWR hold357/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1598 _5698_/X VGND VGND VPWR VPWR hold266/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_168_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5012__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1699_A _7517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3969__A2 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5947__B _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6368__B1 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4570__C _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5591__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4579__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6540__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold3247_A _6898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4854__B1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3930__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5203__A _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output301_A _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5857__B hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6359__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3658__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4510_ _4510_/A0 _5714_/A0 _4514_/S VGND VGND VPWR VPWR _4510_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3593__B1 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5490_ _5158_/A _4952_/B _5052_/B _5489_/X VGND VGND VPWR VPWR _5532_/B sky130_fd_sc_hd__a211oi_2
XFILLER_0_81_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4441_ _4441_/A0 hold464/X _4448_/S VGND VGND VPWR VPWR _4441_/X sky130_fd_sc_hd__mux2_1
Xhold106 hold106/A VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold117 _5936_/X VGND VGND VPWR VPWR _7525_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold128 hold128/A VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold139 hold139/A VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7160_ _7190_/CLK _7160_/D _6871_/A VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4372_ _5940_/A1 _4372_/A1 _4375_/S VGND VGND VPWR VPWR _4372_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_186_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6112_/C _6106_/B _6121_/A _6119_/A VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__and4bb_4
Xfanout608 input164/X VGND VGND VPWR VPWR _6780_/B sky130_fd_sc_hd__buf_12
XANTENNA_hold36_A hold36/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7091_ _7530_/CLK hold79/X fanout605/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 _4743_/A VGND VGND VPWR VPWR _5058_/D sky130_fd_sc_hd__buf_12
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6295__C1 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6042_ _7594_/Q _7593_/Q VGND VGND VPWR VPWR _6434_/B sky130_fd_sc_hd__and2_4
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5113__A _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6598__B1 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6944_ _7278_/CLK _6944_/D fanout580/X VGND VGND VPWR VPWR _7650_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4952__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5767__B _5911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3820__A1 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6875_ _7156_/CLK _6875_/D _6833_/A VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5826_ _5826_/A0 _5997_/A1 _5829_/S VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6365__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5757_ _5757_/A0 _5955_/A1 _5757_/S VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6770__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4708_ _4888_/B _5282_/A _5399_/B VGND VGND VPWR VPWR _5113_/A sky130_fd_sc_hd__and3_4
X_5688_ _5967_/A1 _5688_/A1 _5694_/S VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6117__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7427_ _7471_/CLK _7427_/D fanout593/X VGND VGND VPWR VPWR _7427_/Q sky130_fd_sc_hd__dfrtp_2
X_4639_ _4667_/A _5301_/A1 _4636_/Y VGND VGND VPWR VPWR _4641_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 _5988_/X VGND VGND VPWR VPWR _7571_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7358_ _7555_/CLK _7358_/D fanout594/X VGND VGND VPWR VPWR _7358_/Q sky130_fd_sc_hd__dfrtp_4
Xhold651 hold651/A VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold662 hold662/A VGND VGND VPWR VPWR hold662/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6110__C _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold673 _5805_/X VGND VGND VPWR VPWR _7408_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5007__B _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold684 hold684/A VGND VGND VPWR VPWR hold684/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6309_ _7012_/Q _6136_/B _6120_/B _6110_/A VGND VGND VPWR VPWR _6309_/X sky130_fd_sc_hd__a31o_1
Xhold695 _4487_/X VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmgmt_gpio_30_buff_inst _4164_/X VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__clkbuf_8
X_7289_ _7359_/CLK _7289_/D fanout575/X VGND VGND VPWR VPWR _7289_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6825__A1 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2030 _7200_/Q VGND VGND VPWR VPWR hold442/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3639__B2 _7673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2041 _5786_/X VGND VGND VPWR VPWR _7391_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2052 hold384/X VGND VGND VPWR VPWR _4404_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2063 hold682/X VGND VGND VPWR VPWR _4239_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7416__SET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6119__A _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2074 hold97/X VGND VGND VPWR VPWR _7491_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2085 hold94/X VGND VGND VPWR VPWR _4436_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1340 _4319_/A1 VGND VGND VPWR VPWR hold2806/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6038__C1 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2096 _6878_/Q VGND VGND VPWR VPWR hold143/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1351 _4300_/A1 VGND VGND VPWR VPWR hold2848/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1362 _6790_/A1 VGND VGND VPWR VPWR hold2914/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_169_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1373 hold1905/X VGND VGND VPWR VPWR hold1906/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1384 hold1699/X VGND VGND VPWR VPWR hold1700/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6589__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1395 hold1395/A VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1983_A _7185_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__B1 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5677__B _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4581__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3811__A1 _7289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3478__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6356__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input95_A usr1_vcc_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6761__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3575__B1 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3925__B _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5316__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6513__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3878__A1 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3660__B _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6292__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4248__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4055__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4990_ _5183_/A _5295_/C _5038_/B _5203_/B VGND VGND VPWR VPWR _5037_/C sky130_fd_sc_hd__nand4_1
XANTENNA__5587__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3941_ _7551_/Q _3508_/X _4422_/S input43/X _3940_/X VGND VGND VPWR VPWR _3941_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4491__B _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6660_ _7112_/Q _6651_/B _6426_/X _6659_/X VGND VGND VPWR VPWR _6660_/X sky130_fd_sc_hd__a31o_1
X_3872_ _7568_/Q _5983_/A _5992_/C _3869_/X _3871_/X VGND VGND VPWR VPWR _3872_/X
+ sky130_fd_sc_hd__a311o_2
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5611_ _5611_/A0 _5955_/A1 _5611_/S VGND VGND VPWR VPWR _5611_/X sky130_fd_sc_hd__mux2_1
X_6591_ _7452_/Q _6443_/X _6446_/X _7524_/Q _6574_/X VGND VGND VPWR VPWR _6591_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5807__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5542_ _4622_/Y _4726_/Y _4748_/Y _5512_/A _5462_/X VGND VGND VPWR VPWR _5543_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_121_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6504__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5473_ _4791_/A _5473_/B _5473_/C _5473_/D VGND VGND VPWR VPWR _5518_/A sky130_fd_sc_hd__and4b_1
XANTENNA__3581__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7212_ _7212_/CLK _7212_/D fanout574/X VGND VGND VPWR VPWR _7212_/Q sky130_fd_sc_hd__dfrtp_4
X_4424_ _7102_/Q _6827_/A VGND VGND VPWR VPWR _4424_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7143_ _7266_/CLK _7143_/D fanout567/X VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfrtp_4
X_4355_ _4355_/A0 _5914_/A1 _4357_/S VGND VGND VPWR VPWR _4355_/X sky130_fd_sc_hd__mux2_1
Xfanout416 _3480_/X VGND VGND VPWR VPWR _5938_/B sky130_fd_sc_hd__buf_12
XANTENNA__6268__C1 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7074_ _7075_/CLK _7074_/D _6864_/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout438 _6078_/X VGND VGND VPWR VPWR _6116_/A sky130_fd_sc_hd__buf_8
X_4286_ _4289_/S _6789_/A2 _4285_/Y VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__4666__B _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6025_ _6144_/A _6136_/B _6051_/C VGND VGND VPWR VPWR _6025_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4719__A_N _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _7363_/CLK _6927_/D fanout575/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_162_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6858_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6858_/X sky130_fd_sc_hd__and2_1
XANTENNA__6338__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5809_ _5809_/A0 _5953_/A1 _5811_/S VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6743__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6789_ _6789_/A1 _6789_/A2 _6788_/Y VGND VGND VPWR VPWR _7633_/D sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6121__B _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6510__A3 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold470 _7013_/Q VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold481 hold481/A VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold492 hold492/A VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 hold1170/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
XFILLER_0_169_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input10_A mask_rev_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1181 hold2914/X VGND VGND VPWR VPWR hold1181/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1192 hold1192/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
XFILLER_0_87_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__B1 _5102_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6577__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6734__B1 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3655__B hold36/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6031__B _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3671__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4140_ _4142_/A _4140_/B VGND VGND VPWR VPWR _4140_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__6265__A2 _6073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4071_ hold1/A hold82/A _4075_/S VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4276__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4933__C _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5225__B1 _5102_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4973_ _4709_/Y _4748_/Y _4814_/Y _4826_/Y VGND VGND VPWR VPWR _5200_/C sky130_fd_sc_hd__a211o_2
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_176_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3787__B1 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6712_ _7169_/Q _6408_/D _6427_/X _7119_/Q _6711_/X VGND VGND VPWR VPWR _6712_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_19_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3924_ _3923_/X _3924_/A1 _3996_/A VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3549__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6643_ _7550_/Q _6419_/A _6467_/X _7422_/Q _6642_/X VGND VGND VPWR VPWR _6643_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6725__B1 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3855_ _3855_/A _3855_/B _3855_/C VGND VGND VPWR VPWR _3856_/B sky130_fd_sc_hd__and3_4
XFILLER_0_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3539__B1 _5929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4441__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4200__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3786_ _7165_/Q _3663_/X _3666_/X _7014_/Q _3785_/X VGND VGND VPWR VPWR _3792_/C
+ sky130_fd_sc_hd__a221o_1
X_6574_ _7444_/Q _6574_/B _6574_/C VGND VGND VPWR VPWR _6574_/X sky130_fd_sc_hd__and3_1
XFILLER_0_6_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6740__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3565__B _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5525_ _4817_/X _5453_/C _5395_/X _5521_/Y _5524_/X VGND VGND VPWR VPWR _5525_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4751__A2 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5456_ _5545_/C _5541_/D _5456_/C _5543_/A VGND VGND VPWR VPWR _5457_/A sky130_fd_sc_hd__and4b_1
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4407_ _4422_/S _4215_/X _4406_/Y _5992_/D VGND VGND VPWR VPWR _4423_/S sky130_fd_sc_hd__o211a_4
XANTENNA__5700__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5387_ _4887_/B _5387_/B _5387_/C _5387_/D VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__and4b_1
XANTENNA_fanout497_A hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7126_ _7134_/CLK _7126_/D _6833_/A VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfrtp_4
X_4338_ _4338_/A0 _5852_/A0 _4339_/S VGND VGND VPWR VPWR _4338_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input2_A debug_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6256__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4269_ _4269_/A0 _5647_/A0 _4270_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
X_7057_ _7070_/CLK _7057_/D fanout590/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4267__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6008_ _6005_/Y _6006_/X _6018_/A VGND VGND VPWR VPWR _7584_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_179_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6116__B _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6716__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input58_A mgmt_gpio_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6247__A2 _6116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4258__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5910__S _5910_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5470__A3 _4971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_0__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3410__1 _7075_/CLK VGND VGND VPWR VPWR _6881_/CLK sky130_fd_sc_hd__inv_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6707__B1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3784__A3 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3666__A hold36/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3640_ _7396_/Q _5803_/A _3933_/A _3564_/X _7364_/Q VGND VGND VPWR VPWR _3640_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3571_ _6893_/Q _7073_/Q VGND VGND VPWR VPWR _3996_/A sky130_fd_sc_hd__nand2_8
XANTENNA__3536__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3941__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5310_ _4583_/B _4783_/Y _4789_/Y _4744_/Y _5153_/B VGND VGND VPWR VPWR _5488_/A
+ sky130_fd_sc_hd__o221a_1
X_6290_ _7187_/Q _6119_/A _6106_/B _6136_/B _6121_/C VGND VGND VPWR VPWR _6290_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5241_ _4935_/X _5243_/C _5239_/X VGND VGND VPWR VPWR _5244_/C sky130_fd_sc_hd__a21o_1
XANTENNA__5694__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2607 _5828_/X VGND VGND VPWR VPWR hold851/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5172_ _4877_/A _5180_/B _5018_/B _5180_/A VGND VGND VPWR VPWR _5172_/X sky130_fd_sc_hd__a22o_1
Xhold2618 hold870/X VGND VGND VPWR VPWR _5882_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2629 _4255_/X VGND VGND VPWR VPWR hold648/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6238__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4123_ _6890_/Q _4123_/B _4123_/C VGND VGND VPWR VPWR _4123_/Y sky130_fd_sc_hd__nand3_1
Xhold1906 hold1906/A VGND VGND VPWR VPWR _5963_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5105__B _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1917 _6955_/Q VGND VGND VPWR VPWR hold124/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1928 _5879_/X VGND VGND VPWR VPWR hold401/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5820__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1939 hold360/X VGND VGND VPWR VPWR _5798_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4054_ _6910_/Q _6909_/Q _6908_/Q _4062_/A _4054_/B1 VGND VGND VPWR VPWR _4054_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_127_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5997__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4382__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4956_ _4956_/A _4956_/B VGND VGND VPWR VPWR _4956_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_191_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_163_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3907_ _7408_/Q _5803_/A _5947_/A _4485_/A _7143_/Q VGND VGND VPWR VPWR _3907_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4972__A2 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4887_ _4747_/B _4887_/B _4945_/A _4887_/D VGND VGND VPWR VPWR _4940_/C sky130_fd_sc_hd__and4b_4
XFILLER_0_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3576__A _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6626_ _7534_/Q _6058_/X _6409_/X _7406_/Q VGND VGND VPWR VPWR _6626_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6174__A1 _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3838_ _7377_/Q _4473_/A _5983_/A _3658_/X _7114_/Q VGND VGND VPWR VPWR _3838_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6713__A3 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6557_ _7563_/Q _6419_/C _6434_/X _7467_/Q _6556_/X VGND VGND VPWR VPWR _6557_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3769_ input29/X _3503_/X _3520_/X _7442_/Q _3768_/X VGND VGND VPWR VPWR _3769_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5508_ _5508_/A _5508_/B _5508_/C VGND VGND VPWR VPWR _5575_/A sky130_fd_sc_hd__and3_2
XANTENNA__3932__B1 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6488_ _7472_/Q _6574_/B _6441_/X _6423_/X _7328_/Q VGND VGND VPWR VPWR _6488_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6477__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5439_ _5107_/A _5342_/A _5180_/B _5260_/D _5058_/C VGND VGND VPWR VPWR _5439_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4838__C _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _7207_/CLK _7109_/D _4309_/B VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5730__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f_user_clock clkbuf_0_user_clock/X VGND VGND VPWR VPWR _4163_/A1 sky130_fd_sc_hd__clkbuf_16
XANTENNA__5988__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_187_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4573__C _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input112_A wb_adr_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4412__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3766__A3 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3486__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5912__A1 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_csclk_A _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5905__S _5910_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11__f_wb_clk_i clkbuf_3_5_0_wb_clk_i/X VGND VGND VPWR VPWR _7630_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6640__A2 _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4810_ _5138_/A _5138_/B _4810_/C _5453_/B VGND VGND VPWR VPWR _4812_/B sky130_fd_sc_hd__nand4_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4403__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5790_ _5790_/A0 _5979_/A0 _5793_/S VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4741_ _5074_/B _4814_/C VGND VGND VPWR VPWR _4741_/Y sky130_fd_sc_hd__nand2_8
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7460_ _7581_/CLK _7460_/D fanout584/X VGND VGND VPWR VPWR _7460_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4672_ _4861_/A _4861_/B _4667_/Y _4669_/X VGND VGND VPWR VPWR _4672_/X sky130_fd_sc_hd__a211o_4
XFILLER_0_98_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6411_ _6467_/A _6651_/B _6409_/X _6410_/X _6600_/B VGND VGND VPWR VPWR _6411_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_3623_ _3623_/A _3623_/B _3623_/C _3623_/D VGND VGND VPWR VPWR _3643_/A sky130_fd_sc_hd__nor4_2
XANTENNA__3509__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7391_ _7487_/CLK _7391_/D fanout593/X VGND VGND VPWR VPWR _7391_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_153_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5815__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3914__B1 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6342_ _7058_/Q _6332_/B _6084_/X _6121_/X _6990_/Q VGND VGND VPWR VPWR _6342_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3554_ _4176_/B _4248_/S _4231_/S input42/X _3551_/X VGND VGND VPWR VPWR _3568_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3485_ hold280/X _3485_/B _3511_/A VGND VGND VPWR VPWR _3485_/X sky130_fd_sc_hd__and3b_4
X_6273_ _7462_/Q _6080_/X _6269_/X _6270_/X _6272_/X VGND VGND VPWR VPWR _6280_/A
+ sky130_fd_sc_hd__a2111o_1
Xhold3105 hold3105/A VGND VGND VPWR VPWR _5582_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3116 _7431_/Q VGND VGND VPWR VPWR hold3116/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3127 _5588_/X VGND VGND VPWR VPWR hold3127/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5224_ _5224_/A _5349_/A _5224_/C VGND VGND VPWR VPWR _5228_/B sky130_fd_sc_hd__nor3_1
Xhold3138 _4395_/X VGND VGND VPWR VPWR hold3138/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3562__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2404 hold999/X VGND VGND VPWR VPWR _4269_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5131__A2 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3149 hold3149/A VGND VGND VPWR VPWR _5975_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2415 hold957/X VGND VGND VPWR VPWR _4494_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2426 _7266_/Q VGND VGND VPWR VPWR hold684/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2437 hold987/X VGND VGND VPWR VPWR _4500_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2448 _7128_/Q VGND VGND VPWR VPWR hold653/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5155_ _4956_/A _4690_/Y _4802_/Y _4796_/Y _4706_/Y VGND VGND VPWR VPWR _5156_/C
+ sky130_fd_sc_hd__o32a_1
Xhold1703 hold312/X VGND VGND VPWR VPWR _5941_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1714 hold337/X VGND VGND VPWR VPWR _7253_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2459 _6928_/Q VGND VGND VPWR VPWR hold656/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3693__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1725 hold1725/A VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4106_ _7585_/Q _7584_/Q _7586_/Q _7587_/Q VGND VGND VPWR VPWR _4107_/A sky130_fd_sc_hd__nand4bb_4
XFILLER_0_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1736 _7053_/Q VGND VGND VPWR VPWR hold408/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5086_ _5094_/A _5086_/B VGND VGND VPWR VPWR _5086_/Y sky130_fd_sc_hd__nand2_1
Xhold1747 _7562_/Q VGND VGND VPWR VPWR hold296/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1758 _7576_/Q VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1769 hold1769/A VGND VGND VPWR VPWR _4396_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4166__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4037_ _6901_/Q _6900_/Q _6902_/Q VGND VGND VPWR VPWR _4037_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6631__A2 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _5988_/A0 _5997_/A1 _5991_/S VGND VGND VPWR VPWR _5988_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4939_ _4954_/A _5453_/A _5183_/C _4940_/D VGND VGND VPWR VPWR _4941_/A sky130_fd_sc_hd__and4_1
XFILLER_0_136_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4840__D _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_40 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3737__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7658_ _7658_/A VGND VGND VPWR VPWR _7658_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_191_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_51 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _7174_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_73 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _7301_/Q _6420_/A _6421_/X _7325_/Q _6608_/X VGND VGND VPWR VPWR _6609_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7589_ _7593_/CLK _7589_/D fanout567/X VGND VGND VPWR VPWR _7589_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5725__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6162__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5370__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5658__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput180 _3431_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput191 _3421_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_0_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3684__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2960 _7504_/Q VGND VGND VPWR VPWR hold2960/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold3025_A _7233_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2971 hold2971/A VGND VGND VPWR VPWR _4267_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2982 hold2982/A VGND VGND VPWR VPWR _4511_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2993 _7173_/Q VGND VGND VPWR VPWR hold2993/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6083__B1 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6622__A2 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5399__C _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5291__D1 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5189__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6386__A1 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6386__B2 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5043__D1 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4397__A0 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3739__A3 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4105__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3647__C hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6689__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5897__A0 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7569_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3663__B _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3911__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5649__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__B2 _7123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4321__A0 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7359_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4775__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7078__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4609__D1 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6613__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6960_ _7024_/CLK _6960_/D fanout567/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfstp_2
X_5911_ _5911_/A _5938_/C _5992_/D VGND VGND VPWR VPWR _5919_/S sky130_fd_sc_hd__and3_4
XFILLER_0_76_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6891_ _7075_/CLK _6891_/D _6841_/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3978__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5842_ _5842_/A0 _5914_/A1 _5847_/S VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5773_ _5773_/A0 _5953_/A1 _5775_/S VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__mux2_1
X_7512_ _7513_/CLK _7512_/D fanout602/X VGND VGND VPWR VPWR _7512_/Q sky130_fd_sc_hd__dfstp_4
X_4724_ _4088_/Y _4558_/X _4647_/Y VGND VGND VPWR VPWR _4948_/C sky130_fd_sc_hd__o21a_4
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6129__A1 _7448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7443_ _7505_/CLK _7443_/D fanout601/X VGND VGND VPWR VPWR _7443_/Q sky130_fd_sc_hd__dfrtp_4
X_4655_ _4667_/A _4571_/Y _5387_/B _4657_/C _4657_/B VGND VGND VPWR VPWR _5213_/A
+ sky130_fd_sc_hd__o311a_4
XFILLER_0_32_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_2
X_3606_ _3606_/A _3606_/B _3606_/C _3606_/D VGND VGND VPWR VPWR _3607_/C sky130_fd_sc_hd__nor4_2
Xhold800 hold800/A VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7374_ _7582_/CLK _7374_/D fanout584/X VGND VGND VPWR VPWR _7374_/Q sky130_fd_sc_hd__dfrtp_4
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__buf_2
Xhold811 hold811/A VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4586_ _4675_/A _4675_/B _4586_/C _5089_/B VGND VGND VPWR VPWR _4687_/B sky130_fd_sc_hd__nand4_4
Xinput82 spi_sdoenb VGND VGND VPWR VPWR _4144_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap530 _4888_/Y VGND VGND VPWR VPWR _5528_/A3 sky130_fd_sc_hd__buf_8
Xhold822 _5720_/X VGND VGND VPWR VPWR _7333_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_6
Xmax_cap541 _4715_/Y VGND VGND VPWR VPWR _5357_/B2 sky130_fd_sc_hd__clkbuf_2
Xhold833 hold833/A VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6325_ _7198_/Q _6110_/A _6079_/X _6099_/X _7027_/Q VGND VGND VPWR VPWR _6325_/X
+ sky130_fd_sc_hd__a32o_1
Xhold844 _4339_/X VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold855 _5747_/X VGND VGND VPWR VPWR _7357_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3537_ _3537_/A _4509_/A _4491_/C VGND VGND VPWR VPWR _3537_/X sky130_fd_sc_hd__and3_4
Xhold866 hold866/A VGND VGND VPWR VPWR hold866/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3902__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4388__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold877 hold877/A VGND VGND VPWR VPWR _7341_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold888 hold888/A VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold899 hold899/A VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6256_ _7533_/Q _6092_/X _6252_/X _6253_/X _6255_/X VGND VGND VPWR VPWR _6257_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_149_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6301__B2 _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3468_ _3468_/A1 _3468_/A2 hold154/X _3465_/Y VGND VGND VPWR VPWR _3468_/X sky130_fd_sc_hd__a22o_1
Xhold2201 hold492/X VGND VGND VPWR VPWR _5901_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4312__A0 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2212 hold543/X VGND VGND VPWR VPWR _5874_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2223 _3451_/Y VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5207_ _4956_/A _4709_/Y _4659_/Y VGND VGND VPWR VPWR _5419_/A sky130_fd_sc_hd__a21o_1
Xhold2234 _7536_/Q VGND VGND VPWR VPWR hold540/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6187_ _7490_/Q _6094_/A _6093_/X _6100_/X _7474_/Q VGND VGND VPWR VPWR _6187_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1500 hold173/X VGND VGND VPWR VPWR _5845_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2245 hold536/X VGND VGND VPWR VPWR _5679_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout577_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3399_ _6900_/Q VGND VGND VPWR VPWR _3399_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4863__A1 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2256 _7328_/Q VGND VGND VPWR VPWR hold532/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1511 _5937_/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1522 _7281_/Q VGND VGND VPWR VPWR hold203/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2267 hold555/X VGND VGND VPWR VPWR _5892_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1533 _7438_/Q VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2278 _7454_/Q VGND VGND VPWR VPWR hold557/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5138_ _5138_/A _5138_/B _5138_/C _5138_/D VGND VGND VPWR VPWR _5138_/Y sky130_fd_sc_hd__nand4_1
Xhold1544 hold230/X VGND VGND VPWR VPWR _7514_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_leaf_11_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2289 hold600/X VGND VGND VPWR VPWR _5820_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1555 hold206/X VGND VGND VPWR VPWR _7508_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1566 _7452_/Q VGND VGND VPWR VPWR hold219/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5407__A3 _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1577 _7582_/Q VGND VGND VPWR VPWR hold1577/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5069_ _5091_/A _5072_/B _5260_/C VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__and3_4
XFILLER_0_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1588 hold357/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1599 _7385_/Q VGND VGND VPWR VPWR hold263/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_79_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3969__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5947__C hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6368__B2 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1761_A _7546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4579__B _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6540__A1 _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input40_A mgmt_gpio_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4595__A _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3930__C _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2790 hold2790/A VGND VGND VPWR VPWR hold2790/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6359__A1 _7155_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3658__B _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3674__A _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4440_ _7257_/Q hold284/X _4168_/D _4422_/S _5992_/D VGND VGND VPWR VPWR _4448_/S
+ sky130_fd_sc_hd__o311a_4
Xhold107 hold107/A VGND VGND VPWR VPWR _7339_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6531__B2 _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold118 hold118/A VGND VGND VPWR VPWR hold118/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold129 _5682_/X VGND VGND VPWR VPWR _7299_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4371_ _5840_/A1 _4371_/A1 _4375_/S VGND VGND VPWR VPWR _4371_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3896__A2 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6110_ _6110_/A _6121_/A _6144_/B VGND VGND VPWR VPWR _6110_/X sky130_fd_sc_hd__and3_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 _4860_/A VGND VGND VPWR VPWR _4740_/D sky130_fd_sc_hd__buf_12
X_7090_ _7530_/CLK _7090_/D fanout605/X VGND VGND VPWR VPWR _7669_/A sky130_fd_sc_hd__dfrtp_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6295__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6041_ _7593_/Q _6051_/C _6040_/Y VGND VGND VPWR VPWR _7593_/D sky130_fd_sc_hd__a21oi_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6943_ _7278_/CLK _6943_/D fanout580/X VGND VGND VPWR VPWR _7649_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4444__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5270__B2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6874_ _7201_/CLK _6874_/D _6833_/A VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3820__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5825_ _5825_/A0 _5987_/A1 _5829_/S VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5756_ _5756_/A0 _5954_/A1 _5757_/S VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6770__B2 _7201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4707_ _5091_/C _5260_/C VGND VGND VPWR VPWR _4707_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__3584__B2 _7469_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5687_ _5903_/A0 _5687_/A1 _5694_/S VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7426_ _7556_/CLK _7426_/D fanout594/X VGND VGND VPWR VPWR _7426_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4638_ _4667_/A _5301_/A1 _4636_/Y VGND VGND VPWR VPWR _4801_/C sky130_fd_sc_hd__o21a_4
XFILLER_0_13_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold630 _4366_/X VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7357_ _7429_/CLK _7357_/D fanout583/X VGND VGND VPWR VPWR _7357_/Q sky130_fd_sc_hd__dfrtp_4
X_4569_ _4795_/C _4984_/B _4805_/B VGND VGND VPWR VPWR _4615_/A sky130_fd_sc_hd__and3_2
Xhold641 hold641/A VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold652 _5997_/X VGND VGND VPWR VPWR _7579_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold663 _4305_/X VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold674 hold674/A VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6308_ _7002_/Q _6097_/B _6120_/B _6332_/C _7032_/Q VGND VGND VPWR VPWR _6308_/X
+ sky130_fd_sc_hd__a32o_1
Xhold685 _5645_/X VGND VGND VPWR VPWR _7266_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7288_ _7363_/CLK _7288_/D fanout575/X VGND VGND VPWR VPWR _7288_/Q sky130_fd_sc_hd__dfstp_4
Xhold696 hold696/A VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6286__B1 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6239_ _7373_/Q _6084_/X _6093_/X _7365_/Q VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__a22o_1
Xhold2020 _4374_/X VGND VGND VPWR VPWR hold439/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2031 hold442/X VGND VGND VPWR VPWR _4555_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3639__A2 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2042 _7252_/Q VGND VGND VPWR VPWR hold578/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2053 _7322_/Q VGND VGND VPWR VPWR hold565/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2064 _4239_/X VGND VGND VPWR VPWR hold683/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1330 _5804_/X VGND VGND VPWR VPWR _7407_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2075 _7531_/Q VGND VGND VPWR VPWR hold110/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2086 _4436_/X VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6038__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1341 _4315_/B VGND VGND VPWR VPWR hold2850/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2097 hold143/X VGND VGND VPWR VPWR _4190_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1352 _4294_/B VGND VGND VPWR VPWR hold2816/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1363 _4317_/B VGND VGND VPWR VPWR hold2912/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1374 hold1412/X VGND VGND VPWR VPWR hold1413/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 hold2136/X VGND VGND VPWR VPWR hold2137/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1396 _6938_/Q VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__A1 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5677__C hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4581__C _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3811__A2 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3478__B hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6210__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6761__B2 _7025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input88_A spimemio_flash_io1_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3494__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3925__C _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6513__A1 _7465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5316__A2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6513__B2 _7505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6277__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3660__C _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6292__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3669__A _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5587__C _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3940_ _7567_/Q _5911_/A _5992_/C _3501_/X _7575_/Q VGND VGND VPWR VPWR _3940_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4491__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3871_ input47/X _4248_/S _4467_/A _7128_/Q _3870_/X VGND VGND VPWR VPWR _3871_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6201__B1 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5884__A _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5610_ _5610_/A0 _5954_/A1 _5611_/S VGND VGND VPWR VPWR _5610_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6590_ _7348_/Q _6452_/X _6467_/X _7420_/Q _6589_/X VGND VGND VPWR VPWR _6590_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3566__A1 _7366_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3566__B2 _7470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5541_ _4955_/X _5459_/X _5541_/C _5541_/D VGND VGND VPWR VPWR _5543_/B sky130_fd_sc_hd__and4bb_1
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2457_A _6991_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5472_ _4774_/Y _5471_/X _5386_/X _5256_/X _5267_/X VGND VGND VPWR VPWR _5474_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6504__B2 _7481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7211_ _7211_/CLK _7211_/D fanout574/X VGND VGND VPWR VPWR _7211_/Q sky130_fd_sc_hd__dfstp_1
X_4423_ _4423_/A0 _4422_/X _4423_/S VGND VGND VPWR VPWR _4423_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5823__S _5829_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7142_ _7144_/CLK _7142_/D fanout567/X VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfrtp_4
X_4354_ _4354_/A0 _5583_/A0 _4357_/S VGND VGND VPWR VPWR _4354_/X sky130_fd_sc_hd__mux2_1
Xfanout417 hold21/X VGND VGND VPWR VPWR _5722_/A sky130_fd_sc_hd__buf_12
Xfanout439 _6056_/X VGND VGND VPWR VPWR _6600_/B sky130_fd_sc_hd__buf_12
X_7073_ _4127_/A1 _7073_/D _6863_/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_4
X_4285_ _4289_/S _4285_/B VGND VGND VPWR VPWR _4285_/Y sky130_fd_sc_hd__nand2_1
X_6024_ _7589_/Q _7588_/Q VGND VGND VPWR VPWR _6121_/A sky130_fd_sc_hd__and2_4
XFILLER_0_146_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _6926_/CLK _6926_/D fanout565/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_77_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout442_A _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6857_ _6873_/A _6869_/B VGND VGND VPWR VPWR _6857_/X sky130_fd_sc_hd__and2_1
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5794__A _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5808_ _5808_/A0 hold84/X _5811_/S VGND VGND VPWR VPWR _5808_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6788_ _6792_/S _6788_/B VGND VGND VPWR VPWR _6788_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_161_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5739_ _5739_/A0 _5955_/A1 _5739_/S VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4203__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6121__C _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7409_ _7409_/CLK _7409_/D fanout577/X VGND VGND VPWR VPWR _7409_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5733__S _5739_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold460 hold460/A VGND VGND VPWR VPWR hold460/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6510__A4 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold471 hold471/A VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4857__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold482 hold482/A VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6259__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold493 _5901_/X VGND VGND VPWR VPWR _7494_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5034__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input142_A wb_dat_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6274__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 hold1160/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
Xhold1171 hold3057/X VGND VGND VPWR VPWR hold3058/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1182 hold1182/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
XFILLER_0_169_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 hold2901/X VGND VGND VPWR VPWR hold1193/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__A1 _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5908__S _5910_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6734__B2 _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_180_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3655__C _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_356 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _4150_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3671__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4070_ hold59/A hold1/A _4075_/S VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_58_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2205_A _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4972_ _5113_/A _5094_/A _5399_/C _4846_/B VGND VGND VPWR VPWR _5324_/A sky130_fd_sc_hd__o211a_2
XFILLER_0_176_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3787__A1 _7247_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6711_ _7149_/Q _6408_/A _6424_/X _7129_/Q _6702_/X VGND VGND VPWR VPWR _6711_/X
+ sky130_fd_sc_hd__a221o_2
X_3923_ _7214_/Q _3922_/Y _3923_/S VGND VGND VPWR VPWR _3923_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5818__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6642_ _7486_/Q _6447_/C _6459_/C _6419_/C _7566_/Q VGND VGND VPWR VPWR _6642_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_184_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3854_ _3854_/A _3854_/B _3854_/C _3854_/D VGND VGND VPWR VPWR _3855_/C sky130_fd_sc_hd__and4_1
XFILLER_0_156_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6573_ _6572_/X _6598_/A2 _6573_/S VGND VGND VPWR VPWR _7619_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_116_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3785_ _7180_/Q _5938_/C _5619_/B _3675_/X _7190_/Q VGND VGND VPWR VPWR _3785_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_hold2741_A _7303_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3565__C _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5524_ _5107_/A _5282_/B wire529/X _5559_/C _5523_/X VGND VGND VPWR VPWR _5524_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_131_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6489__B1 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7203__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5455_ _4947_/Y _5245_/X _5366_/X VGND VGND VPWR VPWR _5543_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4406_ _4406_/A1 hold284/X _4168_/D _4422_/S VGND VGND VPWR VPWR _4406_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_0_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5386_ _4703_/Y _4844_/Y _4716_/Y _5563_/A1 VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_1_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3711__A1 input24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7125_ _7134_/CLK _7125_/D _6833_/A VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfrtp_4
X_4337_ hold470/X _5950_/A1 _4339_/S VGND VGND VPWR VPWR _4337_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout392_A hold2225/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7056_ _7170_/CLK _7056_/D fanout573/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_4
X_4268_ _4268_/A0 _5950_/A1 _4270_/S VGND VGND VPWR VPWR _4268_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_157_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6007_ _6932_/Q _6751_/S _6051_/C _7584_/Q _4117_/Y VGND VGND VPWR VPWR _6017_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__6661__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4199_ _4199_/A0 _7643_/Q _7084_/Q VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6116__C _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6909_ _4127_/A1 _6909_/D _6859_/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5728__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5519__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6413__A _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6192__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5029__A _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3055_A _7146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_10__f_wb_clk_i clkbuf_3_5_0_wb_clk_i/X VGND VGND VPWR VPWR _7636_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold290 hold290/A VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6652__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5207__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3769__A1 input29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__B2 _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__C1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3666__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6042__B _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4194__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3570_ _3491_/X _3570_/B _3570_/C VGND VGND VPWR VPWR _3570_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_180_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3682__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5240_ _5091_/A _5072_/B wire533/X _4879_/C VGND VGND VPWR VPWR _5243_/C sky130_fd_sc_hd__a22o_1
XANTENNA__6486__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4497__B _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2608 _7515_/Q VGND VGND VPWR VPWR hold620/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5171_ _5038_/A _4861_/X _5180_/A _5038_/C _4928_/B VGND VGND VPWR VPWR _5171_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2619 _5882_/X VGND VGND VPWR VPWR hold871/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4122_ _4004_/A _4076_/C _4121_/Y _4005_/C _4010_/Y VGND VGND VPWR VPWR _7074_/D
+ sky130_fd_sc_hd__a32o_1
Xhold1907 _5963_/X VGND VGND VPWR VPWR hold134/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5105__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1918 hold124/X VGND VGND VPWR VPWR _4257_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1929 _6916_/Q VGND VGND VPWR VPWR hold354/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6643__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4053_ _3998_/Y _4123_/B _4052_/X _4053_/B2 _4062_/A VGND VGND VPWR VPWR _6895_/D
+ sky130_fd_sc_hd__o221a_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_2
XFILLER_0_143_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4955_ _5248_/A _5248_/B _5094_/A _4953_/X _5222_/A VGND VGND VPWR VPWR _4955_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3906_ input15/X _3503_/X _3666_/X _7012_/Q _3905_/X VGND VGND VPWR VPWR _3913_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4886_ _5222_/A _5213_/B VGND VGND VPWR VPWR _4886_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6625_ _6624_/X _6649_/A1 _6777_/S VGND VGND VPWR VPWR _6625_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_144_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3837_ _3837_/A _3837_/B _3837_/C _3837_/D VGND VGND VPWR VPWR _3854_/B sky130_fd_sc_hd__nor4_1
XFILLER_0_74_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6174__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6713__A4 _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6556_ _7355_/Q _6459_/B _6459_/C _6420_/C _7395_/Q VGND VGND VPWR VPWR _6556_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_144_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3768_ _7418_/Q _5866_/B _4212_/A _3669_/X _6970_/Q VGND VGND VPWR VPWR _3768_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5507_ _4716_/Y _5065_/Y _5210_/X _5185_/C _5355_/A VGND VGND VPWR VPWR _5508_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__3932__B2 _7229_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6487_ _7296_/Q _6420_/A _6467_/X _7416_/Q _6486_/X VGND VGND VPWR VPWR _6494_/A
+ sky130_fd_sc_hd__a221o_1
X_3699_ _7355_/Q _5785_/A _4212_/A _3498_/X _7379_/Q VGND VGND VPWR VPWR _3699_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5438_ _5438_/A _5438_/B _5438_/C _5438_/D VGND VGND VPWR VPWR _5441_/C sky130_fd_sc_hd__and4_1
Xoutput340 hold2769/X VGND VGND VPWR VPWR hold1162/A sky130_fd_sc_hd__buf_6
XFILLER_0_100_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5685__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5369_ _4601_/Y _4956_/A _4956_/B _4960_/B VGND VGND VPWR VPWR _5457_/B sky130_fd_sc_hd__a31o_1
X_7108_ _7644_/CLK _7108_/D _4309_/B VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6634__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7039_ _7189_/CLK _7039_/D fanout572/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6408__A _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4660__A2 _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1791_A _7565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input105_A wb_adr_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3620__B1 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3486__B _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6165__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold3172_A _7407_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input70_A mgmt_gpio_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3923__A1 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6322__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3687__B1 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5222__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6640__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6752__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4780__B _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5600__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4740_ _4831_/A _4786_/C _4909_/D _4740_/D VGND VGND VPWR VPWR _5077_/B sky130_fd_sc_hd__and4bb_4
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3611__B1 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4671_ _4667_/A _4667_/B _4667_/C _4974_/D _4974_/B VGND VGND VPWR VPWR _5339_/D
+ sky130_fd_sc_hd__o311a_4
XFILLER_0_126_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6410_ _7594_/Q _6455_/B _6651_/B VGND VGND VPWR VPWR _6410_/X sky130_fd_sc_hd__and3_1
X_3622_ _7234_/Q _3617_/X _3618_/X _3616_/X _3621_/X VGND VGND VPWR VPWR _3623_/D
+ sky130_fd_sc_hd__a2111o_4
X_7390_ _7582_/CLK _7390_/D fanout584/X VGND VGND VPWR VPWR _7390_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_141_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6341_ _6332_/B _6333_/X _6340_/X _6339_/X VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_24_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3553_ hold22/A _5938_/B _5992_/C VGND VGND VPWR VPWR _4231_/S sky130_fd_sc_hd__and3_4
XANTENNA__4939__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2537_A _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6272_ _7358_/Q _6099_/X _6112_/X _7486_/Q _6271_/X VGND VGND VPWR VPWR _6272_/X
+ sky130_fd_sc_hd__a221o_1
X_3484_ _3507_/A _3576_/C _5830_/C VGND VGND VPWR VPWR _5911_/A sky130_fd_sc_hd__and3_4
XFILLER_0_122_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3106 _7021_/Q VGND VGND VPWR VPWR hold3106/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5667__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3117 hold3117/A VGND VGND VPWR VPWR _5831_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5223_ _5223_/A _5223_/B _5223_/C _5223_/D VGND VGND VPWR VPWR _5224_/C sky130_fd_sc_hd__nand4_1
Xhold3128 _7142_/Q VGND VGND VPWR VPWR hold3128/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3139 _7177_/Q VGND VGND VPWR VPWR hold3139/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2405 _4269_/X VGND VGND VPWR VPWR hold2405/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5831__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2416 _7139_/Q VGND VGND VPWR VPWR hold993/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2427 hold684/X VGND VGND VPWR VPWR _5645_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_44_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5154_ _4687_/Y _4793_/Y _4821_/Y _4796_/Y _4723_/Y VGND VGND VPWR VPWR _5156_/B
+ sky130_fd_sc_hd__o32a_1
Xhold2438 _7236_/Q VGND VGND VPWR VPWR hold645/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_47_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2449 hold653/X VGND VGND VPWR VPWR _4469_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1704 _5941_/X VGND VGND VPWR VPWR hold313/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1715 _7298_/Q VGND VGND VPWR VPWR hold306/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6616__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4105_ _6427_/A _4105_/B VGND VGND VPWR VPWR _4105_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3693__A3 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1726 _4541_/X VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4447__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1737 hold408/X VGND VGND VPWR VPWR _4385_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5085_ _5222_/A _5387_/C _4765_/B _5084_/Y VGND VGND VPWR VPWR _5085_/Y sky130_fd_sc_hd__a31oi_1
Xhold1748 hold296/X VGND VGND VPWR VPWR _5978_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1759 hold67/X VGND VGND VPWR VPWR _5994_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4036_ _4036_/A0 _4035_/X _4040_/A VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3850__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4690__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6395__A2 _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5987_ _5987_/A0 _5987_/A1 _5991_/S VGND VGND VPWR VPWR _5987_/X sky130_fd_sc_hd__mux2_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4938_ _4882_/Y _4936_/Y _4937_/Y _4934_/Y VGND VGND VPWR VPWR _4941_/C sky130_fd_sc_hd__o211ai_1
XANTENNA__3602__B1 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_30 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4646_/A _4869_/A2 _4617_/Y _4860_/B VGND VGND VPWR VPWR _4889_/B sky130_fd_sc_hd__o211ai_4
X_7657_ _7657_/A VGND VGND VPWR VPWR _7657_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_52 _3575_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _7174_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4158__A1 _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _7389_/Q _6413_/C _6426_/X _6451_/X _7485_/Q VGND VGND VPWR VPWR _6608_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_74 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7588_ _7610_/CLK _7588_/D fanout567/X VGND VGND VPWR VPWR _7588_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_105_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3905__A1 _7158_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6539_ _7546_/Q _6419_/A _6435_/X _7514_/Q _6538_/X VGND VGND VPWR VPWR _6544_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4849__C _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5741__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput181 _3430_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3420_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XANTENNA__4330__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6607__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3684__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2950 hold2950/A VGND VGND VPWR VPWR _5867_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2961 hold2961/A VGND VGND VPWR VPWR _5913_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2972 _4267_/X VGND VGND VPWR VPWR hold2972/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2983 _4511_/X VGND VGND VPWR VPWR hold2983/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2994 hold2994/A VGND VGND VPWR VPWR _4523_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6083__B2 _7319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7377__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6386__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3497__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4105__B _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6138__A2 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_170_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4149__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6689__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output274_A _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3663__C _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__A2 _6072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4609__C1 _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4085__B1 _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5910_ _5991_/A1 _5910_/A1 _5910_/S VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_159_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6890_ _7075_/CLK _6890_/D _6840_/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3832__B1 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5841_ _5841_/A0 _5985_/A1 _5847_/S VGND VGND VPWR VPWR _5841_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5585__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2487_A _7138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5772_ _5772_/A0 _5997_/A1 _5775_/S VGND VGND VPWR VPWR _5772_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7511_ _7560_/CLK _7511_/D fanout599/X VGND VGND VPWR VPWR _7511_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4723_ _5387_/C _4815_/B VGND VGND VPWR VPWR _4723_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_29_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6129__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5826__S _5829_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2654_A _7459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7442_ _7513_/CLK _7442_/D fanout600/X VGND VGND VPWR VPWR _7442_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4654_ _4644_/Y _4646_/Y _4823_/C VGND VGND VPWR VPWR _4654_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_142_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5888__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_4
XFILLER_0_4_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3605_ input9/X _3486_/X _3508_/X _7557_/Q _3604_/X VGND VGND VPWR VPWR _3606_/D
+ sky130_fd_sc_hd__a221o_1
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_2
X_7373_ _7429_/CLK _7373_/D fanout583/X VGND VGND VPWR VPWR _7373_/Q sky130_fd_sc_hd__dfrtp_4
X_4585_ _4675_/B _4643_/C _5038_/A _5089_/B VGND VGND VPWR VPWR _4585_/Y sky130_fd_sc_hd__nand4_2
Xhold801 hold801/A VGND VGND VPWR VPWR hold801/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold812 hold812/A VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2821_A _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold823 hold823/A VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_4
Xinput94 uart_enabled VGND VGND VPWR VPWR _4173_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6324_ _7007_/Q _6082_/X _6094_/X _7210_/Q _6323_/X VGND VGND VPWR VPWR _6327_/C
+ sky130_fd_sc_hd__a221o_1
Xhold834 hold834/A VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3536_ _7494_/Q _3496_/Y hold12/A _3535_/X _7486_/Q VGND VGND VPWR VPWR _3536_/X
+ sky130_fd_sc_hd__a32o_1
Xhold845 hold845/A VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap553 _5395_/A1 VGND VGND VPWR VPWR _5401_/A3 sky130_fd_sc_hd__clkbuf_2
Xhold856 hold856/A VGND VGND VPWR VPWR hold856/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold867 hold867/A VGND VGND VPWR VPWR _7254_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold878 hold878/A VGND VGND VPWR VPWR hold878/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4388__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold889 hold889/A VGND VGND VPWR VPWR hold889/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6255_ _7325_/Q _6082_/X _6110_/X _7437_/Q _6254_/X VGND VGND VPWR VPWR _6255_/X
+ sky130_fd_sc_hd__a221o_1
X_3467_ _4429_/B _3468_/A2 hold154/X _3465_/Y VGND VGND VPWR VPWR _3467_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__6301__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2202 _7302_/Q VGND VGND VPWR VPWR hold458/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5206_ _5202_/X _5204_/X _5205_/X VGND VGND VPWR VPWR _5206_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2213 _5874_/X VGND VGND VPWR VPWR hold544/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2224 _3454_/X VGND VGND VPWR VPWR _3485_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_6186_ _7498_/Q _6085_/X _6112_/X _7482_/Q _6185_/X VGND VGND VPWR VPWR _6186_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2235 hold540/X VGND VGND VPWR VPWR _5949_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1501 _5845_/X VGND VGND VPWR VPWR hold174/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2246 _5679_/X VGND VGND VPWR VPWR hold537/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1512 _7564_/Q VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5137_ _4695_/Y _4735_/Y _4821_/Y _4687_/Y VGND VGND VPWR VPWR _5139_/C sky130_fd_sc_hd__a211o_1
Xhold2257 hold532/X VGND VGND VPWR VPWR _5715_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2268 _7539_/Q VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout472_A _4256_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1523 hold203/X VGND VGND VPWR VPWR _5662_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1534 hold29/X VGND VGND VPWR VPWR _5838_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2279 hold557/X VGND VGND VPWR VPWR _5856_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1545 _7580_/Q VGND VGND VPWR VPWR hold207/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1556 _7666_/A VGND VGND VPWR VPWR hold195/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_165_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1567 hold219/X VGND VGND VPWR VPWR _5854_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5068_ _5091_/C _5068_/B _5453_/C VGND VGND VPWR VPWR _5573_/D sky130_fd_sc_hd__nand3_1
XANTENNA__6604__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1578 hold1578/A VGND VGND VPWR VPWR _6000_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1589 _7377_/Q VGND VGND VPWR VPWR hold239/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4019_ _4040_/D _4014_/B _3450_/X _4017_/Y VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_149_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6368__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4379__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5736__S _5739_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5879__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6540__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input33_A mask_rev_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3930__D _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2780 hold2780/A VGND VGND VPWR VPWR _4353_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2791 hold2791/A VGND VGND VPWR VPWR hold2791/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5203__C _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6359__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3658__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4116__A _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5646__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3593__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3674__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6050__B _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold108 hold108/A VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6531__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold119 hold119/A VGND VGND VPWR VPWR _7533_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4542__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4370_ _4370_/A _4551_/D VGND VGND VPWR VPWR _4375_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_21_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _7593_/Q _6051_/C _6929_/Q VGND VGND VPWR VPWR _6040_/Y sky130_fd_sc_hd__nor3_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6942_ _7278_/CLK _6942_/D fanout580/X VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6873_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6873_/X sky130_fd_sc_hd__and2_1
XANTENNA__3820__A3 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5824_ _5824_/A0 _5896_/A0 _5829_/S VGND VGND VPWR VPWR _5824_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_174_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5755_ _5755_/A0 _5953_/A1 _5757_/S VGND VGND VPWR VPWR _5755_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6770__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4706_ _4706_/A _5260_/C VGND VGND VPWR VPWR _4706_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_173_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3584__A2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5686_ _5686_/A hold47/X VGND VGND VPWR VPWR _5694_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_127_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7425_ _7489_/CLK _7425_/D fanout586/X VGND VGND VPWR VPWR _7425_/Q sky130_fd_sc_hd__dfrtp_2
X_4637_ _4984_/B _4814_/C VGND VGND VPWR VPWR _4836_/C sky130_fd_sc_hd__nor2_8
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold620 hold620/A VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold631 hold631/A VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7356_ _7429_/CLK _7356_/D fanout583/X VGND VGND VPWR VPWR _7356_/Q sky130_fd_sc_hd__dfrtp_4
X_4568_ _4795_/C _4984_/B VGND VGND VPWR VPWR _4568_/Y sky130_fd_sc_hd__nand2_4
Xhold642 _4499_/X VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold653 hold653/A VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6307_ _6306_/X _6330_/A2 _6777_/S VGND VGND VPWR VPWR _6307_/X sky130_fd_sc_hd__mux2_1
Xhold664 hold664/A VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3519_ hold22/A _3519_/B _4491_/C VGND VGND VPWR VPWR _3519_/X sky130_fd_sc_hd__and3_2
Xhold675 hold675/A VGND VGND VPWR VPWR _7230_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7287_ _7363_/CLK _7287_/D fanout575/X VGND VGND VPWR VPWR _7287_/Q sky130_fd_sc_hd__dfstp_2
Xhold686 hold686/A VGND VGND VPWR VPWR hold686/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4499_ _5940_/A1 _4499_/A1 _4502_/S VGND VGND VPWR VPWR _4499_/X sky130_fd_sc_hd__mux2_1
Xhold697 _4330_/X VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6238_ _6260_/A2 _4116_/X _6067_/X _6237_/X VGND VGND VPWR VPWR _7607_/D sky130_fd_sc_hd__o31a_1
Xhold2010 _7003_/Q VGND VGND VPWR VPWR hold596/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2021 _7345_/Q VGND VGND VPWR VPWR hold559/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2032 _4555_/X VGND VGND VPWR VPWR hold443/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2043 hold578/X VGND VGND VPWR VPWR _5626_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6649_/S _6169_/A2 _6777_/S _6168_/X VGND VGND VPWR VPWR _6169_/X sky130_fd_sc_hd__a211o_1
Xhold2054 hold565/X VGND VGND VPWR VPWR _5708_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 _4192_/X VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2065 _7528_/Q VGND VGND VPWR VPWR hold542/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1331 hold3168/X VGND VGND VPWR VPWR hold3169/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6119__C _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2076 hold110/X VGND VGND VPWR VPWR _5943_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2087 _7242_/Q VGND VGND VPWR VPWR hold623/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1342 _4310_/B VGND VGND VPWR VPWR hold2819/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2098 _4190_/X VGND VGND VPWR VPWR hold144/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1353 _6784_/B VGND VGND VPWR VPWR hold2824/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1364 _6781_/B VGND VGND VPWR VPWR hold2916/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1375 hold1414/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6589__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1386 hold1926/X VGND VGND VPWR VPWR hold1927/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5797__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1397 hold90/X VGND VGND VPWR VPWR _4228_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7572_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4581__D _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1871_A _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3811__A3 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3478__C _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7309_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6761__A2 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3575__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3494__B _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3925__D _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6513__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3252_A _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5721__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4524__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4742__A_N _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6277__A1 _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4288__A0 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6682__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output237_A _4148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7321__RESET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4772__C _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3669__B _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5587__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4491__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3870_ _7138_/Q _4491_/B _4521_/B hold72/A _7560_/Q VGND VGND VPWR VPWR _3870_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6201__A1 _7451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4280__S _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2185_A _7294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3566__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5540_ _4953_/X _4956_/Y _5248_/X _5371_/X _4959_/X VGND VGND VPWR VPWR _5541_/C
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5471_ _4743_/A _4747_/B _5073_/A _4748_/Y VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__o31a_2
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4422_ _4448_/A0 _5991_/A1 _4422_/S VGND VGND VPWR VPWR _4422_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5712__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7210_ _7213_/CLK _7210_/D fanout590/X VGND VGND VPWR VPWR _7210_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7141_ _7197_/CLK _7141_/D fanout601/X VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_4
X_4353_ _4353_/A0 _5840_/A1 _4357_/S VGND VGND VPWR VPWR _4353_/X sky130_fd_sc_hd__mux2_1
Xfanout407 hold1467/X VGND VGND VPWR VPWR _3931_/D sky130_fd_sc_hd__buf_12
XANTENNA__6000__S hold37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout418 hold21/X VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__buf_8
X_7072_ _4127_/A1 _7072_/D _6862_/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_1
X_4284_ _4289_/S _3795_/B _4283_/Y VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__o21ai_1
X_6023_ _7589_/Q _7588_/Q VGND VGND VPWR VPWR _6023_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5779__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6926_/CLK _6925_/D fanout565/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_159_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout435_A _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6856_ _6873_/A _6872_/B VGND VGND VPWR VPWR _6856_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5794__B hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5807_ _5807_/A0 _5951_/A1 _5811_/S VGND VGND VPWR VPWR _5807_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3999_ _7071_/Q _7074_/Q _7073_/Q _6908_/Q VGND VGND VPWR VPWR _4006_/A sky130_fd_sc_hd__o31a_2
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6743__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6787_ _6792_/S _3795_/B _6786_/Y VGND VGND VPWR VPWR _7632_/D sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout602_A fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5738_ _5738_/A0 _5954_/A1 _5739_/S VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5669_ _5903_/A0 _5669_/A1 _5670_/S VGND VGND VPWR VPWR _5669_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4506__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7408_ _7409_/CLK _7408_/D fanout577/X VGND VGND VPWR VPWR _7408_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_32_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold450 hold450/A VGND VGND VPWR VPWR hold450/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7339_ _7499_/CLK _7339_/D fanout578/X VGND VGND VPWR VPWR _7339_/Q sky130_fd_sc_hd__dfrtp_4
Xhold461 _5739_/X VGND VGND VPWR VPWR _7350_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold472 hold472/A VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold483 hold483/A VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold494 hold494/A VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input135_A wb_dat_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 _4457_/X VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1161 hold2768/X VGND VGND VPWR VPWR hold2769/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1172 _4402_/X VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1183 hold2838/X VGND VGND VPWR VPWR hold1183/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 hold1194/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5050__A _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__A2 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6195__B1 _6116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6734__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3655__D _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7573__RESET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3671__C _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3720__A2 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_max_cap400_A _4758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4971_ _4571_/Y _4843_/A _4709_/Y VGND VGND VPWR VPWR _4971_/X sky130_fd_sc_hd__o21a_4
XFILLER_0_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6710_ _7018_/Q _6425_/X _6454_/X _7068_/Q _6709_/X VGND VGND VPWR VPWR _6710_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3787__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3922_ _3922_/A _3922_/B _3922_/C VGND VGND VPWR VPWR _3922_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3853_ _7023_/Q _3667_/X _3849_/X _3850_/X _3852_/X VGND VGND VPWR VPWR _3854_/D
+ sky130_fd_sc_hd__a2111oi_2
X_6641_ _7326_/Q _6421_/X _6462_/X _7366_/Q _6640_/X VGND VGND VPWR VPWR _6647_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6186__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3619__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5528__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5933__A0 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3539__A2 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6572_ _6649_/S _6572_/A2 _6570_/Y _6571_/X VGND VGND VPWR VPWR _6572_/X sky130_fd_sc_hd__a22o_1
X_3784_ _7538_/Q _3590_/C _5938_/C _3565_/X _7466_/Q VGND VGND VPWR VPWR _3792_/B
+ sky130_fd_sc_hd__a32o_2
XANTENNA__3944__C1 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5523_ _5282_/B _5399_/C _5113_/B _5324_/A VGND VGND VPWR VPWR _5523_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5834__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2734_A _7279_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5454_ _5180_/B _4935_/X _5238_/X _5453_/X _5347_/X VGND VGND VPWR VPWR _5545_/C
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3862__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4405_ _4405_/A0 _5586_/A0 _4405_/S VGND VGND VPWR VPWR _4405_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5161__A1 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5385_ _5222_/A _4702_/Y _4755_/C _5453_/C _5086_/B VGND VGND VPWR VPWR _5385_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_10_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3711__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4336_ _4336_/A0 _5583_/A0 _4339_/S VGND VGND VPWR VPWR _4336_/X sky130_fd_sc_hd__mux2_1
X_7124_ _7134_/CLK _7124_/D _6833_/A VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_5_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7055_ _7213_/CLK _7055_/D fanout590/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4267_ _4267_/A0 _5583_/A0 _4270_/S VGND VGND VPWR VPWR _4267_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout385_A _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6006_ _6006_/A _7584_/Q VGND VGND VPWR VPWR _6006_/X sky130_fd_sc_hd__and2_1
XANTENNA__6661__A1 _6967_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4198_ _4198_/A0 _5863_/A0 _4202_/S VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3475__A1 _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4185__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6908_ _4127_/A1 _6908_/D _6858_/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3778__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6839_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6839_/X sky130_fd_sc_hd__and2_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6177__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6413__B _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6716__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5924__A0 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5744__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3950__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold280 _3500_/C VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3702__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold291 hold291/A VGND VGND VPWR VPWR _7386_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6101__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6652__A1 _7137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6652__B2 _7187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5207__A2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__A2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6707__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3666__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5391__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3941__A2 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4778__B _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3682__B _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6340__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5170_ _5339_/D _5180_/B _5030_/C _5039_/B VGND VGND VPWR VPWR _5170_/X sky130_fd_sc_hd__a31o_1
Xhold2609 hold620/X VGND VGND VPWR VPWR _5925_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4121_ _4121_/A _6882_/Q VGND VGND VPWR VPWR _4121_/Y sky130_fd_sc_hd__nor2_1
Xhold1908 _7418_/Q VGND VGND VPWR VPWR hold366/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1919 _4257_/X VGND VGND VPWR VPWR hold125/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4052_ _7071_/Q _7074_/Q _7073_/Q _6893_/Q VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__o31a_1
XANTENNA__6643__B2 _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3457__A1 _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4406__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5829__S _5829_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4954_ _4954_/A _5248_/A _4954_/C VGND VGND VPWR VPWR _4960_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3905_ _7158_/Q _5947_/B _5632_/B _3544_/X _7416_/Q VGND VGND VPWR VPWR _3905_/X
+ sky130_fd_sc_hd__a32o_1
X_7673_ _7673_/A VGND VGND VPWR VPWR _7673_/X sky130_fd_sc_hd__clkbuf_2
X_4885_ _5222_/A _4942_/A _4948_/C VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__and3_1
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5906__A0 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6624_ _6649_/S _7620_/Q _6622_/X _6623_/X VGND VGND VPWR VPWR _6624_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold2949_A _7463_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3836_ _7237_/Q _3515_/X _4394_/A _7063_/Q _3835_/X VGND VGND VPWR VPWR _3837_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6174__A3 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5382__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3767_ _7330_/Q _5713_/A _3562_/X _7298_/Q _3766_/X VGND VGND VPWR VPWR _3767_/X
+ sky130_fd_sc_hd__a221o_1
X_6555_ _7435_/Q _6747_/B _6645_/C _6460_/X _7387_/Q VGND VGND VPWR VPWR _6555_/X
+ sky130_fd_sc_hd__a32o_1
X_5506_ _5205_/X _5506_/B _5506_/C _5506_/D VGND VGND VPWR VPWR _5550_/C sky130_fd_sc_hd__and4b_2
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3932__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6486_ _7368_/Q _6413_/C _6651_/C _6422_/X _7288_/Q VGND VGND VPWR VPWR _6486_/X
+ sky130_fd_sc_hd__a32o_1
X_3698_ _7395_/Q _3473_/X _4533_/A _7186_/Q _3697_/X VGND VGND VPWR VPWR _3698_/X
+ sky130_fd_sc_hd__a221o_1
X_5437_ _5203_/B _5329_/X _5436_/X VGND VGND VPWR VPWR _5438_/D sky130_fd_sc_hd__a21oi_2
Xoutput330 hold1191/X VGND VGND VPWR VPWR hold1192/A sky130_fd_sc_hd__buf_6
Xoutput341 hold1179/X VGND VGND VPWR VPWR hold1180/A sky130_fd_sc_hd__buf_6
XFILLER_0_11_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5368_ _4654_/Y _4936_/Y _5245_/X _5419_/A VGND VGND VPWR VPWR _5512_/A sky130_fd_sc_hd__o31a_2
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7107_ _4164_/A1 _7107_/D _4309_/B VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_4
X_4319_ _3643_/Y _4319_/A1 _4321_/S VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__mux2_1
X_5299_ _5451_/A1 _4722_/Y _4737_/Y _4746_/Y _5298_/X VGND VGND VPWR VPWR _5538_/A
+ sky130_fd_sc_hd__o311a_1
XANTENNA__6229__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6634__A1 _7334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7038_ _7189_/CLK _7038_/D fanout572/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__6408__B _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3853__D1 _3852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4660__A3 _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5739__S _5739_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__B1 _4940_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3620__A1 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3486__C _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6165__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5373__A1 _4744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4598__B _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input63_A mgmt_gpio_in[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6322__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout590 fanout606/X VGND VGND VPWR VPWR fanout590/X sky130_fd_sc_hd__buf_12
XFILLER_0_88_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5649__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4670_ _4568_/Y _4984_/C _4740_/D VGND VGND VPWR VPWR _4974_/D sky130_fd_sc_hd__o21ai_4
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3621_ _7404_/Q _5794_/A _3542_/X _6924_/Q _3620_/X VGND VGND VPWR VPWR _3621_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5364__A1 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6561__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4789__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3552_ _5640_/B _5612_/C _5614_/B VGND VGND VPWR VPWR _4248_/S sky130_fd_sc_hd__and3_4
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6340_ _7179_/Q _6092_/X _6119_/X _7134_/Q _6334_/X VGND VGND VPWR VPWR _6340_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3914__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6271_ _7430_/Q _7592_/Q _6074_/X _6120_/X _7342_/Q VGND VGND VPWR VPWR _6271_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5116__A1 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6313__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3483_ _3505_/C _3505_/D VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__and2b_1
XANTENNA__5116__B2 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5222_ _5222_/A _5222_/B _5222_/C _5387_/D VGND VGND VPWR VPWR _5223_/C sky130_fd_sc_hd__nand4_1
Xhold3107 hold3107/A VGND VGND VPWR VPWR _4347_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3118 _5831_/X VGND VGND VPWR VPWR hold3118/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3129 hold3129/A VGND VGND VPWR VPWR _4486_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2406 _7441_/Q VGND VGND VPWR VPWR hold943/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5153_ _5153_/A _5153_/B _5153_/C VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__and3_1
Xhold2417 hold993/X VGND VGND VPWR VPWR _4482_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2428 _7184_/Q VGND VGND VPWR VPWR hold937/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2439 hold645/X VGND VGND VPWR VPWR _5605_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1705 _7370_/Q VGND VGND VPWR VPWR hold288/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4104_ _7593_/Q _6462_/D _6435_/B _7594_/Q VGND VGND VPWR VPWR _4105_/B sky130_fd_sc_hd__and4bb_4
Xhold1716 hold306/X VGND VGND VPWR VPWR _5681_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6616__A1 _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5084_ _5084_/A _5467_/A _5084_/C _5084_/D VGND VGND VPWR VPWR _5084_/Y sky130_fd_sc_hd__nand4_1
Xhold1727 hold58/X VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1738 _4385_/X VGND VGND VPWR VPWR hold409/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1749 _5978_/X VGND VGND VPWR VPWR hold297/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_79_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4035_ _6902_/Q _4025_/A _4025_/Y _4034_/X VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_189_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _5986_/A0 _5986_/A1 _5991_/S VGND VGND VPWR VPWR _5986_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6395__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4937_ _4954_/A _5453_/A _4937_/C _4940_/D VGND VGND VPWR VPWR _4937_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_136_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3602__B2 _7309_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7656_ _7656_/A VGND VGND VPWR VPWR _7656_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_31 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4571_/Y _4646_/A _5387_/B _4617_/Y _4860_/B VGND VGND VPWR VPWR _5213_/C
+ sky130_fd_sc_hd__o311a_4
XFILLER_0_47_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_42 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _3583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4158__A2 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _7357_/Q _6413_/C _6459_/C _6408_/B _7381_/Q VGND VGND VPWR VPWR _6607_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_64 input72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ _7497_/Q _5902_/A _3812_/X _3813_/X _3818_/X VGND VGND VPWR VPWR _3855_/B
+ sky130_fd_sc_hd__a2111oi_2
XANTENNA__6552__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4699__A _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7587_ _7601_/CLK _7587_/D _4128_/B VGND VGND VPWR VPWR _7587_/Q sky130_fd_sc_hd__dfrtp_4
X_4799_ _5387_/C _4815_/B _4799_/C VGND VGND VPWR VPWR _4800_/B sky130_fd_sc_hd__and3_1
XFILLER_0_105_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3905__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6538_ _7330_/Q _4105_/B _6459_/B _6420_/B _7306_/Q VGND VGND VPWR VPWR _6538_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6410__C _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6469_ _7367_/Q _6459_/B _6429_/X _6468_/X _7407_/Q VGND VGND VPWR VPWR _6469_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput171 _4175_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
XFILLER_0_100_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput182 _3429_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput193 _3419_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_0_100_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6419__A _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2940 hold2940/A VGND VGND VPWR VPWR _5621_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2951 _5867_/X VGND VGND VPWR VPWR _7463_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2962 _7168_/Q VGND VGND VPWR VPWR hold2962/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2973 _7133_/Q VGND VGND VPWR VPWR hold2973/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4584__D _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2984 _6875_/Q VGND VGND VPWR VPWR hold2984/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2995 _4523_/X VGND VGND VPWR VPWR hold2995/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3841__A1 _7393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3841__B2 _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3497__B _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5594__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6791__A0 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3282_A _7391_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5346__A1 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6543__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__C1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4609__B1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4085__A1 _6895_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5840_ _5840_/A0 _5840_/A1 _5847_/S VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_185_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5771_ _5771_/A0 _5987_/A1 _5775_/S VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_174_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7510_ _7510_/CLK _7510_/D fanout603/X VGND VGND VPWR VPWR _7510_/Q sky130_fd_sc_hd__dfrtp_4
X_4722_ _5399_/A _5399_/B VGND VGND VPWR VPWR _4722_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_72_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6129__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7441_ _7447_/CLK _7441_/D fanout598/X VGND VGND VPWR VPWR _7441_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6534__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4653_ _4644_/Y _4646_/Y _4823_/C VGND VGND VPWR VPWR _5248_/A sky130_fd_sc_hd__o21a_4
XFILLER_0_126_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__buf_2
X_3604_ _7429_/Q _4509_/A hold12/A _3562_/X _7301_/Q VGND VGND VPWR VPWR _3604_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_2
X_7372_ _7478_/CLK _7372_/D fanout583/X VGND VGND VPWR VPWR _7372_/Q sky130_fd_sc_hd__dfrtp_4
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR _3859_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4584_ _4675_/A _4675_/B _4643_/C _5038_/A VGND VGND VPWR VPWR _4593_/A sky130_fd_sc_hd__nand4_4
Xhold802 _5900_/X VGND VGND VPWR VPWR _7493_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3899__A1 _7488_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _4134_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold813 hold813/A VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_4
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_2
Xhold824 hold824/A VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6323_ _7133_/Q _6091_/X _6144_/C _6322_/X VGND VGND VPWR VPWR _6323_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold835 hold835/A VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3535_ hold22/A _5938_/C _3931_/D VGND VGND VPWR VPWR _3535_/X sky130_fd_sc_hd__and3_4
Xmax_cap554 _5134_/A VGND VGND VPWR VPWR _5395_/A1 sky130_fd_sc_hd__clkbuf_2
Xhold846 _5610_/X VGND VGND VPWR VPWR _7241_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold857 _4381_/X VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_149_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold868 hold868/A VGND VGND VPWR VPWR hold868/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6254_ _7405_/Q _6091_/X _6116_/B _7469_/Q _6087_/X VGND VGND VPWR VPWR _6254_/X
+ sky130_fd_sc_hd__a32o_1
X_3466_ hold153/X _4025_/A _4429_/B VGND VGND VPWR VPWR _3466_/X sky130_fd_sc_hd__o21ba_1
Xhold879 hold879/A VGND VGND VPWR VPWR hold879/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6301__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2203 hold458/X VGND VGND VPWR VPWR _5685_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5205_ _5205_/A1 _5107_/A _5061_/B _4969_/Y VGND VGND VPWR VPWR _5205_/X sky130_fd_sc_hd__a31o_1
Xhold2214 _7332_/Q VGND VGND VPWR VPWR hold891/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6185_ _7458_/Q _6094_/A _6079_/X _6094_/X _7506_/Q VGND VGND VPWR VPWR _6185_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2225 _3564_/A VGND VGND VPWR VPWR hold2225/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2236 _7406_/Q VGND VGND VPWR VPWR hold454/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1502 hold174/X VGND VGND VPWR VPWR _7444_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2247 _7398_/Q VGND VGND VPWR VPWR hold610/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5136_ _4687_/Y _5135_/Y _5134_/X VGND VGND VPWR VPWR _5139_/B sky130_fd_sc_hd__o21ba_1
Xhold2258 _7542_/Q VGND VGND VPWR VPWR hold534/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1513 hold209/X VGND VGND VPWR VPWR _5980_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2269 hold92/X VGND VGND VPWR VPWR _5952_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1524 _5662_/X VGND VGND VPWR VPWR hold204/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_165_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1535 _5838_/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1546 hold207/X VGND VGND VPWR VPWR _5998_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1557 hold195/X VGND VGND VPWR VPWR _4434_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5067_ _5091_/C _5260_/C _5453_/C VGND VGND VPWR VPWR _5067_/X sky130_fd_sc_hd__and3_1
Xhold1568 _5854_/X VGND VGND VPWR VPWR hold220/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1579 _6000_/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout465_A hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5273__B1 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_csclk_A _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4018_ hold51/A _6905_/Q _6904_/Q _4025_/B _3451_/Y VGND VGND VPWR VPWR _4018_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3823__A1 _7465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3598__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3823__B2 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6405__C _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6368__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_164_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5969_ _5969_/A0 _5987_/A1 hold13/X VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__mux2_1
X_7639_ _7646_/CLK _7639_/D _4309_/B VGND VGND VPWR VPWR _7639_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6525__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6421__B _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1747_A _7562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4579__D _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input165_A wb_sel_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4854__A3 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input26_A mask_rev_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2770 _6967_/Q VGND VGND VPWR VPWR hold2770/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2781 _6973_/Q VGND VGND VPWR VPWR _4280_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2792 _7182_/Q VGND VGND VPWR VPWR hold2792/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_187_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3814__B2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4116__B _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7180__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3593__A3 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3674__C hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6531__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold109 hold109/A VGND VGND VPWR VPWR _7259_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6295__A2 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_csclk_A _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5255__B1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6941_ _7333_/CLK _6941_/D fanout582/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7268__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5270__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6872_ _6873_/A _6872_/B VGND VGND VPWR VPWR _6872_/X sky130_fd_sc_hd__and2_1
X_5823_ _5823_/A0 _5967_/A1 _5829_/S VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6755__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5558__B2 _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5837__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5754_ _5754_/A0 _5754_/A1 _5757_/S VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3865__B hold36/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4705_ _4825_/A _5115_/A _5089_/B VGND VGND VPWR VPWR _4705_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_0_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6507__B1 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5685_ _5685_/A0 _5955_/A1 _5685_/S VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2931_A _7376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7424_ _7476_/CLK _7424_/D fanout586/X VGND VGND VPWR VPWR _7424_/Q sky130_fd_sc_hd__dfstp_2
X_4636_ _4814_/C _5301_/A1 _4772_/A VGND VGND VPWR VPWR _4636_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold610 hold610/A VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold621 _5925_/X VGND VGND VPWR VPWR _7515_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5730__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7355_ _7563_/CLK _7355_/D fanout599/X VGND VGND VPWR VPWR _7355_/Q sky130_fd_sc_hd__dfrtp_4
X_4567_ _4772_/A _4805_/B VGND VGND VPWR VPWR _4667_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold632 _5670_/X VGND VGND VPWR VPWR _7288_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold643 hold643/A VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap351 _5653_/S VGND VGND VPWR VPWR _5658_/S sky130_fd_sc_hd__buf_2
X_6306_ _6751_/S _7609_/Q _6304_/X _6305_/X VGND VGND VPWR VPWR _6306_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap362 _5127_/A VGND VGND VPWR VPWR _5205_/A1 sky130_fd_sc_hd__clkbuf_2
Xhold654 _4469_/X VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold665 _4205_/X VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3518_ _5785_/A hold22/A _5830_/C VGND VGND VPWR VPWR _5758_/A sky130_fd_sc_hd__and3_4
X_7286_ _7309_/CLK _7286_/D fanout579/X VGND VGND VPWR VPWR _7286_/Q sky130_fd_sc_hd__dfrtp_4
Xhold676 hold676/A VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4498_ _5840_/A1 _4498_/A1 _4502_/S VGND VGND VPWR VPWR _4498_/X sky130_fd_sc_hd__mux2_1
Xhold687 _5751_/X VGND VGND VPWR VPWR _7360_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_110_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap395 _4850_/B VGND VGND VPWR VPWR _4849_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__6286__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold698 hold698/A VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6237_ _6649_/S _6237_/A2 _6777_/S _6236_/X VGND VGND VPWR VPWR _6237_/X sky130_fd_sc_hd__a211o_1
XANTENNA_fanout582_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3449_ _3449_/A0 hold279/X _4429_/B VGND VGND VPWR VPWR _3449_/X sky130_fd_sc_hd__mux2_1
Xhold2000 hold440/X VGND VGND VPWR VPWR _5834_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2011 hold596/X VGND VGND VPWR VPWR _4325_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4297__A1 _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2022 hold559/X VGND VGND VPWR VPWR _5734_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2033 _7120_/Q VGND VGND VPWR VPWR hold486/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2044 _5626_/X VGND VGND VPWR VPWR hold579/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6036_/Y _7281_/Q _6167_/X _6157_/Y _6775_/B1 VGND VGND VPWR VPWR _6168_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 hold3135/X VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2055 _5708_/X VGND VGND VPWR VPWR hold566/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 hold3122/X VGND VGND VPWR VPWR hold3123/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2066 hold542/X VGND VGND VPWR VPWR _5940_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1332 _5604_/X VGND VGND VPWR VPWR _7235_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6119__D _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2077 _5943_/X VGND VGND VPWR VPWR hold111/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2088 hold623/X VGND VGND VPWR VPWR _5611_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1343 _4280_/A1 VGND VGND VPWR VPWR hold2782/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5119_ _5059_/B _5115_/X _5118_/X _5117_/Y VGND VGND VPWR VPWR _5119_/X sky130_fd_sc_hd__a211o_1
Xhold1354 _4302_/A1 VGND VGND VPWR VPWR hold2901/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2099 _6918_/Q VGND VGND VPWR VPWR hold655/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6099_ _6332_/B _6106_/B _6144_/A _6119_/A VGND VGND VPWR VPWR _6099_/X sky130_fd_sc_hd__and4bb_4
XANTENNA__6589__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1365 _4285_/B VGND VGND VPWR VPWR hold2925/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1376 hold1495/X VGND VGND VPWR VPWR hold1496/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1387 hold1744/X VGND VGND VPWR VPWR hold1745/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 _4228_/X VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5549__A1 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6746__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5747__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1864_A _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6210__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4221__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3494__C _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6513__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6277__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5788__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3669__C _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4460__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6737__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6201__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3566__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5960__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5470_ _4605_/Y _5563_/A1 _4971_/X _5265_/A _5469_/Y VGND VGND VPWR VPWR _5564_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_170_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4421_ _4421_/A0 _4420_/X _4423_/S VGND VGND VPWR VPWR _4421_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_151_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3723__B1 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7140_ _7156_/CLK _7140_/D fanout598/X VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_4
X_4352_ _4352_/A _5632_/B _4551_/D VGND VGND VPWR VPWR _4357_/S sky130_fd_sc_hd__and3_2
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6268__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout408 hold1467/X VGND VGND VPWR VPWR _4491_/C sky130_fd_sc_hd__clkbuf_16
X_7071_ _7075_/CLK _7071_/D _6861_/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfstp_4
Xfanout419 _3569_/A VGND VGND VPWR VPWR _5590_/A sky130_fd_sc_hd__buf_12
X_4283_ _4289_/S _4283_/B VGND VGND VPWR VPWR _4283_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4279__A1 _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6022_ _7588_/Q _7589_/Q VGND VGND VPWR VPWR _6022_/X sky130_fd_sc_hd__and2b_4
XANTENNA__3487__C1 _3479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6924_ _6926_/CLK _6924_/D fanout565/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6440__A2 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4451__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6855_ _6871_/A _6872_/B VGND VGND VPWR VPWR _6855_/X sky130_fd_sc_hd__and2_1
XANTENNA__6728__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5806_ _5806_/A0 _5950_/A1 _5811_/S VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6786_ _6792_/S _6786_/B VGND VGND VPWR VPWR _6786_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3998_ _7074_/Q _7073_/Q VGND VGND VPWR VPWR _3998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5737_ _5737_/A0 _5953_/A1 _5739_/S VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5951__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3962__B1 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5668_ _5668_/A _5902_/B VGND VGND VPWR VPWR _5670_/S sky130_fd_sc_hd__nand2_8
XANTENNA__4203__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7407_ _7409_/CLK _7407_/D fanout577/X VGND VGND VPWR VPWR _7407_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_103_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4619_ _4570_/Y _4869_/A2 _4618_/Y VGND VGND VPWR VPWR _4860_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5703__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5599_ _5599_/A0 _5950_/A1 _5602_/S VGND VGND VPWR VPWR _5599_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_142_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold440 hold440/A VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7338_ _7555_/CLK _7338_/D fanout594/X VGND VGND VPWR VPWR _7338_/Q sky130_fd_sc_hd__dfrtp_4
Xhold451 _4338_/X VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold462 hold462/A VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold473 _5616_/X VGND VGND VPWR VPWR _7245_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6259__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold484 hold484/A VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold495 hold495/A VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7269_ _7530_/CLK _7269_/D fanout600/X VGND VGND VPWR VPWR _7269_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6427__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 _4389_/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 hold2809/X VGND VGND VPWR VPWR hold2810/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 hold1162/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
Xhold1173 hold2801/X VGND VGND VPWR VPWR hold2802/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input128_A wb_adr_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 hold1184/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1195 hold2912/X VGND VGND VPWR VPWR hold1195/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5050__B _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4442__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6719__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6195__A1 _7499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6195__B2 _7315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6734__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input93_A trap VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5942__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3953__B1 _3506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5170__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3720__A3 _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6670__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6903__CLK _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5225__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4970_ _5248_/A _5248_/B _5180_/B VGND VGND VPWR VPWR _5052_/A sky130_fd_sc_hd__and3_1
XANTENNA__4433__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3921_ _3897_/X _3904_/X _3921_/C _3921_/D VGND VGND VPWR VPWR _3922_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__3787__A3 _3519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6640_ hold27/A _6424_/C _6771_/A3 _6434_/X _7470_/Q VGND VGND VPWR VPWR _6640_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6186__A1 _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3852_ input37/X _4231_/S _4467_/A _7129_/Q _3851_/X VGND VGND VPWR VPWR _3852_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__6186__B2 _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6571_ _7283_/Q _6431_/Y _6067_/A VGND VGND VPWR VPWR _6571_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3783_ _6914_/Q _5587_/C _5947_/A _3617_/X _7232_/Q VGND VGND VPWR VPWR _3792_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_143_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2462_A _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3944__B1 _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5522_ _4668_/C _4827_/X _5107_/X _5110_/X VGND VGND VPWR VPWR _5559_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6489__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5453_ _5453_/A _5453_/B _5453_/C VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3862__C _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4404_ _4404_/A0 _5951_/A1 _4405_/S VGND VGND VPWR VPWR _4404_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7580_/CLK sky130_fd_sc_hd__clkbuf_16
X_5384_ _5384_/A _5384_/B _5384_/C VGND VGND VPWR VPWR _5390_/A sky130_fd_sc_hd__and3_1
XFILLER_0_100_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5161__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7123_ _7134_/CLK _7123_/D _6833_/A VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_4
X_4335_ _4335_/A0 _5714_/A0 _4339_/S VGND VGND VPWR VPWR _4335_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5850__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7054_ _7170_/CLK _7054_/D fanout573/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfrtp_4
X_4266_ _4266_/A0 _5714_/A0 _4270_/S VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6005_ _7584_/Q _6006_/A VGND VGND VPWR VPWR _6005_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7299_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6661__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4197_ _4197_/A0 _7642_/Q _4429_/B VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__mux2_4
XANTENNA_fanout378_A _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _4127_/A1 _6907_/D _6857_/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3778__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6838_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6838_/X sky130_fd_sc_hd__and2_1
XFILLER_0_49_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6177__A1 _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6177__B2 _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6716__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6769_ _7040_/Q _6459_/B _6651_/C _6421_/X _7010_/Q VGND VGND VPWR VPWR _6769_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3935__B1 hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5688__A0 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3950__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5152__A2 _4758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold270 hold270/A VGND VGND VPWR VPWR _7234_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5045__B _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold281 _3485_/X VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5760__S _5766_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold292 hold292/A VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6652__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5860__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4663__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5061__A _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__A1 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6707__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4179__A0 _6879_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5915__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output297_A _7246_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3926__B1 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5391__A2 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4778__C _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4140__A _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3682__C _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6340__B2 _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4120_ _6882_/Q _7071_/Q _4123_/B _3403_/A VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__a31o_1
Xhold1909 hold366/X VGND VGND VPWR VPWR _5816_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6643__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4051_ _3998_/Y _4062_/A _3403_/A _4051_/B1 VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__a31o_1
XANTENNA__6067__A _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5300__C1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5851__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4953_ _4954_/A _5248_/A _4954_/C VGND VGND VPWR VPWR _4953_/X sky130_fd_sc_hd__and3_4
XFILLER_0_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3904_ _7062_/Q _4394_/A _3899_/X _3901_/X _3903_/X VGND VGND VPWR VPWR _3904_/X
+ sky130_fd_sc_hd__a2111o_1
X_7672_ _7672_/A VGND VGND VPWR VPWR _7672_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4315__A _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4884_ _5213_/B _4884_/B _5213_/C _4937_/C VGND VGND VPWR VPWR _5448_/D sky130_fd_sc_hd__nand4_2
XFILLER_0_46_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6623_ _7285_/Q _6431_/Y _6775_/B1 VGND VGND VPWR VPWR _6623_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_6_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3835_ _7058_/Q hold56/A _5623_/B _3834_/X VGND VGND VPWR VPWR _3835_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_117_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3917__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6554_ _7403_/Q _6409_/X _6549_/X _6553_/X _6430_/X VGND VGND VPWR VPWR _6554_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3766_ _7458_/Q _5785_/B _5866_/B _3537_/X _7426_/Q VGND VGND VPWR VPWR _3766_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5505_ _5342_/A _5094_/A wire536/X _5504_/Y VGND VGND VPWR VPWR _5505_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4135__A_N _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3932__A3 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6485_ _7480_/Q _6451_/X _6480_/X _6482_/X _6484_/X VGND VGND VPWR VPWR _6495_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3697_ _7136_/Q _4473_/A _5619_/B _3661_/X _7035_/Q VGND VGND VPWR VPWR _3697_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5436_ _5339_/D _5339_/C _5425_/X _5170_/X VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput320 hold2783/X VGND VGND VPWR VPWR hold1170/A sky130_fd_sc_hd__buf_6
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput331 hold1211/X VGND VGND VPWR VPWR hold1212/A sky130_fd_sc_hd__buf_6
Xoutput342 hold1199/X VGND VGND VPWR VPWR hold1200/A sky130_fd_sc_hd__buf_6
XANTENNA__4342__A0 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6676__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5367_ _5545_/B _5367_/B _5367_/C _5367_/D VGND VGND VPWR VPWR _5367_/Y sky130_fd_sc_hd__nor4_2
XANTENNA_fanout495_A _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7106_ _7207_/CLK _7106_/D _6780_/B VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4318_ _4321_/S _6789_/A2 _4317_/Y VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__o21ai_2
X_5298_ _4583_/B _4821_/Y _4735_/Y _4687_/Y VGND VGND VPWR VPWR _5298_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6095__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7037_ _7189_/CLK _7037_/D fanout572/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6634__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4249_ _4249_/A0 _4248_/X _4249_/S VGND VGND VPWR VPWR _4249_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6408__C _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4660__A4 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1777_A _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3620__A2 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5373__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6322__A1 _7143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input56_A mgmt_gpio_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3687__A2 _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout580 fanout581/X VGND VGND VPWR VPWR fanout580/X sky130_fd_sc_hd__buf_12
XANTENNA__4636__A1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout591 fanout606/X VGND VGND VPWR VPWR _6833_/A sky130_fd_sc_hd__buf_12
XFILLER_0_189_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3611__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3620_ _5640_/C _5623_/B _3619_/X _3558_/X _7284_/Q VGND VGND VPWR VPWR _3620_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5364__A2 wire533/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3551_ input51/X _4491_/B _5619_/B _5920_/A _7518_/Q VGND VGND VPWR VPWR _3551_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3914__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2258_A _7542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6270_ _7414_/Q _6116_/B _6116_/C _6144_/B VGND VGND VPWR VPWR _6270_/X sky130_fd_sc_hd__o211a_1
X_3482_ _5803_/A _5722_/A _5640_/B VGND VGND VPWR VPWR _5794_/A sky130_fd_sc_hd__and3_4
XANTENNA__4324__A0 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5221_ _5213_/B _5220_/X _5219_/Y VGND VGND VPWR VPWR _5223_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3108 _7551_/Q VGND VGND VPWR VPWR hold3108/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3119 _7423_/Q VGND VGND VPWR VPWR hold3119/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3678__A2 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2407 hold943/X VGND VGND VPWR VPWR _5842_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2418 _7145_/Q VGND VGND VPWR VPWR hold2418/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5152_ _4794_/A _4758_/X _5410_/B _5096_/A wire546/A VGND VGND VPWR VPWR _5153_/C
+ sky130_fd_sc_hd__a32oi_4
XFILLER_0_138_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2429 hold937/X VGND VGND VPWR VPWR _4536_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6077__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4103_ _6462_/D _6435_/B VGND VGND VPWR VPWR _6455_/B sky130_fd_sc_hd__and2b_4
XANTENNA__6616__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1706 hold288/X VGND VGND VPWR VPWR _5762_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1717 _5681_/X VGND VGND VPWR VPWR hold307/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5083_ _5451_/A1 _4720_/Y _4946_/Y _4748_/Y _4717_/Y VGND VGND VPWR VPWR _5083_/X
+ sky130_fd_sc_hd__o32a_1
Xhold1728 _7179_/Q VGND VGND VPWR VPWR hold352/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1739 _7466_/Q VGND VGND VPWR VPWR hold237/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4627__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4034_ _6902_/Q _6901_/Q _6900_/Q _6903_/Q VGND VGND VPWR VPWR _4034_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_78_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3850__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5985_ _5985_/A0 _5985_/A1 _5991_/S VGND VGND VPWR VPWR _5985_/X sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4936_ _4954_/A _4940_/D VGND VGND VPWR VPWR _4936_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3602__A2 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_10 _3921_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7655_ _7655_/A VGND VGND VPWR VPWR _7655_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_21 _7411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4947_/C _4942_/A _4948_/C VGND VGND VPWR VPWR _4933_/B sky130_fd_sc_hd__and3_2
XANTENNA_32 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _4093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _7309_/Q _6420_/B _6425_/X _7341_/Q _6605_/X VGND VGND VPWR VPWR _6606_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_54 _3714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3818_ _7003_/Q _4322_/A _3799_/X _3815_/X _3817_/X VGND VGND VPWR VPWR _3818_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout410_A _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4158__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7586_ _7586_/CLK _7586_/D _4128_/B VGND VGND VPWR VPWR _7586_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_65 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4699__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _5387_/C _4799_/C VGND VGND VPWR VPWR _4798_/Y sky130_fd_sc_hd__nand2_4
X_6537_ _7362_/Q _6462_/X _6468_/X _7410_/Q _6536_/X VGND VGND VPWR VPWR _6544_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3905__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3749_ _7115_/Q _3658_/X _3661_/X _7034_/Q _3748_/X VGND VGND VPWR VPWR _3749_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6468_ _6574_/B _6600_/B _6747_/C VGND VGND VPWR VPWR _6468_/X sky130_fd_sc_hd__and3_4
XFILLER_0_112_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5419_ _5419_/A _5419_/B _5491_/A VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__and3_1
X_6399_ _6961_/Q _6036_/Y _6775_/B1 VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__o21a_1
Xoutput172 _7648_/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
Xoutput183 _3428_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 _3418_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
Xhold2930 hold2930/A VGND VGND VPWR VPWR _4451_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2941 _7065_/Q VGND VGND VPWR VPWR hold700/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2952 _7660_/A VGND VGND VPWR VPWR hold2952/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4618__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2963 hold2963/A VGND VGND VPWR VPWR _4517_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2974 hold2974/A VGND VGND VPWR VPWR _4475_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2985 hold2985/A VGND VGND VPWR VPWR _4184_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2996 _7363_/Q VGND VGND VPWR VPWR hold726/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6083__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5291__A1 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1894_A _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4881__C _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3841__A2 _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input110_A wb_adr_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3497__C _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6543__A1 _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5346__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6543__B2 _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4554__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__B1 _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4609__A1 _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4085__A2 _6879_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5019__D1 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3832__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5770_/A0 _5986_/A1 _5775_/S VGND VGND VPWR VPWR _5770_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6782__A1 _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _5058_/D _4856_/A _5073_/A VGND VGND VPWR VPWR _5059_/B sky130_fd_sc_hd__nor3_4
XFILLER_0_173_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7440_ _7521_/CLK _7440_/D fanout600/X VGND VGND VPWR VPWR _7440_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_56_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4652_ _4648_/A _4591_/Y _5005_/A _4726_/B VGND VGND VPWR VPWR _5222_/C sky130_fd_sc_hd__o211a_4
XANTENNA__6534__A1 _7538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_2
X_3603_ _7445_/Q _3520_/X _5920_/A _7517_/Q _3602_/X VGND VGND VPWR VPWR _3606_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7371_ _7487_/CLK _7371_/D fanout593/X VGND VGND VPWR VPWR _7371_/Q sky130_fd_sc_hd__dfrtp_4
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4583_ _4646_/A _4583_/B VGND VGND VPWR VPWR _4586_/C sky130_fd_sc_hd__nor2_2
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _4174_/A sky130_fd_sc_hd__buf_8
Xhold803 hold803/A VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _4135_/B sky130_fd_sc_hd__clkbuf_4
Xhold814 _5792_/X VGND VGND VPWR VPWR _7397_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6322_ _7143_/Q _6144_/C _6097_/B _6144_/B VGND VGND VPWR VPWR _6322_/X sky130_fd_sc_hd__o211a_1
Xhold825 hold825/A VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3534_ _7534_/Q _3529_/X _5857_/A _7462_/Q _3533_/X VGND VGND VPWR VPWR _3534_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5127__C _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_4
Xmax_cap544 _4704_/Y VGND VGND VPWR VPWR fanout542/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold836 _4405_/X VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap555 _4604_/Y VGND VGND VPWR VPWR _5134_/A sky130_fd_sc_hd__clkbuf_2
Xhold847 hold847/A VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6298__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold858 hold858/A VGND VGND VPWR VPWR hold858/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6253_ _7461_/Q _6112_/C _6079_/X _6094_/X hold76/A VGND VGND VPWR VPWR _6253_/X
+ sky130_fd_sc_hd__a32o_1
Xhold869 hold869/A VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3465_ _4076_/B _4025_/A VGND VGND VPWR VPWR _3465_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_0_149_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4966__C _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5204_ _4605_/Y _4679_/Y _4880_/Y _5203_/Y VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__o31a_1
Xhold2204 _5685_/X VGND VGND VPWR VPWR hold459/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6184_ _7418_/Q _6072_/X _6144_/X _7290_/Q _6183_/X VGND VGND VPWR VPWR _6184_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2215 hold891/X VGND VGND VPWR VPWR _5719_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2226 _5787_/X VGND VGND VPWR VPWR hold531/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2237 hold454/X VGND VGND VPWR VPWR _5802_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5135_ _4790_/B _5077_/B _5297_/B _5138_/D VGND VGND VPWR VPWR _5135_/Y sky130_fd_sc_hd__a22oi_2
Xhold1503 _7500_/Q VGND VGND VPWR VPWR hold225/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2248 hold610/X VGND VGND VPWR VPWR _5793_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2259 hold534/X VGND VGND VPWR VPWR _5955_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1514 _5980_/X VGND VGND VPWR VPWR hold210/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1525 hold204/X VGND VGND VPWR VPWR _7281_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1536 hold30/X VGND VGND VPWR VPWR _7438_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_165_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1547 _5998_/X VGND VGND VPWR VPWR hold208/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1558 _4434_/X VGND VGND VPWR VPWR hold196/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5066_ _5096_/A _5453_/C VGND VGND VPWR VPWR _5444_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_74_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1569 hold220/X VGND VGND VPWR VPWR _7452_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6470__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4017_ hold51/A _4017_/B VGND VGND VPWR VPWR _4017_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3598__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6758__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6222__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6405__D _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5968_ _5968_/A0 _5995_/A1 hold13/X VGND VGND VPWR VPWR _5968_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_177_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4233__C1 hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4919_ _4919_/A _5573_/C _4919_/C VGND VGND VPWR VPWR _4922_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_164_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5899_ _5998_/A1 hold187/X _5901_/S VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6702__B _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7638_ _7646_/CLK _7638_/D _4309_/B VGND VGND VPWR VPWR _7638_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6525__A1 _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6525__B2 _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6421__C _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4536__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7569_ _7569_/CLK _7569_/D fanout597/X VGND VGND VPWR VPWR _7569_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_132_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6828__A2 _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input158_A wb_dat_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5053__B _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3023_A _7025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2760 _7151_/Q VGND VGND VPWR VPWR hold858/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2771 hold2771/A VGND VGND VPWR VPWR _4272_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2782 hold2782/A VGND VGND VPWR VPWR hold2782/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4892__B _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2793 hold2793/A VGND VGND VPWR VPWR _4534_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input19_A mask_rev_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3814__A2 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5016__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6213__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6764__A1 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3750__A1 _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3463__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5255__A1 _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6940_ _6956_/CLK _6940_/D fanout604/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3805__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ _6871_/A _6872_/B VGND VGND VPWR VPWR _6871_/X sky130_fd_sc_hd__and2_1
XFILLER_0_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6204__B1 _6106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5822_ _5822_/A0 _5993_/A1 _5829_/S VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_151_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5753_ _5753_/A0 _5951_/A1 _5757_/S VGND VGND VPWR VPWR _5753_/X sky130_fd_sc_hd__mux2_1
X_4704_ _4825_/A _5071_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _4704_/Y sky130_fd_sc_hd__nor4_4
XANTENNA__3865__C _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5684_ _5684_/A0 _5954_/A1 _5685_/S VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7423_ _7471_/CLK _7423_/D fanout593/X VGND VGND VPWR VPWR _7423_/Q sky130_fd_sc_hd__dfstp_1
X_4635_ _4856_/A _4574_/X _4733_/B VGND VGND VPWR VPWR _4730_/C sky130_fd_sc_hd__a21boi_4
XANTENNA__5853__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold600 hold600/A VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7354_ _7575_/CLK _7354_/D fanout595/X VGND VGND VPWR VPWR _7354_/Q sky130_fd_sc_hd__dfrtp_4
X_4566_ _4772_/A _4805_/B VGND VGND VPWR VPWR _5100_/A sky130_fd_sc_hd__and2_4
Xhold611 _5793_/X VGND VGND VPWR VPWR _7398_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold622 hold622/A VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold633 hold633/A VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold644 _5912_/X VGND VGND VPWR VPWR _7503_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap352 _5653_/S VGND VGND VPWR VPWR _5656_/S sky130_fd_sc_hd__clkbuf_2
X_6305_ _6957_/Q _6036_/Y _6775_/B1 VGND VGND VPWR VPWR _6305_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_13_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3741__A1 _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3517_ _7242_/Q _3515_/X hold72/A _7566_/Q _3513_/X VGND VGND VPWR VPWR _3524_/C
+ sky130_fd_sc_hd__a221o_1
Xmax_cap363 _4836_/A VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__clkbuf_2
Xhold655 hold655/A VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7285_ _7299_/CLK _7285_/D fanout579/X VGND VGND VPWR VPWR _7285_/Q sky130_fd_sc_hd__dfrtp_4
Xhold666 hold666/A VGND VGND VPWR VPWR hold666/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4497_ _4497_/A _4551_/D VGND VGND VPWR VPWR _4502_/S sky130_fd_sc_hd__nand2_4
Xhold677 hold677/A VGND VGND VPWR VPWR _7223_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold688 hold688/A VGND VGND VPWR VPWR hold688/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6236_ _6224_/X _6234_/X _6235_/X VGND VGND VPWR VPWR _6236_/X sky130_fd_sc_hd__o21a_1
Xhold699 _4345_/X VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3448_ _4028_/A0 _6904_/Q _4025_/A VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6286__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2001 _5834_/X VGND VGND VPWR VPWR hold441/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2012 _6921_/Q VGND VGND VPWR VPWR hold494/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4297__A2 _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6691__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5494__B2 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2023 _7130_/Q VGND VGND VPWR VPWR hold510/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2034 hold486/X VGND VGND VPWR VPWR _4459_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6161_/X _6163_/X _6164_/X _6166_/X VGND VGND VPWR VPWR _6167_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4993__A _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 hold3028/X VGND VGND VPWR VPWR hold3029/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout575_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2045 _7115_/Q VGND VGND VPWR VPWR hold482/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 hold3162/X VGND VGND VPWR VPWR hold3163/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2056 _7150_/Q VGND VGND VPWR VPWR hold508/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1322 hold3124/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5118_/A _5118_/B _5118_/C VGND VGND VPWR VPWR _5118_/X sky130_fd_sc_hd__and3_1
Xhold2067 _5940_/X VGND VGND VPWR VPWR _7528_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1333 hold3128/X VGND VGND VPWR VPWR hold3129/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2078 _7259_/Q VGND VGND VPWR VPWR hold108/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2089 _5611_/X VGND VGND VPWR VPWR _7242_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1344 _4313_/B VGND VGND VPWR VPWR hold2787/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6098_ _7407_/Q _6097_/B _6144_/B _6097_/X _7439_/Q VGND VGND VPWR VPWR _6098_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1355 _4291_/B VGND VGND VPWR VPWR hold2877/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1366 _6788_/B VGND VGND VPWR VPWR hold3081/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1377 _7188_/Q VGND VGND VPWR VPWR _4541_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
X_5049_ _5339_/D _5342_/A _5260_/D _5339_/C VGND VGND VPWR VPWR _5051_/C sky130_fd_sc_hd__nand4_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1388 hold2146/X VGND VGND VPWR VPWR hold2147/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1399 hold91/X VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6416__C _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5549__A2 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5763__S _5766_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4887__B _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6131__C1 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3280 _6901_/Q VGND VGND VPWR VPWR _4041_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2590 _5823_/X VGND VGND VPWR VPWR hold713/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3799__A1 _7441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6737__A1 _6991_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6737__B2 _7034_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6201__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4420_ _4447_/A0 hold61/X _4422_/S VGND VGND VPWR VPWR _4420_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4797__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3723__A1 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4351_ _4351_/A0 _5754_/A1 _4351_/S VGND VGND VPWR VPWR _4351_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3723__B2 _7339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4289__S _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7070_ _7070_/CLK _7070_/D fanout590/X VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout409 _4455_/C VGND VGND VPWR VPWR _4388_/B sky130_fd_sc_hd__buf_12
X_4282_ _4289_/S _3856_/B _4281_/Y VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__4279__A2 _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6021_ _7589_/Q _7588_/Q VGND VGND VPWR VPWR _6072_/B sky130_fd_sc_hd__and2b_4
XFILLER_0_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6923_ _6926_/CLK _6923_/D fanout565/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__7489__RESET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6854_ _6871_/A _6872_/B VGND VGND VPWR VPWR _6854_/X sky130_fd_sc_hd__and2_1
XANTENNA__6728__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5805_ _5805_/A0 _5805_/A1 _5811_/S VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6785_ _6792_/S _3856_/B _6784_/Y VGND VGND VPWR VPWR _7631_/D sky130_fd_sc_hd__o21ai_1
X_3997_ _3997_/A1 _3996_/A _3996_/Y _3923_/S VGND VGND VPWR VPWR _7214_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_18_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5736_ _5736_/A0 hold84/X _5739_/S VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__mux2_1
XFILLER_0_134_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5667_ _5667_/A0 _5955_/A1 _5667_/S VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3962__B2 _7399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4203__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4618_ _4667_/A _4869_/A2 _4795_/C VGND VGND VPWR VPWR _4618_/Y sky130_fd_sc_hd__o21bai_4
X_7406_ _7501_/CLK _7406_/D fanout581/X VGND VGND VPWR VPWR _7406_/Q sky130_fd_sc_hd__dfrtp_4
X_5598_ _5598_/A0 _5805_/A1 _5602_/S VGND VGND VPWR VPWR _5598_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7337_ _7539_/CLK _7337_/D fanout578/X VGND VGND VPWR VPWR _7337_/Q sky130_fd_sc_hd__dfrtp_4
Xhold430 hold430/A VGND VGND VPWR VPWR hold430/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4549_ _5951_/A1 _4549_/A1 _4550_/S VGND VGND VPWR VPWR _4549_/X sky130_fd_sc_hd__mux2_1
Xhold441 hold441/A VGND VGND VPWR VPWR _7434_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold452 hold452/A VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold463 hold463/A VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold474 hold474/A VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7268_ _7268_/CLK _7268_/D _6871_/A VGND VGND VPWR VPWR _7268_/Q sky130_fd_sc_hd__dfrtp_1
Xhold485 _5703_/X VGND VGND VPWR VPWR _7318_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold496 hold496/A VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6219_ _7516_/Q _6332_/B _6317_/C _6072_/X _7420_/Q VGND VGND VPWR VPWR _6219_/X
+ sky130_fd_sc_hd__a32o_1
X_7199_ _7201_/CLK _7199_/D _6839_/A VGND VGND VPWR VPWR _7199_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5612__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 _4475_/X VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 hold3021/X VGND VGND VPWR VPWR hold3022/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 hold1152/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 hold2806/X VGND VGND VPWR VPWR hold2807/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1174 hold1174/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
Xhold1185 hold2883/X VGND VGND VPWR VPWR hold1185/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1196 hold1196/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6719__A1 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5059__A _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input86_A spimemio_flash_io0_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3953__A1 _7132_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5458__A1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6655__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4969__B1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5630__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3920_ _7520_/Q _5929_/A _5634_/A _7260_/Q _3919_/X VGND VGND VPWR VPWR _3921_/D
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3851_ _7545_/Q _4491_/B _4212_/A _5643_/A _4174_/A VGND VGND VPWR VPWR _3851_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6186__A2 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6072__B _6072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2288_A _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6570_ _6554_/X _6570_/B _6570_/C VGND VGND VPWR VPWR _6570_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_143_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3782_ _3782_/A _3782_/B _3782_/C _3782_/D VGND VGND VPWR VPWR _3793_/C sky130_fd_sc_hd__nor4_1
XFILLER_0_128_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5521_ _5521_/A _5521_/B _5562_/C _5521_/D VGND VGND VPWR VPWR _5521_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__3944__A1 _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5452_ _5510_/B _5452_/B _5574_/A VGND VGND VPWR VPWR _5456_/C sky130_fd_sc_hd__and3_1
XFILLER_0_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5697__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4403_ _4403_/A0 _5815_/A1 _4405_/S VGND VGND VPWR VPWR _4403_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5383_ _5077_/Y _5255_/X _5378_/X _5380_/X _5382_/X VGND VGND VPWR VPWR _5384_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_100_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7122_ _7134_/CLK _7122_/D _6833_/A VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4334_ _4551_/A _4551_/C _4352_/A hold47/X VGND VGND VPWR VPWR _4339_/S sky130_fd_sc_hd__and4_4
XANTENNA__5449__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7053_ _7211_/CLK _7053_/D fanout572/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_10_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4265_ _5632_/B _5659_/B _4551_/D VGND VGND VPWR VPWR _4270_/S sky130_fd_sc_hd__and3_4
X_6004_ _6751_/S _4107_/A _6932_/Q _6006_/A VGND VGND VPWR VPWR _6018_/A sky130_fd_sc_hd__a211o_1
X_4196_ _4196_/A0 _5754_/A1 _4202_/S VGND VGND VPWR VPWR _4196_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2991_A _7352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4990__B _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5621__A1 hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6906_ _4127_/A1 _6906_/D _6856_/X VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6837_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6837_/X sky130_fd_sc_hd__and2_1
XFILLER_0_18_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6177__A2 _6116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4188__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6768_ _7045_/Q _6408_/B _6425_/X _7020_/Q _6767_/X VGND VGND VPWR VPWR _6773_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5719_ _5953_/A1 _5719_/A1 _5721_/S VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3935__B2 _7559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6699_ _6958_/Q _6431_/Y _6775_/B1 VGND VGND VPWR VPWR _6699_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5137__B1 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6334__C1 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3699__B1 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold260 hold260/A VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4360__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold271 hold271/A VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold282 _5587_/C VGND VGND VPWR VPWR _5619_/A sky130_fd_sc_hd__buf_2
Xhold293 hold293/A VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6101__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5342__A _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input140_A wb_dat_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3926__A1 _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5391__A3 _4744_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_user_clock_A user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5679__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6340__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4351__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6628__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4050_ _4050_/A0 _3400_/A _4050_/S VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__mux2_1
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_189_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4406__A2 hold284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4952_ _5222_/A _4952_/B VGND VGND VPWR VPWR _4958_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3614__B1 hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3903_ _7448_/Q _5848_/A _3520_/X _7440_/Q _3902_/X VGND VGND VPWR VPWR _3903_/X
+ sky130_fd_sc_hd__a221o_1
X_7671_ _7671_/A VGND VGND VPWR VPWR _7671_/X sky130_fd_sc_hd__clkbuf_2
X_4883_ _5180_/A _5216_/A _5342_/B VGND VGND VPWR VPWR _4904_/A sky130_fd_sc_hd__and3_2
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6622_ _7293_/Q _6422_/X _6604_/X _6615_/X _6621_/X VGND VGND VPWR VPWR _6622_/X
+ sky130_fd_sc_hd__a2111o_2
X_3834_ _7053_/Q _4509_/A _5619_/B _3544_/X _7417_/Q VGND VGND VPWR VPWR _3834_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_171_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6553_ _7531_/Q _6058_/X _6551_/X _6552_/X VGND VGND VPWR VPWR _6553_/X sky130_fd_sc_hd__a211o_1
X_3765_ _7160_/Q hold56/A _5632_/B _4394_/A _7064_/Q VGND VGND VPWR VPWR _3765_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5382__A3 _4971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5504_ _5572_/A _5504_/B _5550_/A _5550_/B VGND VGND VPWR VPWR _5504_/Y sky130_fd_sc_hd__nand4_1
X_6484_ _7304_/Q _6420_/B _6454_/X _7488_/Q _6483_/X VGND VGND VPWR VPWR _6484_/X
+ sky130_fd_sc_hd__a221o_1
X_3696_ _7196_/Q _4545_/A _3690_/X _3691_/X _3695_/X VGND VGND VPWR VPWR _3733_/C
+ sky130_fd_sc_hd__a2111oi_1
Xpad_flashh_clk_buff_inst _4127_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_8
X_5435_ _5499_/A _5435_/B _5501_/A _5435_/D VGND VGND VPWR VPWR _5438_/A sky130_fd_sc_hd__nor4_1
Xoutput310 _7673_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 hold2791/X VGND VGND VPWR VPWR hold1176/A sky130_fd_sc_hd__buf_6
XANTENNA__5861__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput332 hold1215/X VGND VGND VPWR VPWR hold1216/A sky130_fd_sc_hd__buf_6
XFILLER_0_168_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput343 hold2802/X VGND VGND VPWR VPWR hold1174/A sky130_fd_sc_hd__buf_6
X_5366_ _5248_/B _5453_/A _5243_/C _5367_/D VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4985__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6619__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7105_ _7644_/CLK _7105_/D _4309_/B VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_2
X_4317_ _4321_/S _4317_/B VGND VGND VPWR VPWR _4317_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout390_A hold2225/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5297_ _5297_/A _5297_/B VGND VGND VPWR VPWR _5297_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout488_A _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6095__A1 _7487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7036_ _7144_/CLK _7036_/D fanout572/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6095__B2 _7503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4248_ _5658_/A1 _5955_/A1 _4248_/S VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5842__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6408__D _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7433__RESET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4179_ _6879_/Q _4179_/A1 _4429_/B VGND VGND VPWR VPWR _4179_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_41_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_179_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3605__B1 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__C _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3620__A3 _3619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4879__C _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6322__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5771__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold3053_A _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4333__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3687__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input49_A mgmt_gpio_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5072__A _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout570 _6871_/A VGND VGND VPWR VPWR _6873_/A sky130_fd_sc_hd__buf_6
Xfanout581 fanout582/X VGND VGND VPWR VPWR fanout581/X sky130_fd_sc_hd__buf_12
XANTENNA__5833__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout592 fanout606/X VGND VGND VPWR VPWR _6839_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_189_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7103__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6389__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7555_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4135__B _4135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7542_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6561__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5364__A3 _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3550_ _4551_/A hold22/A _5938_/C VGND VGND VPWR VPWR _5920_/A sky130_fd_sc_hd__and3_4
XANTENNA__6777__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3481_ _5722_/A _5938_/B VGND VGND VPWR VPWR _3481_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6313__A2 _6072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5220_ _5213_/A _5213_/C _5342_/B _5248_/C _5077_/B VGND VGND VPWR VPWR _5220_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3109 hold3109/A VGND VGND VPWR VPWR _5966_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_121_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3678__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5151_ _5563_/A1 _4722_/Y _4787_/Y _4821_/Y _4783_/Y VGND VGND VPWR VPWR _5153_/B
+ sky130_fd_sc_hd__o32a_1
Xhold2408 _5842_/X VGND VGND VPWR VPWR hold944/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2419 hold2419/A VGND VGND VPWR VPWR _4489_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6077__A1 _7343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4102_ _7597_/Q _7598_/Q VGND VGND VPWR VPWR _6427_/A sky130_fd_sc_hd__and2b_4
XANTENNA_hold2418_A _7145_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1707 _5762_/X VGND VGND VPWR VPWR hold289/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_138_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5082_ _4717_/Y _4748_/Y _4946_/Y _4727_/Y _5081_/Y VGND VGND VPWR VPWR _5084_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__6616__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1718 _7578_/Q VGND VGND VPWR VPWR hold277/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1729 hold352/X VGND VGND VPWR VPWR _4530_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5824__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4033_ _4033_/A0 _4032_/X _4040_/A VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4872__A_N _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5984_ _5984_/A0 _5993_/A1 _5991_/S VGND VGND VPWR VPWR _5984_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4935_ _4954_/A _5453_/A _4940_/D VGND VGND VPWR VPWR _4935_/X sky130_fd_sc_hd__and3_1
XFILLER_0_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7267_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__5856__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3602__A3 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 _3961_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7654_ _7654_/A VGND VGND VPWR VPWR _7654_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_22 _7411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _5183_/C _4929_/A _5180_/A VGND VGND VPWR VPWR _4927_/A sky130_fd_sc_hd__and3_1
XFILLER_0_62_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_33 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_44 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ _7493_/Q _6463_/A _6441_/X _6409_/X _7405_/Q VGND VGND VPWR VPWR _6605_/X
+ sky130_fd_sc_hd__a32o_1
X_3817_ _7281_/Q _3558_/X _3659_/X _7008_/Q _3816_/X VGND VGND VPWR VPWR _3817_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_55 _3961_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4797_ _5260_/A _4797_/B _5260_/C VGND VGND VPWR VPWR _4797_/X sky130_fd_sc_hd__and3_1
XANTENNA__4158__A4 _6881_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7585_ _7601_/CLK _7585_/D _4128_/B VGND VGND VPWR VPWR _7585_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_66 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6552__A2 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4699__C _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5760__A0 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _7466_/Q _6434_/B _6574_/C _6446_/X _7522_/Q VGND VGND VPWR VPWR _6536_/X
+ sky130_fd_sc_hd__a32o_1
X_3748_ _7354_/Q _3506_/X _5776_/A _7386_/Q _3738_/X VGND VGND VPWR VPWR _3748_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_15_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3679_ _7191_/Q _4551_/A _4551_/C hold56/A _3678_/X VGND VGND VPWR VPWR _3679_/X
+ sky130_fd_sc_hd__a41o_1
X_6467_ _6467_/A _6600_/B _6747_/C VGND VGND VPWR VPWR _6467_/X sky130_fd_sc_hd__and3_4
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5418_ _5532_/A _5531_/D _5531_/A VGND VGND VPWR VPWR _5491_/A sky130_fd_sc_hd__and3_1
X_6398_ _6383_/X _6385_/X _6397_/Y VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__a21bo_4
XFILLER_0_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput173 _4176_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
Xoutput184 _3427_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
X_5349_ _5349_/A _5349_/B VGND VGND VPWR VPWR _5355_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_11_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput195 _3417_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XANTENNA__6068__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3405__A _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6419__C _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2920 hold2920/A VGND VGND VPWR VPWR _5985_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2931 _7376_/Q VGND VGND VPWR VPWR hold2931/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6607__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2942 hold700/X VGND VGND VPWR VPWR _4399_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2953 hold2953/A VGND VGND VPWR VPWR _4417_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5815__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2964 _7367_/Q VGND VGND VPWR VPWR hold2964/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2975 _7193_/Q VGND VGND VPWR VPWR hold2975/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7019_ _7170_/CLK _7019_/D fanout573/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2986 _4184_/X VGND VGND VPWR VPWR hold2986/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2997 hold726/X VGND VGND VPWR VPWR _5754_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_168_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3841__A3 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input103_A wb_adr_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5766__S _5766_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6543__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4306__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4609__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5806__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4490__A0 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5019__C1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3832__A3 _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6231__B2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6782__A2 _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3596__A2 _3543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _4836_/C _5079_/B VGND VGND VPWR VPWR _4720_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4651_ _4591_/Y _4648_/A _4726_/B VGND VGND VPWR VPWR _4948_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__6080__B _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6534__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR _3930_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3602_ _7241_/Q _5612_/B _5603_/B _5686_/A _7309_/Q VGND VGND VPWR VPWR _3602_/X
+ sky130_fd_sc_hd__a32o_4
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_9_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4582_ _4887_/D _4747_/B _4887_/B _4879_/C VGND VGND VPWR VPWR _4583_/B sky130_fd_sc_hd__nand4_4
X_7370_ _7575_/CLK _7370_/D fanout595/X VGND VGND VPWR VPWR _7370_/Q sky130_fd_sc_hd__dfrtp_4
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__buf_2
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_2
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold804 hold804/A VGND VGND VPWR VPWR _7557_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3533_ input60/X _5785_/B _5965_/A _3531_/X _7342_/Q VGND VGND VPWR VPWR _3533_/X
+ sky130_fd_sc_hd__a32o_1
X_6321_ _7022_/Q _6070_/X _6110_/X _7173_/Q _6320_/X VGND VGND VPWR VPWR _6327_/B
+ sky130_fd_sc_hd__a221o_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _4129_/B sky130_fd_sc_hd__buf_4
Xhold815 hold815/A VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold826 hold826/A VGND VGND VPWR VPWR _7081_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap534 _4856_/Y VGND VGND VPWR VPWR _5199_/C sky130_fd_sc_hd__clkbuf_4
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__clkbuf_2
Xmax_cap545 _4704_/Y VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold837 hold837/A VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap556 _4748_/C VGND VGND VPWR VPWR _5091_/A sky130_fd_sc_hd__buf_12
Xhold848 hold848/A VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6252_ _7413_/Q _6116_/B _6116_/C _6144_/B VGND VGND VPWR VPWR _6252_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6298__B2 _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3464_ hold34/X _3505_/C VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__and2b_1
Xhold859 _4496_/X VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5203_ _5342_/A _5203_/B _5295_/C _5339_/D VGND VGND VPWR VPWR _5203_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_0_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7096__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6183_ _7386_/Q _6109_/X _6110_/X _7434_/Q _6182_/X VGND VGND VPWR VPWR _6183_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2205 _6917_/Q VGND VGND VPWR VPWR hold878/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2216 _7503_/Q VGND VGND VPWR VPWR hold643/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5134_ _5134_/A _5260_/C _5134_/C VGND VGND VPWR VPWR _5134_/X sky130_fd_sc_hd__and3_1
Xhold2227 hold531/X VGND VGND VPWR VPWR _7392_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2238 _5802_/X VGND VGND VPWR VPWR hold455/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2249 _7245_/Q VGND VGND VPWR VPWR hold472/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1504 hold225/X VGND VGND VPWR VPWR _5908_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1515 _7513_/Q VGND VGND VPWR VPWR hold183/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1526 _7558_/Q VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1537 _7545_/Q VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5065_ _5213_/B _5453_/C VGND VGND VPWR VPWR _5065_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__3808__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1548 _7428_/Q VGND VGND VPWR VPWR hold271/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1559 _7258_/Q VGND VGND VPWR VPWR hold223/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_74_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4016_ _6905_/Q _6904_/Q _4025_/B VGND VGND VPWR VPWR _4017_/B sky130_fd_sc_hd__and3_1
XANTENNA__6470__A1 _7503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5273__A2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3598__C _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6222__B2 _7508_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5967_ _5967_/A0 _5967_/A1 hold13/X VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4233__B1 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5981__A0 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4918_ _5213_/A _4932_/B _4929_/A _5342_/B VGND VGND VPWR VPWR _4919_/C sky130_fd_sc_hd__nand4_1
XANTENNA_fanout618_A _4945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6702__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5898_ _5979_/A0 hold96/X _5901_/S VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__mux2_1
X_7637_ _7646_/CLK _7637_/D _4309_/B VGND VGND VPWR VPWR _7637_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4503__B _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6525__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4849_ _5342_/A _4849_/B _5138_/D VGND VGND VPWR VPWR _4849_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4768__A_N _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1468_A _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7568_ _7580_/CLK _7568_/D fanout596/X VGND VGND VPWR VPWR _7568_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6519_ _7457_/Q _6455_/X _6463_/X _7425_/Q _6518_/X VGND VGND VPWR VPWR _6519_/X
+ sky130_fd_sc_hd__a221o_1
X_7499_ _7499_/CLK _7499_/D fanout578/X VGND VGND VPWR VPWR _7499_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6289__A1 _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2750 _5651_/X VGND VGND VPWR VPWR hold2750/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2761 hold858/X VGND VGND VPWR VPWR _4496_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2772 _7132_/Q VGND VGND VPWR VPWR hold2772/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2783 hold2783/A VGND VGND VPWR VPWR hold2783/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2794 _4534_/X VGND VGND VPWR VPWR hold2794/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4472__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3814__A3 _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6213__A1 _7283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6764__A2 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6516__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3750__A2 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4786__D _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3443__2 _3443__2/A VGND VGND VPWR VPWR _6823_/A3 sky130_fd_sc_hd__inv_2
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5255__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6075__B _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3805__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6790__S _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6870_ _6871_/A _6872_/B VGND VGND VPWR VPWR _6870_/X sky130_fd_sc_hd__and2_1
XFILLER_0_135_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6204__A1 _7363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5821_ _5866_/B hold12/X hold48/A VGND VGND VPWR VPWR _5829_/S sky130_fd_sc_hd__and3_4
XANTENNA__6755__A2 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4215__B1 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4604__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5752_ _5752_/A0 _5950_/A1 _5757_/S VGND VGND VPWR VPWR _5752_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4910__A_N _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4703_ _5399_/B _5072_/B VGND VGND VPWR VPWR _4703_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3865__D _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5683_ _5683_/A0 _5953_/A1 _5685_/S VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6507__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5715__A0 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7422_ _7478_/CLK _7422_/D fanout583/X VGND VGND VPWR VPWR _7422_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4518__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4634_ _4743_/A _4856_/A _4888_/B _5282_/A _4805_/B VGND VGND VPWR VPWR _4733_/B
+ sky130_fd_sc_hd__a41o_4
XANTENNA__7267__CLK _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3726__C1 _3725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4565_ _4565_/A _4565_/B VGND VGND VPWR VPWR _4675_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_25_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold601 hold601/A VGND VGND VPWR VPWR _7422_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7353_ _7478_/CLK _7353_/D fanout583/X VGND VGND VPWR VPWR _7353_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5191__A1 _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold612 hold612/A VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4977__C _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold623 hold623/A VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold634 hold634/A VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6304_ _6289_/X _6291_/X _6303_/Y VGND VGND VPWR VPWR _6304_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold645 hold645/A VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7206__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3741__A2 _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3516_ hold22/A _5830_/C _5992_/C VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__and3_4
X_7284_ _7309_/CLK _7284_/D fanout579/X VGND VGND VPWR VPWR _7284_/Q sky130_fd_sc_hd__dfrtp_4
Xhold656 hold656/A VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4496_ _4496_/A0 _5586_/A0 _4496_/S VGND VGND VPWR VPWR _4496_/X sky130_fd_sc_hd__mux2_1
Xhold667 _4348_/X VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold678 hold678/A VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6235_ _7284_/Q _6036_/Y _6775_/B1 VGND VGND VPWR VPWR _6235_/X sky130_fd_sc_hd__o21a_1
X_3447_ _6904_/Q _4025_/A VGND VGND VPWR VPWR _3447_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6140__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold689 hold689/A VGND VGND VPWR VPWR _7555_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2002 _7099_/Q VGND VGND VPWR VPWR hold135/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_176_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2013 hold494/X VGND VGND VPWR VPWR _4206_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5494__A2 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2024 hold510/X VGND VGND VPWR VPWR _4471_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2035 _4459_/X VGND VGND VPWR VPWR hold487/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6166_ _7345_/Q _6070_/X _6072_/X _7417_/Q _6165_/X VGND VGND VPWR VPWR _6166_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 hold3030/X VGND VGND VPWR VPWR _7224_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2046 hold482/X VGND VGND VPWR VPWR _4453_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 _5948_/X VGND VGND VPWR VPWR _7535_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2057 hold508/X VGND VGND VPWR VPWR _4495_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2068 _6886_/Q VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 hold3170/X VGND VGND VPWR VPWR hold3171/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5117_ _4826_/Y _4832_/Y _5528_/A3 _5116_/X _5112_/X VGND VGND VPWR VPWR _5117_/Y
+ sky130_fd_sc_hd__o311ai_4
Xhold1334 _4486_/X VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6097_ _6110_/A _6097_/B _6120_/B VGND VGND VPWR VPWR _6097_/X sky130_fd_sc_hd__and3_4
Xhold2079 hold108/X VGND VGND VPWR VPWR _5636_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1345 _4301_/A1 VGND VGND VPWR VPWR hold2883/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout568_A fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5246__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1356 _6792_/A1 VGND VGND VPWR VPWR hold2861/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5048_ _5339_/D _5339_/A _5203_/B _5260_/D VGND VGND VPWR VPWR _5051_/B sky130_fd_sc_hd__nand4_1
Xhold1367 _6954_/Q VGND VGND VPWR VPWR _4256_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1378 hold1768/X VGND VGND VPWR VPWR hold1769/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1389 _7392_/Q VGND VGND VPWR VPWR _5787_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6999_ _6999_/CLK _6999_/D VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6746__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5706__A0 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4887__C _4945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input170_A wb_we_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6131__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3270 _7584_/Q VGND VGND VPWR VPWR _4099_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input31_A mask_rev_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3281 _6895_/Q VGND VGND VPWR VPWR _4053_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2580 hold805/X VGND VGND VPWR VPWR _5837_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2591 _7311_/Q VGND VGND VPWR VPWR hold2591/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1890 _4254_/X VGND VGND VPWR VPWR hold405/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_81_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3799__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6198__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6737__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5173__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6370__B1 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5173__B2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4350_ _4350_/A0 _5647_/A0 _4351_/S VGND VGND VPWR VPWR _4350_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3723__A2 _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4281_ _4289_/S _4281_/B VGND VGND VPWR VPWR _4281_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_190_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6673__A1 _7182_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6020_ _6051_/C _6019_/Y _6020_/S VGND VGND VPWR VPWR _7588_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3487__A1 _7406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3503__A _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6922_ _7255_/CLK _6922_/D fanout565/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_89_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6853_ _6871_/A _6872_/B VGND VGND VPWR VPWR _6853_/X sky130_fd_sc_hd__and2_1
XANTENNA__6728__A2 _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5804_ _5804_/A0 _5948_/A1 _5811_/S VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5936__A0 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4334__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6784_ _6792_/S _6784_/B VGND VGND VPWR VPWR _6784_/Y sky130_fd_sc_hd__nand2_1
X_3996_ _3996_/A _3996_/B VGND VGND VPWR VPWR _3996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5735_ _5735_/A0 _5735_/A1 _5739_/S VGND VGND VPWR VPWR _5735_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7458__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5864__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3962__A2 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5666_ _5666_/A0 _5954_/A1 _5667_/S VGND VGND VPWR VPWR _5666_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_1_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7405_ _7577_/CLK _7405_/D fanout584/X VGND VGND VPWR VPWR _7405_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4617_ _4570_/Y _4869_/A2 _4740_/D VGND VGND VPWR VPWR _4617_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6361__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5597_ _5597_/A0 _5948_/A1 _5602_/S VGND VGND VPWR VPWR _5597_/X sky130_fd_sc_hd__mux2_1
Xhold420 hold420/A VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7336_ _7412_/CLK _7336_/D fanout580/X VGND VGND VPWR VPWR _7336_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__3714__A2 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold431 hold431/A VGND VGND VPWR VPWR _7426_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4548_ _5815_/A1 _4548_/A1 _4550_/S VGND VGND VPWR VPWR _4548_/X sky130_fd_sc_hd__mux2_1
Xhold442 hold442/A VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold453 hold453/A VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold464 hold464/A VGND VGND VPWR VPWR hold464/X sky130_fd_sc_hd__buf_12
XANTENNA__6113__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold475 _5885_/X VGND VGND VPWR VPWR _7479_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7267_ _7267_/CLK _7267_/D fanout605/X VGND VGND VPWR VPWR _7670_/A sky130_fd_sc_hd__dfrtp_1
Xhold486 hold486/A VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4479_ _4491_/B _4521_/B _4551_/D VGND VGND VPWR VPWR _4484_/S sky130_fd_sc_hd__and3_2
XFILLER_0_187_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold497 hold497/A VGND VGND VPWR VPWR _7374_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6664__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6218_ _7412_/Q _6121_/C _6116_/C _6136_/C VGND VGND VPWR VPWR _6218_/X sky130_fd_sc_hd__o211a_1
X_7198_ _7201_/CLK _7198_/D _6839_/A VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5612__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1120 _5913_/X VGND VGND VPWR VPWR _7504_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _7529_/Q _6092_/X _6120_/X _7337_/Q _6148_/X VGND VGND VPWR VPWR _6149_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4509__A _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3413__A _7538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6427__C _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1131 hold3019/X VGND VGND VPWR VPWR hold3020/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 _4378_/X VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 hold2763/X VGND VGND VPWR VPWR hold2764/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 hold1164/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
Xhold1175 hold2790/X VGND VGND VPWR VPWR hold2791/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 hold1186/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
Xhold1197 hold2916/X VGND VGND VPWR VPWR hold1197/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6443__B _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6719__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5927__A0 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6195__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5774__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3953__A2 _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5155__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input79_A spi_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold3250_A _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6104__B1 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5803__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output235_A _4147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3641__B2 _6916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3850_ input22/X _3488_/X _3542_/X _6921_/Q VGND VGND VPWR VPWR _3850_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6072__C _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3781_ _7410_/Q _5803_/A _3590_/C _3780_/X VGND VGND VPWR VPWR _3782_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6591__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5520_ _5521_/A _5521_/B _5521_/D VGND VGND VPWR VPWR _5520_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_171_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5451_ _5451_/A1 _4720_/Y _4844_/Y _5448_/D _5223_/C VGND VGND VPWR VPWR _5508_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4601__B _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2350_A _7283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4402_ _4402_/A0 _5583_/A0 _4405_/S VGND VGND VPWR VPWR _4402_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_151_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5382_ _4605_/Y _5563_/A1 _4971_/X _5265_/A _5381_/X VGND VGND VPWR VPWR _5382_/X
+ sky130_fd_sc_hd__o311a_1
X_7121_ _7447_/CLK _7121_/D fanout598/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4333_ _4333_/A0 _5754_/A1 _4333_/S VGND VGND VPWR VPWR _4333_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5713__A _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4264_ _4264_/A0 _5754_/A1 _4264_/S VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__mux2_1
X_7052_ _7196_/CLK _7052_/D fanout590/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6003_ _6932_/Q _6751_/S _6051_/C _4117_/Y VGND VGND VPWR VPWR _6006_/A sky130_fd_sc_hd__o31ai_4
X_4195_ _4195_/A0 _5647_/A0 _4202_/S VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3880__A1 _7376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5859__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5082__B1 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5621__A2 _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6905_ _4127_/A1 _6905_/D _6855_/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5909__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6836_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6836_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout433_A _6404_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5385__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6582__B1 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6767_ _7030_/Q _6459_/B _6459_/C _6462_/X _7035_/Q VGND VGND VPWR VPWR _6767_/X
+ sky130_fd_sc_hd__a32o_1
X_3979_ _7439_/Q _3520_/X _3932_/X _3977_/X _3978_/X VGND VGND VPWR VPWR _3988_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_73_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5718_ _5754_/A1 _5718_/A1 _5721_/S VGND VGND VPWR VPWR _5718_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3935__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6698_ _6682_/X _6698_/B _6698_/C VGND VGND VPWR VPWR _6698_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5649_ _5998_/A1 _5649_/A1 _5649_/S VGND VGND VPWR VPWR _5649_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6334__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3408__A _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold250 hold250/A VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7319_ _7499_/CLK _7319_/D fanout578/X VGND VGND VPWR VPWR _7319_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold261 hold261/A VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold272 hold272/A VGND VGND VPWR VPWR hold272/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5623__A _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold283 hold283/A VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold294 hold294/A VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1715_A _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6637__A1 _7302_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5342__B _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input133_A wb_dat_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3871__A1 input47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5769__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6270__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5376__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3926__A2 _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4702__A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5391__A4 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6325__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output185_A _3426_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6628__A1 _7310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5300__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_2
XFILLER_0_188_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6800__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4406__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4951_ _4853_/Y _4936_/Y _4950_/Y _4681_/Y _4949_/Y VGND VGND VPWR VPWR _4958_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3902_ _7255_/Q _3557_/X _4521_/B _4340_/A _7017_/Q VGND VGND VPWR VPWR _3902_/X
+ sky130_fd_sc_hd__a32o_1
X_7670_ _7670_/A VGND VGND VPWR VPWR _7670_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4882_ _4932_/B _5342_/B VGND VGND VPWR VPWR _4882_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6159__A3 _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6621_ _7469_/Q _6434_/X _6616_/X _6617_/X _6620_/X VGND VGND VPWR VPWR _6621_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_157_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3833_ _7537_/Q _3590_/C _5947_/B _3675_/X _7189_/Q VGND VGND VPWR VPWR _3837_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6564__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3917__A2 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6552_ _7427_/Q _6463_/X _6467_/X _7419_/Q VGND VGND VPWR VPWR _6552_/X sky130_fd_sc_hd__a22o_1
X_3764_ input14/X _3490_/X _3760_/X _3761_/X _3763_/X VGND VGND VPWR VPWR _3764_/X
+ sky130_fd_sc_hd__a2111o_4
X_5503_ _4672_/X _4873_/X _4893_/Y _5340_/D _5438_/C VGND VGND VPWR VPWR _5550_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__6316__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6483_ _7352_/Q _6459_/B _6459_/C _6462_/X _7360_/Q VGND VGND VPWR VPWR _6483_/X
+ sky130_fd_sc_hd__a32o_1
X_3695_ _7467_/Q _3565_/X _3692_/X _3694_/X VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput300 _4173_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
XFILLER_0_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5434_ _4996_/A _5329_/X _5426_/X _5053_/C _5191_/X VGND VGND VPWR VPWR _5501_/A
+ sky130_fd_sc_hd__a221o_1
Xoutput311 _7628_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
Xoutput322 hold1177/X VGND VGND VPWR VPWR hold1178/A sky130_fd_sc_hd__buf_6
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput333 hold1181/X VGND VGND VPWR VPWR hold1182/A sky130_fd_sc_hd__buf_6
XFILLER_0_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5365_ _4601_/Y _4947_/Y _4949_/A VGND VGND VPWR VPWR _5367_/D sky130_fd_sc_hd__o21bai_2
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7496_/CLK sky130_fd_sc_hd__clkbuf_8
X_7104_ _7207_/CLK _7104_/D _4309_/B VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_4
X_4316_ _4321_/S _3795_/B _4315_/Y VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5296_ _4720_/Y _4755_/Y _4761_/Y _4692_/Y _5143_/A VGND VGND VPWR VPWR _5303_/A
+ sky130_fd_sc_hd__o221a_1
X_7035_ _7196_/CLK _7035_/D fanout588/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_4
X_4247_ _4247_/A0 _4246_/X _4249_/S VGND VGND VPWR VPWR _4247_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout383_A _3492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4178_ _4178_/A _7111_/Q VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__and2_1
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6252__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6819_ _6818_/X _6819_/A1 _6822_/S VGND VGND VPWR VPWR _7643_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6555__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3908__A2 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire427 _4753_/C VGND VGND VPWR VPWR _4694_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4879__D _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5530__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5072__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout571 fanout587/X VGND VGND VPWR VPWR _6871_/A sky130_fd_sc_hd__buf_12
Xfanout582 fanout587/X VGND VGND VPWR VPWR fanout582/X sky130_fd_sc_hd__buf_8
Xfanout593 fanout597/X VGND VGND VPWR VPWR fanout593/X sky130_fd_sc_hd__buf_12
XANTENNA__3844__A1 _7513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5597__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6546__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6561__A3 _6429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3480_ _3505_/C _3505_/D VGND VGND VPWR VPWR _3480_/X sky130_fd_sc_hd__and2_1
XANTENNA__6313__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _5150_/A _5150_/B _5150_/C VGND VGND VPWR VPWR _5153_/A sky130_fd_sc_hd__and3_1
Xhold2409 _7552_/Q VGND VGND VPWR VPWR hold618/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6078__B _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4101_ _7593_/Q _7594_/Q VGND VGND VPWR VPWR _6463_/A sky130_fd_sc_hd__and2b_4
XANTENNA__6077__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5081_ _5081_/A _5387_/D _5260_/C _5091_/A VGND VGND VPWR VPWR _5081_/Y sky130_fd_sc_hd__nand4_2
Xhold1708 _7164_/Q VGND VGND VPWR VPWR hold332/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1719 hold277/X VGND VGND VPWR VPWR _5996_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4032_ _6903_/Q _7074_/Q _4030_/Y _4031_/X VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_5_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5588__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5983_ _5983_/A _5992_/C hold48/X VGND VGND VPWR VPWR _5991_/S sky130_fd_sc_hd__and3_4
XANTENNA__3599__B1 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4934_ _4934_/A _4934_/B _4934_/C VGND VGND VPWR VPWR _4934_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4260__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7653_ _7653_/A VGND VGND VPWR VPWR _7653_/X sky130_fd_sc_hd__buf_2
X_4865_ _5183_/A _5053_/C VGND VGND VPWR VPWR _4865_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6537__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 _3972_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_34 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6604_ _7373_/Q _6413_/C _6651_/C _6603_/X VGND VGND VPWR VPWR _6604_/X sky130_fd_sc_hd__a31o_1
X_3816_ _7179_/Q _5947_/B _5619_/B _7401_/Q _5794_/A VGND VGND VPWR VPWR _3816_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7584_ _7586_/CLK _7584_/D _4128_/B VGND VGND VPWR VPWR _7584_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_45 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 _3965_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4796_ _5260_/A _4797_/B VGND VGND VPWR VPWR _4796_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_7_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_67 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6535_ _7298_/Q _6420_/A _6530_/X _6532_/X _6534_/X VGND VGND VPWR VPWR _6545_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_104_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3747_ _7185_/Q _4533_/A _3670_/X _7135_/Q _3746_/X VGND VGND VPWR VPWR _3747_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6466_ _7596_/Q _7595_/Q _6574_/B _6600_/B VGND VGND VPWR VPWR _6466_/X sky130_fd_sc_hd__and4_4
X_3678_ _7181_/Q _5938_/C _5619_/B _3647_/X _7171_/Q VGND VGND VPWR VPWR _3678_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5417_ _4695_/Y _4732_/Y _5317_/A VGND VGND VPWR VPWR _5532_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6397_ _6397_/A _6397_/B _6397_/C _6397_/D VGND VGND VPWR VPWR _6397_/Y sky130_fd_sc_hd__nor4_1
XANTENNA_fanout598_A fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput174 _4177_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
X_5348_ _5094_/A _5183_/C _5213_/C _4954_/C _5213_/B VGND VGND VPWR VPWR _5349_/B
+ sky130_fd_sc_hd__o2111a_1
Xoutput185 _3426_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 _3416_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XANTENNA__6068__A2 _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2910 hold2910/A VGND VGND VPWR VPWR _5795_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6419__D _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2921 _7432_/Q VGND VGND VPWR VPWR hold2921/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2932 hold2932/A VGND VGND VPWR VPWR _5769_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2943 _4399_/X VGND VGND VPWR VPWR hold701/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5279_ _4667_/B _4828_/Y _5278_/X VGND VGND VPWR VPWR _5279_/Y sky130_fd_sc_hd__o21ai_1
Xhold2954 _4417_/X VGND VGND VPWR VPWR hold2954/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7018_ _7211_/CLK _7018_/D fanout572/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfstp_2
Xhold2965 hold2965/A VGND VGND VPWR VPWR _5759_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2976 hold2976/A VGND VGND VPWR VPWR _4547_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2987 _7123_/Q VGND VGND VPWR VPWR hold2987/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2998 _7257_/Q VGND VGND VPWR VPWR _4078_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3421__A _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6435__C _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6776__B1 _6774_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6240__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4251__A1 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6451__B _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_191_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5751__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5782__S hold49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3762__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input61_A mgmt_gpio_in[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6700__B1 _6698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5267__B1 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout390 hold2225/X VGND VGND VPWR VPWR _5803_/A sky130_fd_sc_hd__buf_12
XFILLER_0_108_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6767__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6231__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4242__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6519__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5990__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2096_A _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4650_ _4591_/Y _4648_/A _4726_/B VGND VGND VPWR VPWR _4942_/A sky130_fd_sc_hd__o21a_4
XFILLER_0_182_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6080__C _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3601_ _6917_/Q _3527_/X _3597_/X _3598_/X _3600_/X VGND VGND VPWR VPWR _3606_/B
+ sky130_fd_sc_hd__a2111o_1
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR _3863_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5742__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4581_ _4887_/D _4747_/B _4887_/B _4879_/C VGND VGND VPWR VPWR _4626_/B sky130_fd_sc_hd__and4_4
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6320_ _7037_/Q _6144_/C _6084_/X _6072_/X _7153_/Q VGND VGND VPWR VPWR _6320_/X
+ sky130_fd_sc_hd__a32o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7672_/A sky130_fd_sc_hd__buf_4
XFILLER_0_24_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold805 hold805/A VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3532_ _4551_/A _3537_/A _5965_/A VGND VGND VPWR VPWR _3532_/X sky130_fd_sc_hd__and3_1
Xinput76 qspi_enabled VGND VGND VPWR VPWR _4142_/A sky130_fd_sc_hd__buf_12
Xhold816 hold816/A VGND VGND VPWR VPWR _7176_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7671_/A sky130_fd_sc_hd__buf_4
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold827 hold827/A VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6298__A2 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold838 hold838/A VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap557 _4583_/B VGND VGND VPWR VPWR _5301_/A1 sky130_fd_sc_hd__buf_8
X_6251_ _7349_/Q _6070_/X _6112_/X _7485_/Q _6250_/X VGND VGND VPWR VPWR _6257_/C
+ sky130_fd_sc_hd__a221o_1
Xhold849 hold849/A VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_150_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6089__A _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3463_ _3462_/X _3463_/A1 _4429_/B VGND VGND VPWR VPWR _3463_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3506__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5202_ _5202_/A _5202_/B _5202_/C VGND VGND VPWR VPWR _5202_/X sky130_fd_sc_hd__and3_1
XANTENNA__4848__A3 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6182_ _7426_/Q _6094_/A _6074_/X _6120_/X _7338_/Q VGND VGND VPWR VPWR _6182_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2206 hold878/X VGND VGND VPWR VPWR _4200_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2217 hold643/X VGND VGND VPWR VPWR _5912_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2228 _7326_/Q VGND VGND VPWR VPWR hold570/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5133_ _4888_/B _4879_/C _5091_/A _4940_/C VGND VGND VPWR VPWR _5134_/C sky130_fd_sc_hd__a31o_1
Xhold2239 _7344_/Q VGND VGND VPWR VPWR hold561/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1505 _5908_/X VGND VGND VPWR VPWR hold226/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1516 hold183/X VGND VGND VPWR VPWR _5923_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1527 hold31/X VGND VGND VPWR VPWR _5973_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5064_ _5064_/A _5064_/B _5064_/C VGND VGND VPWR VPWR _5064_/Y sky130_fd_sc_hd__nand3_1
Xhold1538 hold199/X VGND VGND VPWR VPWR _5959_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1549 hold271/X VGND VGND VPWR VPWR _5827_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4982__D _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4015_ _6903_/Q _6902_/Q _6901_/Q _6900_/Q VGND VGND VPWR VPWR _4025_/B sky130_fd_sc_hd__and4_2
XANTENNA__6470__A2 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4481__A1 _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7648__A _7648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5966_ _5966_/A0 _5993_/A1 hold13/X VGND VGND VPWR VPWR _5966_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4233__A1 _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4917_ _5213_/A _5213_/B _4929_/A _4937_/C VGND VGND VPWR VPWR _5573_/C sky130_fd_sc_hd__nand4_2
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5897_ _5987_/A1 _5897_/A1 _5901_/S VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7636_ _7636_/CLK _7636_/D VGND VGND VPWR VPWR _7636_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout513_A _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4848_ _5205_/A1 _4849_/B _5295_/C _4847_/X VGND VGND VPWR VPWR _4851_/B sky130_fd_sc_hd__a31oi_1
XFILLER_0_117_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4503__C _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6525__A3 _6429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5733__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7567_ _7572_/CLK _7567_/D fanout596/X VGND VGND VPWR VPWR _7567_/Q sky130_fd_sc_hd__dfstp_1
X_4779_ _4700_/Y _4774_/Y _4778_/Y _4776_/Y VGND VGND VPWR VPWR _4781_/B sky130_fd_sc_hd__o211ai_1
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6518_ _7393_/Q _6420_/C _6467_/X _7417_/Q _6517_/X VGND VGND VPWR VPWR _6518_/X
+ sky130_fd_sc_hd__a221o_1
X_7498_ _7513_/CLK _7498_/D fanout602/X VGND VGND VPWR VPWR _7498_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6289__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6449_ _7311_/Q _6419_/D _6425_/X _7335_/Q _6448_/X VGND VGND VPWR VPWR _6449_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3416__A _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7556_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5631__A _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2740 hold835/X VGND VGND VPWR VPWR _4405_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2751 _6923_/Q VGND VGND VPWR VPWR hold744/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2762 _6978_/Q VGND VGND VPWR VPWR _4288_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2773 hold2773/A VGND VGND VPWR VPWR _4474_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_55_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7501_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2784 _6977_/Q VGND VGND VPWR VPWR _4287_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5264__A3 _5102_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2795 _6994_/Q VGND VGND VPWR VPWR _4312_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6461__A2 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5777__S hold49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6213__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5724__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6401__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4710__A _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4160__B1 _4159_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6906__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4463__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6075__C _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6204__A2 _6093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5820_ _5820_/A0 _5955_/A1 _5820_/S VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5751_ _5751_/A0 _5967_/A1 _5757_/S VGND VGND VPWR VPWR _5751_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4604__B _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5963__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3974__B1 _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4702_ _4887_/D _4856_/A _4888_/B _4879_/C VGND VGND VPWR VPWR _4702_/Y sky130_fd_sc_hd__nor4_4
XFILLER_0_155_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5682_ _5682_/A0 hold84/X _5685_/S VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6507__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7421_ _7581_/CLK _7421_/D fanout585/X VGND VGND VPWR VPWR _7421_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4633_ _4768_/B _4694_/B VGND VGND VPWR VPWR _4802_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_71_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5138__D _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7352_ _7563_/CLK _7352_/D fanout598/X VGND VGND VPWR VPWR _7352_/Q sky130_fd_sc_hd__dfstp_2
X_4564_ _4564_/A _4564_/B _4564_/C _4564_/D VGND VGND VPWR VPWR _4565_/B sky130_fd_sc_hd__nand4_4
XANTENNA__5191__A2 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold602 hold602/A VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold613 hold613/A VGND VGND VPWR VPWR _6956_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold624 hold624/A VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6303_ _6303_/A _6303_/B _6303_/C _6303_/D VGND VGND VPWR VPWR _6303_/Y sky130_fd_sc_hd__nor4_1
X_3515_ _5640_/B _5612_/B _4388_/B VGND VGND VPWR VPWR _3515_/X sky130_fd_sc_hd__and3_4
Xhold635 hold635/A VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7283_ _7309_/CLK _7283_/D fanout576/X VGND VGND VPWR VPWR _7283_/Q sky130_fd_sc_hd__dfrtp_4
Xhold646 hold646/A VGND VGND VPWR VPWR _7236_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4495_ _4495_/A0 _5852_/A0 _4496_/S VGND VGND VPWR VPWR _4495_/X sky130_fd_sc_hd__mux2_1
Xhold657 hold657/A VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_100_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold668 hold668/A VGND VGND VPWR VPWR hold668/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold679 hold679/A VGND VGND VPWR VPWR _7225_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6234_ _6228_/X _6230_/X _6231_/X _6233_/X VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__a211o_1
X_3446_ _6910_/Q _6909_/Q _6908_/Q VGND VGND VPWR VPWR _3856_/A sky130_fd_sc_hd__nor3_4
XFILLER_0_100_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6140__B2 _7440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2003 hold135/X VGND VGND VPWR VPWR _4447_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6691__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5494__A3 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2014 _4206_/X VGND VGND VPWR VPWR hold495/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6165_ _7497_/Q _6332_/B _6084_/X _6100_/X _7473_/Q VGND VGND VPWR VPWR _6165_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_176_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 _4471_/X VGND VGND VPWR VPWR hold511/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2036 _7637_/Q VGND VGND VPWR VPWR hold462/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4993__C _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 hold3125/X VGND VGND VPWR VPWR hold3126/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2047 _4453_/X VGND VGND VPWR VPWR hold483/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1313 hold3062/X VGND VGND VPWR VPWR hold3063/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5116_ _4709_/Y _4826_/Y _4832_/Y _4828_/Y _4703_/Y VGND VGND VPWR VPWR _5116_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2058 _4495_/X VGND VGND VPWR VPWR hold509/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2069 hold82/X VGND VGND VPWR VPWR _4189_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1324 _4204_/X VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6096_ _7375_/Q _6090_/X _6092_/X _7527_/Q _6095_/X VGND VGND VPWR VPWR _6102_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1335 _4289_/A1 VGND VGND VPWR VPWR hold2809/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1346 _4281_/B VGND VGND VPWR VPWR hold2790/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1357 _4278_/B VGND VGND VPWR VPWR hold2853/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5246__A3 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5047_ _5047_/A _5047_/B _5047_/C VGND VGND VPWR VPWR _5051_/A sky130_fd_sc_hd__nor3_1
Xhold1368 hold1394/X VGND VGND VPWR VPWR hold1395/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5651__A0 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4454__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1379 hold1506/X VGND VGND VPWR VPWR hold1507/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4206__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6998_ _6999_/CLK _6998_/D VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6746__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5954__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5949_ _5949_/A0 _5967_/A1 _5955_/S VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold1480_A _7468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7619_ _7621_/CLK _7619_/D fanout579/X VGND VGND VPWR VPWR _7619_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5048__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4390__A0 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4887__D _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input163_A wb_dat_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6682__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3260 _6779_/X VGND VGND VPWR VPWR _7628_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3271 _4099_/Y VGND VGND VPWR VPWR _4112_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3282 _7391_/Q VGND VGND VPWR VPWR hold567/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2570 _7476_/Q VGND VGND VPWR VPWR hold2570/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input24_A mask_rev_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2581 _5837_/X VGND VGND VPWR VPWR hold806/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2592 hold2592/A VGND VGND VPWR VPWR _5696_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4445__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1880 _7194_/Q VGND VGND VPWR VPWR hold448/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_leaf_32_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1891 _7261_/Q VGND VGND VPWR VPWR hold348/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3799__A3 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6198__A1 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5945__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5173__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3723__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5970__S hold13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2059_A _7447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4280_ _3922_/Y _4280_/A1 _4289_/S VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4133__A0 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6673__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3487__A2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3503__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4436__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6921_ _7255_/CLK _6921_/D fanout565/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_77_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4615__A _4615_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6852_ _6871_/A _6872_/B VGND VGND VPWR VPWR _6852_/X sky130_fd_sc_hd__and2_1
XFILLER_0_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6728__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5803_ _5803_/A _5947_/A _5902_/B VGND VGND VPWR VPWR _5811_/S sky130_fd_sc_hd__and3_4
XFILLER_0_18_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6783_ _3922_/Y _6783_/A1 _6792_/S VGND VGND VPWR VPWR _7630_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4334__B _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3995_ _3926_/X _3995_/B _3995_/C _3995_/D VGND VGND VPWR VPWR _3996_/B sky130_fd_sc_hd__and4b_4
XANTENNA__3947__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5734_ _5734_/A0 _5950_/A1 _5739_/S VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5665_ _5665_/A0 _5953_/A1 _5667_/S VGND VGND VPWR VPWR _5665_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3962__A3 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4988__C _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7404_ _7501_/CLK _7404_/D fanout581/X VGND VGND VPWR VPWR _7404_/Q sky130_fd_sc_hd__dfrtp_4
X_4616_ _4643_/C _4645_/D VGND VGND VPWR VPWR _4616_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_13_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7498__RESET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5596_ _5612_/C _5596_/B _5640_/C _5640_/D VGND VGND VPWR VPWR _5602_/S sky130_fd_sc_hd__and4_4
XANTENNA__6361__B2 _6991_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold410 hold410/A VGND VGND VPWR VPWR hold410/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4372__A0 _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7335_ _7539_/CLK _7335_/D fanout577/X VGND VGND VPWR VPWR _7335_/Q sky130_fd_sc_hd__dfstp_2
Xhold421 hold421/A VGND VGND VPWR VPWR _7433_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4547_ _5583_/A0 _4547_/A1 _4550_/S VGND VGND VPWR VPWR _4547_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3714__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5880__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold432 hold432/A VGND VGND VPWR VPWR hold432/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7427__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold443 hold443/A VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold454 hold454/A VGND VGND VPWR VPWR hold454/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_3_5_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold465 hold465/A VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7266_ _7266_/CLK _7266_/D _6865_/A VGND VGND VPWR VPWR _7266_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6113__A1 _7367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4478_ _4478_/A0 _5586_/A0 _4478_/S VGND VGND VPWR VPWR _4478_/X sky130_fd_sc_hd__mux2_1
Xhold476 hold476/A VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold487 hold487/A VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold498 hold498/A VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6217_ _7460_/Q _6080_/X _6085_/X _7500_/Q _6216_/X VGND VGND VPWR VPWR _6217_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3429_ _7410_/Q VGND VGND VPWR VPWR _3429_/Y sky130_fd_sc_hd__clkinv_2
X_7197_ _7197_/CLK _7197_/D _6839_/A VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5612__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6148_ _7489_/Q _6112_/C _6332_/C _6116_/X _7313_/Q VGND VGND VPWR VPWR _6148_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _5904_/X VGND VGND VPWR VPWR _7496_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4509__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1121 hold2975/X VGND VGND VPWR VPWR hold2976/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1132 _4360_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 hold2987/X VGND VGND VPWR VPWR hold2988/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _7588_/Q _6119_/A _6106_/B _7589_/Q VGND VGND VPWR VPWR _6079_/X sky130_fd_sc_hd__and4bb_4
Xhold1154 hold1154/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 hold2787/X VGND VGND VPWR VPWR hold2788/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1176 hold1176/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
Xhold1187 hold2848/X VGND VGND VPWR VPWR hold1187/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 hold1198/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6443__C _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3953__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6352__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5155__A2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5790__S _5793_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6104__B2 _7399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5803__B _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6655__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5458__A3 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7107__CLK _4164_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5863__A0 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3090 _7192_/Q VGND VGND VPWR VPWR hold3090/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4418__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4969__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3641__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5918__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3780_ _7450_/Q _5848_/A _4545_/A _7195_/Q _3779_/X VGND VGND VPWR VPWR _3780_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6591__A1 _7452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6591__B2 _7524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2176_A _7334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5450_ _5226_/X _5450_/B _5450_/C VGND VGND VPWR VPWR _5574_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4401_ _4401_/A0 _5714_/A0 _4405_/S VGND VGND VPWR VPWR _4401_/X sky130_fd_sc_hd__mux2_1
X_5381_ _4700_/Y _5451_/A1 _4720_/Y _5081_/Y VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__o31a_1
X_7120_ _7447_/CLK _7120_/D fanout601/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfstp_2
Xclkbuf_3_2_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4332_ _4332_/A0 _5647_/A0 _4333_/S VGND VGND VPWR VPWR _4332_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5713__B hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7051_ _7189_/CLK _7051_/D fanout572/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6646__A2 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4263_ _4263_/A0 _5647_/A0 _4264_/S VGND VGND VPWR VPWR _4263_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3514__A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5854__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6002_ _6065_/C _6929_/Q _7256_/Q _6001_/Y _6002_/B2 VGND VGND VPWR VPWR _7583_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA_hold2608_A _7515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4194_ _4194_/A0 _5950_/A1 _4202_/S VGND VGND VPWR VPWR _4194_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3880__A2 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6904_ _4150_/A1 _6904_/D _6854_/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6835_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6835_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6766_ _7171_/Q _6408_/D _6454_/X _7070_/Q _6765_/X VGND VGND VPWR VPWR _6773_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3978_ _7172_/Q _4509_/A _5623_/B _3649_/X _7066_/Q VGND VGND VPWR VPWR _3978_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_175_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5717_ _5951_/A1 _5717_/A1 _5721_/S VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6697_ _6697_/A _6697_/B _6697_/C _6697_/D VGND VGND VPWR VPWR _6698_/C sky130_fd_sc_hd__nor4_2
XANTENNA__3935__A3 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _7075_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5648_ _5997_/A1 _5648_/A1 _5649_/S VGND VGND VPWR VPWR _5648_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4345__A0 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5579_ _5385_/X _5520_/Y _5564_/Y _5578_/Y _5560_/X VGND VGND VPWR VPWR _5579_/X
+ sky130_fd_sc_hd__o41a_2
XANTENNA__3699__A2 _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7318_ _7582_/CLK _7318_/D fanout584/X VGND VGND VPWR VPWR _7318_/Q sky130_fd_sc_hd__dfrtp_4
Xhold240 hold240/A VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold251 hold251/A VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold262 hold262/A VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold273 hold273/A VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6098__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold284 _4078_/B VGND VGND VPWR VPWR hold284/X sky130_fd_sc_hd__buf_6
XANTENNA__5623__B _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6637__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7249_ _7266_/CLK _7249_/D fanout567/X VGND VGND VPWR VPWR _7648_/A sky130_fd_sc_hd__dfrtp_4
Xhold295 _5672_/X VGND VGND VPWR VPWR _7290_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3424__A _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3871__A2 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input126_A wb_adr_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6454__B _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6270__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5376__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input91_A spimemio_flash_io3_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3926__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4702__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5086__A _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6325__A1 _7198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6325__B2 _7027_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6628__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4639__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5300__A2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_188_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4950_ _4966_/A _5222_/B _5222_/C _5094_/A VGND VGND VPWR VPWR _4950_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_188_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3614__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3901_ _7052_/Q _4509_/A _3548_/X _3900_/X VGND VGND VPWR VPWR _3901_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_47_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _4942_/A _4948_/C _5342_/B VGND VGND VPWR VPWR _4943_/B sky130_fd_sc_hd__and3_2
XFILLER_0_143_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6159__A4 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6620_ _7413_/Q _6468_/X _6618_/X _6619_/X _6430_/X VGND VGND VPWR VPWR _6620_/X
+ sky130_fd_sc_hd__a2111o_1
X_3832_ _7457_/Q _3933_/A _5875_/A _3537_/X _7425_/Q VGND VGND VPWR VPWR _3837_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_172_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6564__A1 _7299_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6551_ _7331_/Q _6423_/X _6452_/X _7347_/Q _6550_/X VGND VGND VPWR VPWR _6551_/X
+ sky130_fd_sc_hd__a221o_1
X_3763_ input23/X _3488_/X _3521_/X _7314_/Q _3762_/X VGND VGND VPWR VPWR _3763_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5502_ _4679_/Y _4832_/Y _5528_/A3 _5438_/B _5200_/B VGND VGND VPWR VPWR _5550_/A
+ sky130_fd_sc_hd__o311a_1
XANTENNA_clkbuf_leaf_1_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6482_ _7392_/Q _6420_/C _6419_/A _7544_/Q _6481_/X VGND VGND VPWR VPWR _6482_/X
+ sky130_fd_sc_hd__a221o_2
X_3694_ _7020_/Q _3669_/C _5619_/B _3693_/X VGND VGND VPWR VPWR _3694_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6316__B2 _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4327__A0 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5433_ _5331_/Y _5554_/B _5433_/C VGND VGND VPWR VPWR _5435_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput301 _4117_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
XFILLER_0_11_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput312 hold2820/X VGND VGND VPWR VPWR hold1168/A sky130_fd_sc_hd__buf_6
Xoutput323 hold2797/X VGND VGND VPWR VPWR hold1160/A sky130_fd_sc_hd__buf_6
Xoutput334 hold2788/X VGND VGND VPWR VPWR hold1166/A sky130_fd_sc_hd__buf_6
X_5364_ _5094_/A wire533/X _5248_/C _4935_/X VGND VGND VPWR VPWR _5545_/B sky130_fd_sc_hd__o31a_1
X_7103_ _7207_/CLK _7103_/D _6780_/B VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6619__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4315_ _4321_/S _4315_/B VGND VGND VPWR VPWR _4315_/Y sky130_fd_sc_hd__nand2_1
X_5295_ _5295_/A _5295_/B _5295_/C _5295_/D VGND VGND VPWR VPWR _5422_/D sky130_fd_sc_hd__nand4_2
X_7034_ _7112_/CLK _7034_/D fanout589/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_4
X_4246_ _5657_/A1 _5954_/A1 _4248_/S VGND VGND VPWR VPWR _4246_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6095__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4177_ _7264_/Q _4177_/B VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__and2_2
XFILLER_0_93_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6252__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6818_ _7109_/Q _6818_/A2 _6818_/B1 wire463/A _6817_/X VGND VGND VPWR VPWR _6818_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5358__A2 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire406 _3505_/Y VGND VGND VPWR VPWR wire406/X sky130_fd_sc_hd__buf_2
XFILLER_0_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6749_ _6749_/A _6749_/B _6749_/C _6749_/D VGND VGND VPWR VPWR _6749_/Y sky130_fd_sc_hd__nor4_4
XANTENNA__3419__A _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout561 _4747_/B VGND VGND VPWR VPWR _4856_/A sky130_fd_sc_hd__buf_12
Xfanout572 fanout574/X VGND VGND VPWR VPWR fanout572/X sky130_fd_sc_hd__buf_12
XANTENNA__6491__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout583 fanout585/X VGND VGND VPWR VPWR fanout583/X sky130_fd_sc_hd__buf_12
Xfanout594 fanout597/X VGND VGND VPWR VPWR fanout594/X sky130_fd_sc_hd__buf_12
XANTENNA__3844__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4819__A_N _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output295_A _7244_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3780__A1 _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4100_ _7584_/Q _7586_/Q _7587_/Q _4099_/D _6932_/Q VGND VGND VPWR VPWR _4100_/X
+ sky130_fd_sc_hd__o41a_1
X_5080_ _5563_/A1 _4737_/Y _4946_/Y _5077_/Y _4748_/Y VGND VGND VPWR VPWR _5084_/C
+ sky130_fd_sc_hd__o32a_1
Xhold1709 hold332/X VGND VGND VPWR VPWR _4512_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6482__B1 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4031_ _6903_/Q _6902_/Q _6901_/Q _6900_/Q _6904_/Q VGND VGND VPWR VPWR _4031_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__3835__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6785__A1 _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5982_ hold17/X _5982_/A1 _5982_/S VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_189_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4933_ _4933_/A _4933_/B _5260_/D VGND VGND VPWR VPWR _4934_/B sky130_fd_sc_hd__and3_1
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7652_ _7652_/A VGND VGND VPWR VPWR _7652_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4864_ _5328_/A _5328_/B _5053_/C VGND VGND VPWR VPWR _5180_/A sky130_fd_sc_hd__and3_4
XANTENNA__6537__A1 _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6537__B2 _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_13 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4548__A0 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3815_ _6913_/Q _3527_/X _4340_/A _7018_/Q _3814_/X VGND VGND VPWR VPWR _3815_/X
+ sky130_fd_sc_hd__a221o_1
X_6603_ _7477_/Q _6574_/B _6441_/X _6058_/X _7533_/Q VGND VGND VPWR VPWR _6603_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_24 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7583_ _7586_/CLK _7583_/D _6865_/A VGND VGND VPWR VPWR _7583_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_35 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_46 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _4740_/D _4984_/B _4795_/C _4814_/C VGND VGND VPWR VPWR _4799_/C sky130_fd_sc_hd__and4bb_4
XFILLER_0_55_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_57 _4859_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_68 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _7538_/Q _6408_/D _6425_/X _7338_/Q _6533_/X VGND VGND VPWR VPWR _6534_/X
+ sky130_fd_sc_hd__a221o_1
X_3746_ _7394_/Q _4473_/A _5785_/B _3665_/X _7125_/Q VGND VGND VPWR VPWR _3746_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3771__A1 _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6465_ _7303_/Q _6420_/B _6462_/X _7359_/Q _6464_/X VGND VGND VPWR VPWR _6471_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3677_ _7539_/Q _3590_/C _5947_/B _3569_/X hold96/A VGND VGND VPWR VPWR _3677_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4996__C _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5416_ _5535_/A _5416_/B _5535_/B VGND VGND VPWR VPWR _5419_/B sky130_fd_sc_hd__and3_1
XFILLER_0_11_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6396_ _7025_/Q _6070_/X _6080_/X _7201_/Q _6395_/X VGND VGND VPWR VPWR _6397_/D
+ sky130_fd_sc_hd__a221o_1
X_5347_ _4947_/C _4933_/A _5346_/X _5208_/Y VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout493_A hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput175 _4160_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput186 _4158_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3442_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
Xhold2900 _6987_/Q VGND VGND VPWR VPWR _4302_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2911 _6997_/Q VGND VGND VPWR VPWR _4317_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2922 hold2922/A VGND VGND VPWR VPWR _5832_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5278_ _5277_/X _5278_/B _5278_/C _5278_/D VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__and4b_1
Xhold2933 _7027_/Q VGND VGND VPWR VPWR hold2933/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2944 _7656_/A VGND VGND VPWR VPWR hold2944/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6473__B1 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2955 _7331_/Q VGND VGND VPWR VPWR hold716/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_7017_ _7170_/CLK hold66/X fanout573/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2966 _5759_/X VGND VGND VPWR VPWR _7367_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4229_ _4257_/A0 hold61/X _4231_/S VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__mux2_1
Xhold2977 _4547_/X VGND VGND VPWR VPWR hold2977/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3826__A2 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2988 hold2988/A VGND VGND VPWR VPWR _4463_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2999 _4406_/A1 VGND VGND VPWR VPWR _5633_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6225__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6435__D _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6776__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6240__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6528__A1 _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6451__C _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5067__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3762__A1 _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3762__B2 _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input54_A mgmt_gpio_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6464__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout380 _4491_/B VGND VGND VPWR VPWR _5992_/C sky130_fd_sc_hd__buf_8
XANTENNA__4708__A _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3817__A2 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout391 hold2225/X VGND VGND VPWR VPWR _4473_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4427__B _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6216__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output308_A _4135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6231__A3 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5973__S hold13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3600_ _7341_/Q _3531_/X _3545_/X _7349_/Q _3599_/X VGND VGND VPWR VPWR _3600_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4580_ _4795_/C _4740_/D _4772_/A _4805_/B VGND VGND VPWR VPWR _4646_/A sky130_fd_sc_hd__nand4_4
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__buf_2
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_2
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_2
X_3531_ _5722_/A _5640_/B _5731_/B VGND VGND VPWR VPWR _3531_/X sky130_fd_sc_hd__and3_4
XFILLER_0_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3753__A1 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7673_/A sky130_fd_sc_hd__buf_6
XFILLER_0_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3753__B2 _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold806 hold806/A VGND VGND VPWR VPWR _7437_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold817 hold817/A VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _4131_/B sky130_fd_sc_hd__buf_4
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold828 _5999_/X VGND VGND VPWR VPWR _7581_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold839 hold839/A VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2256_A _7328_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6250_ _7493_/Q _6112_/C _6332_/C _6097_/X _7445_/Q VGND VGND VPWR VPWR _6250_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap547 _4810_/C VGND VGND VPWR VPWR wire546/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3462_ _6902_/Q _6901_/Q _4025_/A VGND VGND VPWR VPWR _3462_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6089__B _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5201_ _5342_/A _5113_/A wire536/X _5058_/C _5158_/A VGND VGND VPWR VPWR _5202_/B
+ sky130_fd_sc_hd__a32oi_2
XFILLER_0_149_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3506__B hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6181_ _7530_/Q _6091_/X _6179_/X _6180_/X VGND VGND VPWR VPWR _6181_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5132_ _4722_/Y _4727_/Y _4761_/Y _4978_/Y VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__o22a_1
Xhold2207 _4200_/X VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2218 _7286_/Q VGND VGND VPWR VPWR hold522/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2229 hold570/X VGND VGND VPWR VPWR _5712_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1506 _7566_/Q VGND VGND VPWR VPWR hold1506/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1517 _5923_/X VGND VGND VPWR VPWR hold184/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5063_ _5342_/A _5203_/B _5183_/C _5339_/D VGND VGND VPWR VPWR _5064_/C sky130_fd_sc_hd__nand4_1
Xhold1528 _5973_/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3808__A2 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1539 _5959_/X VGND VGND VPWR VPWR hold200/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4014_ _4040_/D _4014_/B VGND VGND VPWR VPWR _4040_/A sky130_fd_sc_hd__nand2_4
XANTENNA__6207__B1 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2792_A _7182_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6222__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5965_ _5965_/A hold12/X hold48/A VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__and3_1
XFILLER_0_149_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4916_ _4916_/A _4916_/B _4916_/C VGND VGND VPWR VPWR _4919_/A sky130_fd_sc_hd__nor3_1
X_5896_ _5896_/A0 _5896_/A1 _5901_/S VGND VGND VPWR VPWR _5896_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3992__A1 _7367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7635_ _7636_/CLK _7635_/D VGND VGND VPWR VPWR _7635_/Q sky130_fd_sc_hd__dfxtp_1
X_4847_ _5107_/A _5118_/B _5453_/C VGND VGND VPWR VPWR _4847_/X sky130_fd_sc_hd__and3_2
XANTENNA__5883__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4778_ _4778_/A _5387_/C _5113_/A _5410_/B VGND VGND VPWR VPWR _4778_/Y sky130_fd_sc_hd__nand4_1
X_7566_ _7566_/CLK hold18/X fanout603/X VGND VGND VPWR VPWR _7566_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_133_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3744__A1 _7546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6517_ _7497_/Q _6600_/B _6651_/C _6452_/X _7345_/Q VGND VGND VPWR VPWR _6517_/X
+ sky130_fd_sc_hd__a32o_1
X_3729_ _7131_/Q _5830_/C _4491_/A _4491_/B _3728_/X VGND VGND VPWR VPWR _3729_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7497_ _7539_/CLK _7497_/D fanout577/X VGND VGND VPWR VPWR _7497_/Q sky130_fd_sc_hd__dfrtp_4
X_6448_ _7439_/Q _6424_/C _6771_/A3 _6446_/X _7519_/Q VGND VGND VPWR VPWR _6448_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6694__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6379_ _7015_/Q _6136_/B _6120_/B _6379_/B1 _7126_/Q VGND VGND VPWR VPWR _6379_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2730 _4538_/X VGND VGND VPWR VPWR hold838/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2741 _7303_/Q VGND VGND VPWR VPWR hold2741/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2752 hold744/X VGND VGND VPWR VPWR _4208_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2763 hold2763/A VGND VGND VPWR VPWR hold2763/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6446__C _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2774 _7172_/Q VGND VGND VPWR VPWR hold2774/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2785 hold2785/A VGND VGND VPWR VPWR hold2785/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2796 hold2796/A VGND VGND VPWR VPWR hold2796/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6462__B _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3578__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5421__B2 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3983__A1 _7343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5793__S _5793_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5094__A _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6685__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3499__B1 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output258_A _7243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6437__B1 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5660__A1 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5968__S hold13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3996__B _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4215__A2 _4078_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5750_ _5750_/A0 _5903_/A0 _5757_/S VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4173__A _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6091__C _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4701_ _4888_/B _5282_/A VGND VGND VPWR VPWR _5072_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_127_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_173_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5681_ _5681_/A0 _5951_/A1 _5685_/S VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4632_ _4740_/D _4984_/C _4628_/Y _4631_/Y VGND VGND VPWR VPWR _4753_/C sky130_fd_sc_hd__o31ai_4
X_7420_ _7581_/CLK _7420_/D fanout584/X VGND VGND VPWR VPWR _7420_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_170_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6373__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3726__A1 _7307_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4563_ _4563_/A _4563_/B _4563_/C _4563_/D VGND VGND VPWR VPWR _4565_/A sky130_fd_sc_hd__nand4_4
XANTENNA__3726__B2 _7025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7351_ _7395_/CLK _7351_/D fanout598/X VGND VGND VPWR VPWR _7351_/Q sky130_fd_sc_hd__dfstp_2
Xhold603 _5811_/X VGND VGND VPWR VPWR _7414_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5191__A3 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold614 hold614/A VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6302_ _7162_/Q _6075_/X _6099_/X _7026_/Q _6301_/X VGND VGND VPWR VPWR _6303_/D
+ sky130_fd_sc_hd__a221o_1
X_3514_ _5938_/B _3576_/B _3576_/C VGND VGND VPWR VPWR _3514_/X sky130_fd_sc_hd__and3_2
XFILLER_0_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold625 hold625/A VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7282_ _7309_/CLK _7282_/D fanout576/X VGND VGND VPWR VPWR _7282_/Q sky130_fd_sc_hd__dfrtp_4
X_4494_ _4494_/A0 _5914_/A1 _4496_/S VGND VGND VPWR VPWR _4494_/X sky130_fd_sc_hd__mux2_1
Xhold636 _4481_/X VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3741__A4 _3502_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold647 hold647/A VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5479__A1 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold658 hold658/A VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6233_ _7340_/Q _6120_/X _6121_/X _7308_/Q _6232_/X VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__a221o_1
X_3445_ _4805_/B VGND VGND VPWR VPWR _4814_/C sky130_fd_sc_hd__inv_16
Xhold669 _4324_/X VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6140__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap399 _4997_/B VGND VGND VPWR VPWR _4932_/B sky130_fd_sc_hd__buf_6
XANTENNA__4151__A1 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2004 _4447_/X VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6121_/C _6071_/X _7289_/Q _6097_/X _7441_/Q VGND VGND VPWR VPWR _6164_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2015 _7426_/Q VGND VGND VPWR VPWR hold430/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2026 _7144_/Q VGND VGND VPWR VPWR hold608/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2037 hold462/X VGND VGND VPWR VPWR _4181_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_176_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5115_/A _5115_/B _5282_/D VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__and3_2
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 hold3127/X VGND VGND VPWR VPWR _7222_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2048 _7140_/Q VGND VGND VPWR VPWR hold490/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 _5644_/X VGND VGND VPWR VPWR _7265_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6095_ _7487_/Q _6110_/A _6332_/C _6094_/X _7503_/Q VGND VGND VPWR VPWR _6095_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2059 _7447_/Q VGND VGND VPWR VPWR hold622/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 hold3155/X VGND VGND VPWR VPWR hold3156/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1336 _4288_/A1 VGND VGND VPWR VPWR hold2763/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1347 _4293_/A1 VGND VGND VPWR VPWR hold2801/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5046_ _5046_/A _5046_/B VGND VGND VPWR VPWR _5047_/B sky130_fd_sc_hd__nor2_1
Xhold1358 _4298_/B VGND VGND VPWR VPWR hold2871/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1369 hold2118/X VGND VGND VPWR VPWR hold2119/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5878__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6997_ _7633_/CLK _6997_/D VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5403__B2 _4428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5948_ _5948_/A0 _5948_/A1 _5955_/S VGND VGND VPWR VPWR _5948_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_164_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5879_ _5879_/A0 _5987_/A1 _5883_/S VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7618_ _7621_/CLK _7618_/D fanout576/X VGND VGND VPWR VPWR _7618_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3717__A1 _7459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7549_ _7555_/CLK _7549_/D fanout594/X VGND VGND VPWR VPWR _7549_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_133_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6667__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6131__A2 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input156_A wb_dat_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3250 _6896_/Q VGND VGND VPWR VPWR _4051_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6457__B _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3261 _6902_/Q VGND VGND VPWR VPWR _4039_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5890__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3272 _4112_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3283 _7074_/Q VGND VGND VPWR VPWR hold3283/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2560 hold2560/A VGND VGND VPWR VPWR _5746_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2571 hold2571/A VGND VGND VPWR VPWR _5881_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2582 _7397_/Q VGND VGND VPWR VPWR hold813/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2593 _7301_/Q VGND VGND VPWR VPWR hold807/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5788__S _5793_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5642__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1870 _5855_/X VGND VGND VPWR VPWR hold121/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input17_A mask_rev_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1881 hold448/X VGND VGND VPWR VPWR _4548_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1892 hold348/X VGND VGND VPWR VPWR _5638_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4705__B _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6198__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__B2 _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3708__A1 input7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3708__B2 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5173__A3 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4381__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6658__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4133__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6673__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5881__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6086__C _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3503__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5633__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6920_ _6926_/CLK _6920_/D fanout565/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6851_ _6873_/A _6872_/B VGND VGND VPWR VPWR _6851_/X sky130_fd_sc_hd__and2_1
XANTENNA__4615__B _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5802_ _5955_/A1 _5802_/A1 _5802_/S VGND VGND VPWR VPWR _5802_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3994_ input34/X _3486_/X _3990_/X _3992_/X _3993_/X VGND VGND VPWR VPWR _3995_/D
+ sky130_fd_sc_hd__a2111oi_4
X_6782_ _6792_/S _3996_/B _6781_/Y VGND VGND VPWR VPWR _7629_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5733_ _5733_/A0 _5967_/A1 _5739_/S VGND VGND VPWR VPWR _5733_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5664_ _5664_/A0 hold84/X _5667_/S VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7403_ _7432_/CLK _7403_/D fanout593/X VGND VGND VPWR VPWR _7403_/Q sky130_fd_sc_hd__dfrtp_4
X_4615_ _4615_/A _4645_/D VGND VGND VPWR VPWR _4615_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_54_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7366_/CLK sky130_fd_sc_hd__clkbuf_16
X_5595_ _5595_/A0 _5754_/A1 _5595_/S VGND VGND VPWR VPWR _5595_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_142_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold400 _3477_/Y VGND VGND VPWR VPWR hold400/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_111_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7334_ _7366_/CLK _7334_/D fanout579/X VGND VGND VPWR VPWR _7334_/Q sky130_fd_sc_hd__dfrtp_4
X_4546_ _5714_/A0 _4546_/A1 _4550_/S VGND VGND VPWR VPWR _4546_/X sky130_fd_sc_hd__mux2_1
Xhold411 hold411/A VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold422 hold422/A VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold433 hold433/A VGND VGND VPWR VPWR _7321_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold444 hold444/A VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold455 hold455/A VGND VGND VPWR VPWR _7406_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7265_ _7266_/CLK _7265_/D _6865_/A VGND VGND VPWR VPWR _7265_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6113__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4477_ _4477_/A0 _5852_/A0 _4478_/S VGND VGND VPWR VPWR _4477_/X sky130_fd_sc_hd__mux2_1
Xhold466 hold466/A VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold477 hold477/A VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold488 hold488/A VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3428_ _7418_/Q VGND VGND VPWR VPWR _3428_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_69_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7363_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold499 hold499/A VGND VGND VPWR VPWR _7425_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6216_ _7492_/Q _6094_/A _6332_/C _6097_/X _7444_/Q VGND VGND VPWR VPWR _6216_/X
+ sky130_fd_sc_hd__a32o_1
X_7196_ _7196_/CLK _7196_/D fanout590/X VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6664__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5872__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6146_/X _6145_/Y _6069_/X _6169_/A2 VGND VGND VPWR VPWR _7603_/D sky130_fd_sc_hd__o2bb2a_1
XANTENNA_input9_A mask_rev_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5612__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1100 hold2931/X VGND VGND VPWR VPWR hold2932/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 hold2991/X VGND VGND VPWR VPWR hold2992/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4509__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1122 hold2977/X VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1133 hold2909/X VGND VGND VPWR VPWR hold2910/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _6119_/A _6106_/B VGND VGND VPWR VPWR _6078_/X sky130_fd_sc_hd__and2b_4
Xhold1144 _4463_/X VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 hold2785/X VGND VGND VPWR VPWR hold1155/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5624__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1166 hold1166/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
X_5029_ _5138_/D _5038_/B _5030_/C VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__and3_1
Xhold1177 hold2828/X VGND VGND VPWR VPWR hold1177/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1188 hold1188/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4806__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1199 hold2877/X VGND VGND VPWR VPWR hold1199/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3938__A1 _7243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_192_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6352__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4899__C1 wire533/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4363__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6468__A _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6104__A2 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5803__C _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6655__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5091__B _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3080 _7633_/Q VGND VGND VPWR VPWR _6788_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3091 hold3091/A VGND VGND VPWR VPWR _4546_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2390 hold945/X VGND VGND VPWR VPWR _4326_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5615__A1 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3626__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_184_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6591__A2 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4170__B _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6343__A2 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4400_ _5612_/C hold56/X _5596_/B _5640_/D VGND VGND VPWR VPWR _4405_/S sky130_fd_sc_hd__and4_4
XFILLER_0_2_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4354__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5380_ _5255_/X _4844_/Y _4703_/Y _4737_/Y _5451_/A1 VGND VGND VPWR VPWR _5380_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_23_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4331_ _4331_/A0 _5815_/A1 _4333_/S VGND VGND VPWR VPWR _4331_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5282__A _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7050_ _7151_/CLK _7050_/D fanout593/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_4
X_4262_ _4262_/A0 _5950_/A1 _4264_/S VGND VGND VPWR VPWR _4262_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6097__B _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6001_ _6932_/Q _6929_/Q _4100_/X VGND VGND VPWR VPWR _6001_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4193_ _4193_/A0 _5805_/A1 _4202_/S VGND VGND VPWR VPWR _4193_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5606__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4626__A _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3530__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5082__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6903_ _4150_/A1 _6903_/D _6853_/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_173_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6834_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6834_/X sky130_fd_sc_hd__and2_1
XFILLER_0_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6765_ _6992_/Q _6420_/B _6460_/X _7116_/Q VGND VGND VPWR VPWR _6765_/X sky130_fd_sc_hd__a22o_1
X_3977_ _6927_/Q _4212_/A _5659_/B _3682_/X _7224_/Q VGND VGND VPWR VPWR _3977_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__6582__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5716_ _5896_/A0 _5716_/A1 _5721_/S VGND VGND VPWR VPWR _5716_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_190_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6696_ _6989_/Q _6420_/B _6422_/X _6963_/Q _6695_/X VGND VGND VPWR VPWR _6697_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout419_A _3569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5647_ _5647_/A0 _5647_/A1 _5649_/S VGND VGND VPWR VPWR _5647_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6334__A2 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7672__A _7672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5578_ _4707_/Y _4722_/Y _5089_/Y _5254_/X _5474_/C VGND VGND VPWR VPWR _5578_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA_clkbuf_leaf_75_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold230 hold230/A VGND VGND VPWR VPWR hold230/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3699__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold241 hold241/A VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7317_ _7478_/CLK _7317_/D fanout580/X VGND VGND VPWR VPWR _7317_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4529_ _4529_/A0 _5805_/A1 _4532_/S VGND VGND VPWR VPWR _4529_/X sky130_fd_sc_hd__mux2_1
Xhold252 hold252/A VGND VGND VPWR VPWR _7436_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold263 hold263/A VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6098__A1 _7407_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold274 hold274/A VGND VGND VPWR VPWR _7240_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6098__B2 _7439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold285 hold285/A VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4300__S _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7248_ _7266_/CLK _7248_/D _6865_/A VGND VGND VPWR VPWR _7248_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5623__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold296 hold296/A VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5845__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7179_ _7268_/CLK _7179_/D _6871_/A VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5920__A _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3440__A _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6454__C _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A wb_adr_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4271__A _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5781__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4702__C _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input84_A spimemio_flash_csb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4336__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5836__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6645__B _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_188_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_176_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3614__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3900_ _7067_/Q _3649_/X _3675_/X _7188_/Q VGND VGND VPWR VPWR _3900_/X sky130_fd_sc_hd__a22o_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ _5282_/A _5199_/C VGND VGND VPWR VPWR _4880_/Y sky130_fd_sc_hd__nand2_4
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3831_ _7409_/Q _3493_/X _3657_/X _6959_/Q _3830_/X VGND VGND VPWR VPWR _3837_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6564__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2286_A _7347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3762_ _7474_/Q _3494_/X _5704_/A _7322_/Q _3737_/X VGND VGND VPWR VPWR _3762_/X
+ sky130_fd_sc_hd__a221o_4
X_6550_ _7451_/Q _6467_/A _6771_/A3 _6446_/X _7523_/Q VGND VGND VPWR VPWR _6550_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5501_ _5501_/A _5501_/B VGND VGND VPWR VPWR _5504_/B sky130_fd_sc_hd__nor2_1
X_3693_ _7347_/Q _3590_/C _3669_/C _3659_/X _7010_/Q VGND VGND VPWR VPWR _3693_/X
+ sky130_fd_sc_hd__a32o_1
X_6481_ _7456_/Q _6463_/A _6574_/C _6425_/X _7336_/Q VGND VGND VPWR VPWR _6481_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6316__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5432_ _4667_/B _4821_/Y _5174_/Y _5012_/Y VGND VGND VPWR VPWR _5433_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput302 _3619_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
Xoutput313 hold2817/X VGND VGND VPWR VPWR hold1190/A sky130_fd_sc_hd__buf_6
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput324 hold1209/X VGND VGND VPWR VPWR hold1210/A sky130_fd_sc_hd__buf_6
X_5363_ _5347_/X _5363_/B _5510_/A VGND VGND VPWR VPWR _5367_/C sky130_fd_sc_hd__nand3b_1
Xoutput335 hold1207/X VGND VGND VPWR VPWR hold1208/A sky130_fd_sc_hd__buf_6
XFILLER_0_50_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3525__A hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7102_ _7207_/CLK _7102_/D _4309_/B VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfrtp_4
X_4314_ _4321_/S _3856_/B _4313_/Y VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__o21ai_1
X_5294_ _5294_/A _5294_/B _5294_/C VGND VGND VPWR VPWR _5294_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__5827__A1 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4245_ _4245_/A0 _4244_/X _4249_/S VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
X_7033_ _7176_/CLK _7033_/D fanout588/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5740__A _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4176_ _7263_/Q _4176_/B VGND VGND VPWR VPWR _4176_/X sky130_fd_sc_hd__and2_2
XFILLER_0_93_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_184_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6004__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ _7111_/Q _6817_/A2 _6817_/B1 _7110_/Q VGND VGND VPWR VPWR _6817_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_77_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6555__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5358__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5763__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6748_ _7024_/Q _6452_/X _6747_/X _6746_/X _6745_/X VGND VGND VPWR VPWR _6749_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire429 _4614_/Y VGND VGND VPWR VPWR _4947_/C sky130_fd_sc_hd__buf_6
X_6679_ _7148_/Q _6408_/A _6451_/X _6875_/Q _6678_/X VGND VGND VPWR VPWR _6679_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7423__SET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4318__A1 _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7482__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3435__A _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5818__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3829__B1 _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6491__A1 _7464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout562 input99/X VGND VGND VPWR VPWR _4747_/B sky130_fd_sc_hd__buf_12
Xfanout573 fanout574/X VGND VGND VPWR VPWR fanout573/X sky130_fd_sc_hd__buf_12
Xmgmt_gpio_14_buff_inst _4162_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_8
Xfanout584 fanout585/X VGND VGND VPWR VPWR fanout584/X sky130_fd_sc_hd__buf_12
Xfanout595 fanout596/X VGND VGND VPWR VPWR fanout595/X sky130_fd_sc_hd__buf_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5796__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6546__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3780__A2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5809__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4030_ _6904_/Q _4025_/B _4025_/A VGND VGND VPWR VPWR _4030_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6482__A1 _7392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3835__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_23_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5981_ hold61/X _5981_/A1 _5982_/S VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6785__A2 _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3599__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4932_ _4947_/C _4932_/B _4933_/A _4940_/C VGND VGND VPWR VPWR _4932_/X sky130_fd_sc_hd__and4_1
XFILLER_0_86_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7651_ _7651_/A VGND VGND VPWR VPWR _7651_/X sky130_fd_sc_hd__clkbuf_2
X_4863_ _4805_/B _4668_/C _4660_/Y VGND VGND VPWR VPWR _5053_/C sky130_fd_sc_hd__o21a_4
XANTENNA__4623__B _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6537__A2 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6602_ _7349_/Q _6452_/X _6463_/X _7429_/Q VGND VGND VPWR VPWR _6602_/X sky130_fd_sc_hd__a22o_1
XANTENNA_14 _6111_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3814_ _7297_/Q hold12/A _5731_/B input26/X _3503_/X VGND VGND VPWR VPWR _3814_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_25 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7582_ _7582_/CLK hold38/X fanout585/X VGND VGND VPWR VPWR _7582_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_172_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_36 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4794_/A _4803_/A _5410_/B VGND VGND VPWR VPWR _4800_/A sky130_fd_sc_hd__and3_1
XANTENNA_47 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _6086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 wire346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _7354_/Q _6459_/B _6459_/C _6451_/X _7482_/Q VGND VGND VPWR VPWR _6533_/X
+ sky130_fd_sc_hd__a32o_1
X_3745_ _7370_/Q _5758_/A _4370_/A _7044_/Q VGND VGND VPWR VPWR _3745_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3771__A2 _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6464_ _7375_/Q _6408_/B _6463_/X _7423_/Q VGND VGND VPWR VPWR _6464_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3676_ _7060_/Q hold56/A _4521_/B _4322_/A _7005_/Q VGND VGND VPWR VPWR _3676_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7559__SET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5415_ _4706_/Y _4796_/Y _4802_/Y _4759_/Y _5414_/Y VGND VGND VPWR VPWR _5535_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_179_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6395_ _7050_/Q _7592_/Q _6317_/C _6072_/X _7156_/Q VGND VGND VPWR VPWR _6395_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3523__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5346_ _5094_/A _5183_/C _4942_/A _4948_/C VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__o211a_4
Xoutput176 _3435_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3425_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3415_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
Xhold2901 hold2901/A VGND VGND VPWR VPWR hold2901/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2912 hold2912/A VGND VGND VPWR VPWR hold2912/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2923 _5832_/X VGND VGND VPWR VPWR hold2923/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5277_ _5222_/A _4743_/Y _5399_/C _5387_/C VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__o211a_1
XANTENNA_fanout486_A _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2934 hold2934/A VGND VGND VPWR VPWR _4354_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2945 hold2945/A VGND VGND VPWR VPWR _4409_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5276__A2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7016_ _7211_/CLK _7016_/D fanout572/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2956 hold716/X VGND VGND VPWR VPWR _5718_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4228_ _4228_/A0 _4227_/X _4232_/S VGND VGND VPWR VPWR _4228_/X sky130_fd_sc_hd__mux2_1
Xhold2967 _7655_/A VGND VGND VPWR VPWR hold989/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2978 _7183_/Q VGND VGND VPWR VPWR hold2978/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2989 _7005_/Q VGND VGND VPWR VPWR hold722/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4159_ input1/X input2/X VGND VGND VPWR VPWR _4159_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_69_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6225__A1 _7292_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4814__A _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6528__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4533__B _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5197__D1 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_191_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1935_A _7247_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3762__A2 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input47_A mgmt_gpio_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout370 _3576_/X VGND VGND VPWR VPWR _5623_/B sky130_fd_sc_hd__buf_12
XANTENNA__4708__B _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout381 _5965_/A VGND VGND VPWR VPWR _4491_/B sky130_fd_sc_hd__buf_8
Xfanout392 hold2225/X VGND VGND VPWR VPWR _5785_/A sky130_fd_sc_hd__buf_6
XANTENNA__4427__C _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6216__A1 _7492_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6216__B2 _7444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6767__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5975__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output203_A wire365/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6519__A2 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_4
X_3530_ hold36/X _5590_/A _4509_/A VGND VGND VPWR VPWR _5857_/A sky130_fd_sc_hd__and3_4
XANTENNA__3753__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_2
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _4168_/D sky130_fd_sc_hd__buf_12
Xhold807 hold807/A VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_2
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_4
Xhold818 hold818/A VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold829 hold829/A VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3461_ _3460_/X _3461_/A1 _4429_/B VGND VGND VPWR VPWR _3461_/X sky130_fd_sc_hd__mux2_1
Xmax_cap537 _5282_/D VGND VGND VPWR VPWR _5118_/C sky130_fd_sc_hd__buf_2
Xmax_cap548 _4702_/Y VGND VGND VPWR VPWR _5118_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6089__C _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5200_ _5200_/A _5200_/B _5200_/C VGND VGND VPWR VPWR _5202_/A sky130_fd_sc_hd__and3_1
XANTENNA__3506__C _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6180_ _7466_/Q _6121_/A _6116_/A _6379_/B1 _7522_/Q VGND VGND VPWR VPWR _6180_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2208 _7310_/Q VGND VGND VPWR VPWR hold514/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5131_ _4703_/Y _5451_/A1 _4716_/Y _5028_/C VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__o31a_1
Xhold2219 hold522/X VGND VGND VPWR VPWR _5667_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2416_A _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5062_ _4605_/Y _4654_/Y _4880_/Y _4846_/Y _4744_/Y VGND VGND VPWR VPWR _5064_/B
+ sky130_fd_sc_hd__o32a_1
Xhold1507 hold1507/A VGND VGND VPWR VPWR _5982_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1518 hold184/X VGND VGND VPWR VPWR _7513_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1529 _7532_/Q VGND VGND VPWR VPWR hold211/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4013_ _6892_/Q _6891_/Q _3401_/Y _4062_/A _4011_/X VGND VGND VPWR VPWR _4014_/B
+ sky130_fd_sc_hd__o311ai_4
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6833__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6758__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5964_ _5964_/A0 _5991_/A1 _5964_/S VGND VGND VPWR VPWR _5964_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4915_ _5213_/B _5260_/D _4915_/C VGND VGND VPWR VPWR _4916_/B sky130_fd_sc_hd__and3_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5895_ _5985_/A1 _5895_/A1 _5901_/S VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5718__A0 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7634_ _7636_/CLK _7634_/D VGND VGND VPWR VPWR _7634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4846_ _5107_/A _4846_/B VGND VGND VPWR VPWR _4846_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__3992__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6391__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7565_ _7565_/CLK hold73/X fanout603/X VGND VGND VPWR VPWR _7565_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4777_ _4733_/A _4733_/B _4641_/B _4768_/Y VGND VGND VPWR VPWR _4777_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_16_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6516_ _7545_/Q _6419_/A _6512_/X _6515_/X VGND VGND VPWR VPWR _6516_/X sky130_fd_sc_hd__a211o_4
X_3728_ _7141_/Q _4491_/B _4521_/B hold72/A _7563_/Q VGND VGND VPWR VPWR _3728_/X
+ sky130_fd_sc_hd__a32o_1
X_7496_ _7496_/CLK _7496_/D fanout586/X VGND VGND VPWR VPWR _7496_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6447_ _6455_/B _6574_/B _6447_/C VGND VGND VPWR VPWR _6447_/X sky130_fd_sc_hd__and3_4
X_3659_ _4449_/B _4388_/B _4346_/C VGND VGND VPWR VPWR _3659_/X sky130_fd_sc_hd__and3_2
XFILLER_0_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6694__B2 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6378_ _6377_/X _6376_/Y _6069_/X _6378_/B2 VGND VGND VPWR VPWR _7613_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5329_ _5011_/B _5183_/C _5260_/D _4861_/X _5183_/A VGND VGND VPWR VPWR _5329_/X
+ sky130_fd_sc_hd__o311a_2
Xhold2720 _7201_/Q VGND VGND VPWR VPWR hold823/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5249__A2 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2731 _6966_/Q VGND VGND VPWR VPWR hold848/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2742 hold2742/A VGND VGND VPWR VPWR _5687_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2753 _7652_/A VGND VGND VPWR VPWR hold2753/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2764 hold2764/A VGND VGND VPWR VPWR hold2764/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6446__D _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2775 hold2775/A VGND VGND VPWR VPWR _4522_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2786 _6995_/Q VGND VGND VPWR VPWR _4313_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2797 hold2797/A VGND VGND VPWR VPWR hold2797/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3680__A1 _7363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6462__C _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input101_A wb_adr_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5421__A2 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5709__A0 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3983__A2 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6382__B1 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6134__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4160__A2 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3623__A _3623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6437__B2 _7463_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5260__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4215__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7514__RESET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4700_ _4887_/B _5399_/B VGND VGND VPWR VPWR _4700_/Y sky130_fd_sc_hd__nand2b_4
XANTENNA__4604__D _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5680_ _5680_/A0 _5896_/A0 _5685_/S VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4631_ _4570_/Y _5301_/A1 _4740_/D VGND VGND VPWR VPWR _4631_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5176__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6373__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7350_ _7412_/CLK _7350_/D fanout581/X VGND VGND VPWR VPWR _7350_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3726__A2 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4562_ _4562_/A _4562_/B _4562_/C _4562_/D VGND VGND VPWR VPWR _4562_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_69_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6301_ _7046_/Q _6332_/B _6317_/C _6072_/X _7152_/Q VGND VGND VPWR VPWR _6301_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold604 hold604/A VGND VGND VPWR VPWR hold604/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold615 _5930_/X VGND VGND VPWR VPWR _7519_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3513_ _7574_/Q _5983_/A _5965_/A _5686_/A _7310_/Q VGND VGND VPWR VPWR _3513_/X
+ sky130_fd_sc_hd__a32o_1
Xhold626 hold626/A VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7281_ _7359_/CLK _7281_/D fanout576/X VGND VGND VPWR VPWR _7281_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6125__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4493_ _4493_/A0 _5940_/A1 _4496_/S VGND VGND VPWR VPWR _4493_/X sky130_fd_sc_hd__mux2_1
Xhold637 hold637/A VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2533_A _7158_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold648 hold648/A VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold659 hold659/A VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6232_ _7436_/Q _6110_/X _6116_/X _7316_/Q VGND VGND VPWR VPWR _6232_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3444_ _6332_/B VGND VGND VPWR VPWR _3444_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_21_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _7449_/Q _6081_/X _6089_/X _7505_/Q _6162_/X VGND VGND VPWR VPWR _6163_/X
+ sky130_fd_sc_hd__a221o_2
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 _7537_/Q VGND VGND VPWR VPWR hold551/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 hold430/X VGND VGND VPWR VPWR _5825_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2027 hold608/X VGND VGND VPWR VPWR _4488_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2038 _4181_/X VGND VGND VPWR VPWR hold463/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5118_/A _5399_/C _5113_/B _5113_/X VGND VGND VPWR VPWR _5559_/A sky130_fd_sc_hd__a31o_1
Xhold1304 hold3157/X VGND VGND VPWR VPWR hold3158/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6094_/A _6112_/D _6119_/B _6116_/C VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__and4_4
Xhold2049 hold490/X VGND VGND VPWR VPWR _4483_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 hold3164/X VGND VGND VPWR VPWR hold3165/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _4304_/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1337 _4287_/A1 VGND VGND VPWR VPWR hold2785/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5045_ _5339_/D _5183_/C _5203_/B VGND VGND VPWR VPWR _5046_/B sky130_fd_sc_hd__nand3_1
Xhold1348 _4283_/B VGND VGND VPWR VPWR hold2828/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1359 _6791_/A1 VGND VGND VPWR VPWR hold2869/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4364__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6996_ _6999_/CLK _6996_/D VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5947_ _5947_/A _5947_/B hold47/X VGND VGND VPWR VPWR _5955_/S sky130_fd_sc_hd__and3_4
XANTENNA__7255__RESET_B fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5894__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6796__B1_N _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3965__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5878_ _5878_/A0 _5896_/A0 _5883_/S VGND VGND VPWR VPWR _5878_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7617_ _7621_/CLK _7617_/D fanout576/X VGND VGND VPWR VPWR _7617_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6364__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4829_ _5094_/A _5399_/C _5113_/B VGND VGND VPWR VPWR _4830_/B sky130_fd_sc_hd__and3_1
XFILLER_0_173_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7548_ _7556_/CLK _7548_/D fanout597/X VGND VGND VPWR VPWR _7548_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7479_ _7566_/CLK _7479_/D fanout599/X VGND VGND VPWR VPWR _7479_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6667__A1 _7197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4539__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3240 _7208_/Q VGND VGND VPWR VPWR _5580_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6457__C _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3251 _7101_/Q VGND VGND VPWR VPWR _4114_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3262 _6894_/Q VGND VGND VPWR VPWR _4054_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3273 _7598_/Q VGND VGND VPWR VPWR _6060_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input149_A wb_dat_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3284 _6909_/Q VGND VGND VPWR VPWR _4002_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2550 _5655_/X VGND VGND VPWR VPWR hold152/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2561 _7264_/Q VGND VGND VPWR VPWR hold702/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2572 _5881_/X VGND VGND VPWR VPWR hold2572/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2583 hold813/X VGND VGND VPWR VPWR _5792_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2594 hold807/X VGND VGND VPWR VPWR _5684_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1860 _7282_/Q VGND VGND VPWR VPWR hold346/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1871 _7445_/Q VGND VGND VPWR VPWR hold122/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1882 _4548_/X VGND VGND VPWR VPWR hold449/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1893 _5638_/X VGND VGND VPWR VPWR hold349/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3956__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4721__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_163_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3708__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6107__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4118__C1 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6658__B2 _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4669__B1 _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5330__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5330__B2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4168__B _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3892__A1 _7360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3644__A1 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6850_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6850_/X sky130_fd_sc_hd__and2_1
X_5801_ _5999_/A1 _5801_/A1 _5802_/S VGND VGND VPWR VPWR _5801_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_187_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6781_ _6792_/S _6781_/B VGND VGND VPWR VPWR _6781_/Y sky130_fd_sc_hd__nand2_1
X_3993_ _6988_/Q _5731_/B _5623_/B _5704_/A _7319_/Q VGND VGND VPWR VPWR _3993_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4334__D hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5732_ _5732_/A0 _5948_/A1 _5739_/S VGND VGND VPWR VPWR _5732_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3947__A2 _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5663_ _5663_/A0 _5951_/A1 _5667_/S VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6346__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7402_ _7555_/CLK _7402_/D fanout594/X VGND VGND VPWR VPWR _7402_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_142_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4614_ _4657_/D _4657_/C _4909_/C _4909_/A VGND VGND VPWR VPWR _4614_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5594_ _5594_/A0 _5647_/A0 _5595_/S VGND VGND VPWR VPWR _5594_/X sky130_fd_sc_hd__mux2_1
Xhold401 hold401/A VGND VGND VPWR VPWR _7474_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7333_ _7333_/CLK _7333_/D fanout579/X VGND VGND VPWR VPWR _7333_/Q sky130_fd_sc_hd__dfrtp_4
X_4545_ _4545_/A _5902_/B VGND VGND VPWR VPWR _4550_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_170_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold412 hold412/A VGND VGND VPWR VPWR hold412/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold423 hold423/A VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold434 hold434/A VGND VGND VPWR VPWR hold434/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold445 hold445/A VGND VGND VPWR VPWR _7518_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3580__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7264_ _7264_/CLK _7264_/D fanout567/X VGND VGND VPWR VPWR _7264_/Q sky130_fd_sc_hd__dfrtp_1
Xhold456 hold456/A VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4476_ _4476_/A0 _5914_/A1 _4478_/S VGND VGND VPWR VPWR _4476_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6113__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold467 hold467/A VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold478 hold478/A VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold489 hold489/A VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6215_ _6214_/X _6237_/A2 _6573_/S VGND VGND VPWR VPWR _6215_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3427_ _7426_/Q VGND VGND VPWR VPWR _3427_/Y sky130_fd_sc_hd__inv_2
X_7195_ _7212_/CLK _7195_/D fanout574/X VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6649_/S _7602_/Q _4116_/X _6067_/X VGND VGND VPWR VPWR _6146_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4078__B _4078_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3883__A1 _7123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1101 _5769_/X VGND VGND VPWR VPWR _7376_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 _5742_/X VGND VGND VPWR VPWR _7352_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4509__D _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1123 hold2981/X VGND VGND VPWR VPWR hold2982/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _5795_/X VGND VGND VPWR VPWR _7399_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6077_ _7343_/Q _6070_/X _6072_/X _7415_/Q _6076_/X VGND VGND VPWR VPWR _6102_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6574__A _7444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1145 hold2952/X VGND VGND VPWR VPWR hold2953/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout566_A fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 hold1156/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
XANTENNA__6821__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1167 hold2819/X VGND VGND VPWR VPWR hold2820/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5028_ _5028_/A _5028_/B _5028_/C VGND VGND VPWR VPWR _5031_/C sky130_fd_sc_hd__nand3_1
Xhold1178 hold1178/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
XANTENNA__3635__A1 _7492_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 hold2816/X VGND VGND VPWR VPWR hold2817/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3635__B2 _7468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_71_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6585__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6979_ _7636_/CLK _6979_/D VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3938__A2 _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6337__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1750_A _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6468__B _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5312__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold990 hold990/A VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3070 hold3070/A VGND VGND VPWR VPWR _4401_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5799__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3081 hold3081/A VGND VGND VPWR VPWR hold3081/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3092 _4546_/X VGND VGND VPWR VPWR hold3092/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2380 _5883_/X VGND VGND VPWR VPWR hold607/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6812__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2391 _7019_/Q VGND VGND VPWR VPWR hold915/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7177__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3626__B2 _7324_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1690 hold78/X VGND VGND VPWR VPWR _4438_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4969__A4 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7106__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5379__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6576__B1 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4732__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4330_ _4330_/A0 _5805_/A1 _4333_/S VGND VGND VPWR VPWR _4330_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4261_ _4261_/A0 _5805_/A1 _4264_/S VGND VGND VPWR VPWR _4261_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6500__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6097__C _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6000_ _6000_/A0 hold17/X hold37/X VGND VGND VPWR VPWR _6000_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4192_ _4192_/A0 _5948_/A1 _4202_/S VGND VGND VPWR VPWR _4192_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6803__A1 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3530__B _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6902_ _4150_/A1 _6902_/D _6852_/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6833_ _6833_/A _6839_/B VGND VGND VPWR VPWR _6833_/X sky130_fd_sc_hd__and2_1
XANTENNA__6567__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6764_ _6878_/Q _6451_/X _6759_/X _6761_/X _6763_/X VGND VGND VPWR VPWR _6774_/B
+ sky130_fd_sc_hd__a2111oi_4
X_3976_ _7583_/Q _5640_/C _5623_/B _3973_/X _3975_/X VGND VGND VPWR VPWR _3988_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5385__A4 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5715_ _5967_/A1 _5715_/A1 _5721_/S VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_162_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5790__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6695_ _7138_/Q _6419_/C _6446_/X _7188_/Q VGND VGND VPWR VPWR _6695_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5646_ _5986_/A1 _5646_/A1 _5649_/S VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5577_ _5533_/Y _5569_/X _5576_/X VGND VGND VPWR VPWR _5577_/Y sky130_fd_sc_hd__o21ai_1
Xhold220 hold220/A VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7316_ _7478_/CLK _7316_/D fanout580/X VGND VGND VPWR VPWR _7316_/Q sky130_fd_sc_hd__dfrtp_4
Xhold231 hold231/A VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4528_ _4528_/A0 _5714_/A0 _4532_/S VGND VGND VPWR VPWR _4528_/X sky130_fd_sc_hd__mux2_1
Xhold242 hold242/A VGND VGND VPWR VPWR _7498_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold253 hold253/A VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold264 hold264/A VGND VGND VPWR VPWR _7385_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6098__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold275 hold275/A VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7247_ _7333_/CLK _7247_/D fanout582/X VGND VGND VPWR VPWR _7247_/Q sky130_fd_sc_hd__dfrtp_4
X_4459_ _4459_/A0 _5852_/A0 _4460_/S VGND VGND VPWR VPWR _4459_/X sky130_fd_sc_hd__mux2_1
Xhold286 hold286/A VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold297 hold297/A VGND VGND VPWR VPWR _7562_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7178_ _7178_/CLK _7178_/D fanout606/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _7448_/Q _6144_/A _6116_/A _6379_/B1 _7520_/Q VGND VGND VPWR VPWR _6129_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__A _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__A1 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7270__RESET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6270__A2 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6558__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5230__B1 _5102_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4271__B _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4702__D _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6325__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input77_A ser_tx VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6730__B1 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3847__A1 _7246_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5830__B _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6645__C _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7333_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6261__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6100__A_N _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4272__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6549__B1 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _6964_/Q _5603_/B _5640_/C _3829_/X VGND VGND VPWR VPWR _3830_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_68_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7537_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3761_ input6/X _5983_/A _5612_/B _3542_/X _6922_/Q VGND VGND VPWR VPWR _3761_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5772__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5500_ _5053_/C _5329_/X _5426_/X _5203_/B _5171_/X VGND VGND VPWR VPWR _5501_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_172_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3783__B1 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6480_ _7432_/Q _6747_/B _6645_/C _6421_/X _7320_/Q VGND VGND VPWR VPWR _6480_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4980__C1 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3692_ _7055_/Q _5866_/B _5619_/B _3649_/X _7070_/Q VGND VGND VPWR VPWR _3692_/X
+ sky130_fd_sc_hd__a32o_1
X_5431_ _5342_/B _4956_/Y _5180_/A _5553_/A1 VGND VGND VPWR VPWR _5499_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_30_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5524__A1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6721__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput303 _3578_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
Xoutput314 hold1183/X VGND VGND VPWR VPWR hold1184/A sky130_fd_sc_hd__buf_6
XANTENNA_hold2446_A _7393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5362_ _4954_/C _4929_/A _5346_/X _5233_/X VGND VGND VPWR VPWR _5510_/A sky130_fd_sc_hd__a31oi_2
Xoutput325 hold1155/X VGND VGND VPWR VPWR hold1156/A sky130_fd_sc_hd__buf_6
XANTENNA__4842__A_N _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput336 hold1201/X VGND VGND VPWR VPWR hold1202/A sky130_fd_sc_hd__buf_6
X_7101_ _7644_/CLK _7101_/D _4309_/B VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfstp_2
X_4313_ _4321_/S _4313_/B VGND VGND VPWR VPWR _4313_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3525__B _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5293_ _5168_/X _5206_/Y _5292_/Y _4428_/Y hold19/A VGND VGND VPWR VPWR _7203_/D
+ sky130_fd_sc_hd__o32a_1
X_7032_ _7112_/CLK _7032_/D fanout589/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_4
X_4244_ _5656_/A1 _5953_/A1 _4248_/S VGND VGND VPWR VPWR _4244_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3838__A1 _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6836__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3838__B2 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4175_ _4175_/A input1/X VGND VGND VPWR VPWR _4175_/X sky130_fd_sc_hd__and2_1
XANTENNA__3541__A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6252__A2 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7519__SET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6852__A _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4263__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6816_ _6815_/X _6816_/A1 _6822_/S VGND VGND VPWR VPWR _7642_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout431_A _6429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6555__A3 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6747_ _7175_/Q _6747_/B _6747_/C VGND VGND VPWR VPWR _6747_/X sky130_fd_sc_hd__and3_1
XFILLER_0_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3959_ _7503_/Q _5911_/A _3496_/Y _3955_/X _3958_/X VGND VGND VPWR VPWR _3959_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_758 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6678_ _7037_/Q _6459_/B _6651_/C _6423_/X _7012_/Q VGND VGND VPWR VPWR _6678_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5629_ _5629_/A0 _5805_/A1 _5629_/S VGND VGND VPWR VPWR _5629_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6712__B1 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout552 _5401_/A3 VGND VGND VPWR VPWR _5107_/A sky130_fd_sc_hd__clkbuf_16
Xfanout563 _4128_/B VGND VGND VPWR VPWR _6865_/A sky130_fd_sc_hd__buf_8
XANTENNA__6491__A2 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout574 fanout587/X VGND VGND VPWR VPWR fanout574/X sky130_fd_sc_hd__buf_8
Xfanout585 fanout586/X VGND VGND VPWR VPWR fanout585/X sky130_fd_sc_hd__clkbuf_16
Xfanout596 fanout597/X VGND VGND VPWR VPWR fanout596/X sky130_fd_sc_hd__buf_12
XANTENNA_input131_A wb_cyc_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6243__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_9__f_wb_clk_i clkbuf_3_4_0_wb_clk_i/X VGND VGND VPWR VPWR _7206_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4254__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5754__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3765__B1 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6701__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6703__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3517__B1 hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4221__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6909__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6482__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5690__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4493__A1 _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4176__B _4176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6094__D _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5980_ _5998_/A1 _5980_/A1 _5982_/S VGND VGND VPWR VPWR _5980_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4931_ _5183_/C _4933_/A _4933_/B VGND VGND VPWR VPWR _4934_/A sky130_fd_sc_hd__and3_1
XANTENNA__3599__A3 _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5993__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7650_ _7650_/A VGND VGND VPWR VPWR _7650_/X sky130_fd_sc_hd__clkbuf_2
X_4862_ _4984_/B _4574_/X _4797_/B _4669_/X _4974_/B VGND VGND VPWR VPWR _4862_/X
+ sky130_fd_sc_hd__a311o_2
XANTENNA__4623__C _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6601_ _7517_/Q _6435_/X _6446_/X _7525_/Q VGND VGND VPWR VPWR _6601_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_28_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3813_ _7473_/Q _4509_/A _5947_/A _3617_/X _7231_/Q VGND VGND VPWR VPWR _3813_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_15 _6516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7581_ _7581_/CLK _7581_/D fanout584/X VGND VGND VPWR VPWR _7581_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5745__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4793_ _4794_/A _5410_/B VGND VGND VPWR VPWR _4793_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_37 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_48 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6532_ _7290_/Q _6422_/X _6443_/X _7450_/Q _6531_/X VGND VGND VPWR VPWR _6532_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__3756__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_59 _6212_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3744_ _7546_/Q _5992_/C _4212_/A _3741_/X _3743_/X VGND VGND VPWR VPWR _3744_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_82_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6463_ _6463_/A _6600_/B _6747_/C VGND VGND VPWR VPWR _6463_/X sky130_fd_sc_hd__and3_4
X_3675_ hold36/A _5612_/C hold56/A VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__and3_4
XFILLER_0_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5414_ _5113_/A _5295_/C _5404_/C _4802_/A _5410_/A VGND VGND VPWR VPWR _5414_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_179_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6394_ _7055_/Q _6087_/X _6119_/X _7136_/Q _6393_/X VGND VGND VPWR VPWR _6397_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4181__A0 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5345_ _5343_/Y _5506_/C _4969_/Y VGND VGND VPWR VPWR _5345_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput177 _3434_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3424_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
Xhold2902 _7122_/Q VGND VGND VPWR VPWR hold2902/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xoutput199 _3414_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
Xhold2913 _7634_/Q VGND VGND VPWR VPWR _6790_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5276_ _5563_/A1 _4709_/Y _4814_/Y _5102_/Y VGND VGND VPWR VPWR _5278_/B sky130_fd_sc_hd__o31a_1
Xhold2924 _6976_/Q VGND VGND VPWR VPWR _4285_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2935 _7210_/Q VGND VGND VPWR VPWR hold2935/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7015_ _7070_/CLK _7015_/D fanout590/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2946 _4409_/X VGND VGND VPWR VPWR hold2946/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6473__A2 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4227_ _4256_/A0 _4256_/A1 _4231_/S VGND VGND VPWR VPWR _4227_/X sky130_fd_sc_hd__mux2_1
Xhold2957 _7511_/Q VGND VGND VPWR VPWR hold2957/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout381_A _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4484__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2968 hold989/X VGND VGND VPWR VPWR _4226_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout479_A _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2979 hold2979/A VGND VGND VPWR VPWR _4535_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4158_ _7257_/Q _7306_/Q _4168_/D _6881_/Q _4157_/Y VGND VGND VPWR VPWR _4158_/X
+ sky130_fd_sc_hd__o41a_2
XANTENNA__5897__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6225__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4089_ input118/X input119/X _4089_/C _4089_/D VGND VGND VPWR VPWR _4093_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__4236__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5984__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4888__A_N _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5736__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_191_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1830_A _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6464__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5121__C1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout360 _5453_/A VGND VGND VPWR VPWR _5213_/B sky130_fd_sc_hd__buf_12
XANTENNA__5672__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout371 _3576_/X VGND VGND VPWR VPWR _4521_/B sky130_fd_sc_hd__buf_8
XANTENNA__4475__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout382 _5614_/B VGND VGND VPWR VPWR _5965_/A sky130_fd_sc_hd__buf_8
XANTENNA__4708__C _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4427__D _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4227__A1 _4256_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5424__B1 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6767__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5727__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_4
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3753__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _4173_/A sky130_fd_sc_hd__buf_4
Xhold808 _5684_/X VGND VGND VPWR VPWR _7301_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput79 spi_enabled VGND VGND VPWR VPWR _4174_/B sky130_fd_sc_hd__buf_6
Xhold819 hold819/A VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_150_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6152__A1 _7481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3460_ hold396/X _6902_/Q _4025_/A VGND VGND VPWR VPWR _3460_/X sky130_fd_sc_hd__mux2_2
Xmax_cap549 _4702_/Y VGND VGND VPWR VPWR _4810_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5130_ _4703_/Y _4707_/Y _4783_/Y _4956_/A VGND VGND VPWR VPWR _5150_/A sky130_fd_sc_hd__o22a_1
Xhold2209 hold514/X VGND VGND VPWR VPWR _5694_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5061_ _5107_/A _5061_/B _5399_/D VGND VGND VPWR VPWR _5061_/X sky130_fd_sc_hd__and3_1
Xhold1508 _5982_/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1519 _7095_/Q VGND VGND VPWR VPWR hold217/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4466__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4012_ _6892_/Q _6891_/Q VGND VGND VPWR VPWR _4123_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5963_ _5963_/A0 hold61/X _5964_/S VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5966__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4914_ _5213_/B _5183_/C _4929_/A _4940_/D VGND VGND VPWR VPWR _4916_/A sky130_fd_sc_hd__and4_1
XFILLER_0_48_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5894_ _5993_/A1 _5894_/A1 _5901_/S VGND VGND VPWR VPWR _5894_/X sky130_fd_sc_hd__mux2_1
X_7633_ _7633_/CLK _7633_/D VGND VGND VPWR VPWR _7633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4845_ _5115_/A _5115_/B _5107_/A VGND VGND VPWR VPWR _4845_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7564_ _7566_/CLK _7564_/D fanout603/X VGND VGND VPWR VPWR _7564_/Q sky130_fd_sc_hd__dfrtp_4
X_4776_ _4776_/A _4776_/B VGND VGND VPWR VPWR _4776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_99_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6515_ _7561_/Q _6419_/C _6443_/X _7449_/Q _6514_/X VGND VGND VPWR VPWR _6515_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3727_ _7315_/Q _3521_/X _3723_/X _3724_/X _3726_/X VGND VGND VPWR VPWR _3727_/X
+ sky130_fd_sc_hd__a2111o_4
X_7495_ _7537_/CLK _7495_/D fanout577/X VGND VGND VPWR VPWR _7495_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3744__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6446_ _6462_/D _7595_/Q _6463_/A _6600_/B VGND VGND VPWR VPWR _6446_/X sky130_fd_sc_hd__and4_4
XANTENNA__6143__A1 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3658_ _4473_/A _5830_/C _4388_/B VGND VGND VPWR VPWR _3658_/X sky130_fd_sc_hd__and3_2
XFILLER_0_141_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6694__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6377_ _6751_/S _7612_/Q _4116_/X _6067_/X VGND VGND VPWR VPWR _6377_/X sky130_fd_sc_hd__o2bb2a_1
X_3589_ _7581_/Q _3501_/X _5776_/A _7389_/Q _3588_/X VGND VGND VPWR VPWR _3589_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout596_A fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5328_ _5328_/A _5328_/B _5339_/B VGND VGND VPWR VPWR _5328_/X sky130_fd_sc_hd__and3_2
Xhold2710 _7166_/Q VGND VGND VPWR VPWR hold833/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2721 hold823/X VGND VGND VPWR VPWR _4556_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2732 hold848/X VGND VGND VPWR VPWR _4270_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5259_ _4605_/Y _5451_/A1 _4744_/Y _5072_/Y VGND VGND VPWR VPWR _5265_/A sky130_fd_sc_hd__o31a_1
XANTENNA__4457__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5654__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2743 _7359_/Q VGND VGND VPWR VPWR hold2743/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2754 hold2754/A VGND VGND VPWR VPWR _4245_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2765 _7050_/Q VGND VGND VPWR VPWR hold856/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2776 _4522_/X VGND VGND VPWR VPWR hold2776/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2787 hold2787/A VGND VGND VPWR VPWR hold2787/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2798 _7112_/Q VGND VGND VPWR VPWR hold2798/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4209__A1 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5406__B1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3680__A2 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5957__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3968__B1 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5421__A3 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6382__A1 _7116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4393__A0 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3259_A _7628_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6134__A1 _7360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6134__B2 _7392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_csclk_A _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6685__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3499__A2 _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6437__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4448__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5645__A0 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5948__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4630_ _4570_/Y _5301_/A1 _4627_/Y VGND VGND VPWR VPWR _4767_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5176__A2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6373__A1 _7145_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4384__A0 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4561_ _4562_/A _4562_/B _4562_/C _4562_/D VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__and4_4
X_6300_ _7006_/Q _6082_/X _6111_/X _7036_/Q _6299_/X VGND VGND VPWR VPWR _6303_/C
+ sky130_fd_sc_hd__a221o_1
X_3512_ _5722_/A _4449_/B _5731_/B VGND VGND VPWR VPWR _5686_/A sky130_fd_sc_hd__and3_4
XANTENNA_hold2359_A _7339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7280_ _7309_/CLK _7280_/D fanout576/X VGND VGND VPWR VPWR _7280_/Q sky130_fd_sc_hd__dfstp_2
Xhold605 _5697_/X VGND VGND VPWR VPWR _7312_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6125__A1 _7464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6125__B2 _7352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4492_ _4492_/A0 _5840_/A1 _4496_/S VGND VGND VPWR VPWR _4492_/X sky130_fd_sc_hd__mux2_1
Xhold616 hold616/A VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold627 _5648_/X VGND VGND VPWR VPWR _7269_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold638 _5781_/X VGND VGND VPWR VPWR _7387_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold649 hold649/A VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6231_ _7404_/Q _6091_/X _6116_/B _7356_/Q _6099_/X VGND VGND VPWR VPWR _6231_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_hold48_A hold48/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5479__A3 _4971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _7521_/Q _6112_/D _6119_/B _6136_/B _6144_/C VGND VGND VPWR VPWR _6162_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 hold551/X VGND VGND VPWR VPWR _5950_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2017 _5825_/X VGND VGND VPWR VPWR hold431/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5113_ _5113_/A _5113_/B _5282_/D VGND VGND VPWR VPWR _5113_/X sky130_fd_sc_hd__and3_1
Xhold2028 _4488_/X VGND VGND VPWR VPWR hold609/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2039 hold463/X VGND VGND VPWR VPWR hold2039/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _7588_/Q _6106_/B _6119_/A _7589_/Q VGND VGND VPWR VPWR _6093_/X sky130_fd_sc_hd__and4bb_4
Xhold1305 hold3130/X VGND VGND VPWR VPWR hold3131/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4439__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 _5732_/X VGND VGND VPWR VPWR _7343_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_85_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1327 hold3106/X VGND VGND VPWR VPWR hold3107/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5044_/B _5044_/C VGND VGND VPWR VPWR _5047_/C sky130_fd_sc_hd__nand3_1
Xhold1338 _4312_/A1 VGND VGND VPWR VPWR hold2796/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1349 _4296_/B VGND VGND VPWR VPWR hold2838/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5939__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4364__B _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6995_ _6999_/CLK _6995_/D VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5946_ _5946_/A0 hold17/X hold23/X VGND VGND VPWR VPWR _5946_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4611__A1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5877_ _5877_/A0 _5967_/A1 _5883_/S VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3965__A3 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7616_ _7621_/CLK _7616_/D fanout576/X VGND VGND VPWR VPWR _7616_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout511_A _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4828_ _5399_/C _5118_/B VGND VGND VPWR VPWR _4828_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_118_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4375__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4759_ _5158_/A _5183_/A VGND VGND VPWR VPWR _4759_/Y sky130_fd_sc_hd__nand2_8
X_7547_ _7555_/CLK _7547_/D fanout597/X VGND VGND VPWR VPWR _7547_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_133_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1459_A _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7478_ _7478_/CLK _7478_/D fanout581/X VGND VGND VPWR VPWR _7478_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4127__A0 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6667__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6429_ _6435_/B _6462_/D _7593_/Q _7594_/Q VGND VGND VPWR VPWR _6429_/X sky130_fd_sc_hd__and4b_4
XFILLER_0_101_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3230 _7105_/Q VGND VGND VPWR VPWR _6827_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4539__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3241 _7627_/Q VGND VGND VPWR VPWR _6777_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3252 _7107_/Q VGND VGND VPWR VPWR _4427_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3263 _6891_/Q VGND VGND VPWR VPWR _4064_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3274 _6908_/Q VGND VGND VPWR VPWR _4005_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2540 hold704/X VGND VGND VPWR VPWR _4529_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3285 _7257_/Q VGND VGND VPWR VPWR _4250_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2551 _7581_/Q VGND VGND VPWR VPWR hold827/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2562 hold702/X VGND VGND VPWR VPWR _5642_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2573 _7285_/Q VGND VGND VPWR VPWR hold839/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2584 _6922_/Q VGND VGND VPWR VPWR hold967/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_188_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2595 _7416_/Q VGND VGND VPWR VPWR hold769/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1850 _4367_/X VGND VGND VPWR VPWR hold507/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1861 hold346/X VGND VGND VPWR VPWR _5663_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1872 hold122/X VGND VGND VPWR VPWR _5846_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1883 _7449_/Q VGND VGND VPWR VPWR hold310/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_168_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1894 _7378_/Q VGND VGND VPWR VPWR hold328/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_94_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3708__A3 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6107__B2 _7391_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6658__A2 _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4669__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5330__A2 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__B _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3892__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4168__C _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__buf_8
XFILLER_0_176_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6291__B1 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5995__S hold37/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5800_ _5953_/A1 _5800_/A1 _5802_/S VGND VGND VPWR VPWR _5800_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6780_ _7102_/Q _6780_/B VGND VGND VPWR VPWR _6792_/S sky130_fd_sc_hd__nand2_8
XANTENNA__6594__A1 _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3992_ _7367_/Q _5758_/A _5634_/A _7262_/Q _3991_/X VGND VGND VPWR VPWR _3992_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_187_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5731_ _5947_/A _5731_/B hold47/X VGND VGND VPWR VPWR _5739_/S sky130_fd_sc_hd__and3_4
XFILLER_0_45_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3947__A3 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5662_ _5662_/A0 _5896_/A0 _5667_/S VGND VGND VPWR VPWR _5662_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6346__B2 _7184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4613_ _4909_/A _4909_/C VGND VGND VPWR VPWR _4657_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_170_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7401_ _7476_/CLK _7401_/D fanout586/X VGND VGND VPWR VPWR _7401_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5593_ _5593_/A0 _5950_/A1 _5595_/S VGND VGND VPWR VPWR _5593_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7332_ _7366_/CLK _7332_/D fanout579/X VGND VGND VPWR VPWR _7332_/Q sky130_fd_sc_hd__dfrtp_4
X_4544_ _4544_/A0 _5754_/A1 hold57/X VGND VGND VPWR VPWR _4544_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold402 hold402/A VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6839__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold413 hold413/A VGND VGND VPWR VPWR _7457_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold424 hold424/A VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3580__B2 _6925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7263_ _7264_/CLK _7263_/D fanout569/X VGND VGND VPWR VPWR _7263_/Q sky130_fd_sc_hd__dfrtp_1
Xhold435 hold435/A VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold446 hold446/A VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4475_ _4475_/A0 _5583_/A0 _4478_/S VGND VGND VPWR VPWR _4475_/X sky130_fd_sc_hd__mux2_1
Xhold457 hold457/A VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3544__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold468 hold468/A VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_187_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6214_ _6213_/Y _6212_/Y _7605_/Q _6649_/S VGND VGND VPWR VPWR _6214_/X sky130_fd_sc_hd__a2bb2o_1
X_3426_ _7434_/Q VGND VGND VPWR VPWR _3426_/Y sky130_fd_sc_hd__inv_2
Xhold479 hold479/A VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7194_ _7211_/CLK _7194_/D fanout574/X VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5321__A2 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6145_ _6036_/Y _7280_/Q _6143_/X _6133_/X _6775_/B1 VGND VGND VPWR VPWR _6145_/Y
+ sky130_fd_sc_hd__o221ai_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6855__A _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4078__C _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3883__A2 _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 hold2857/X VGND VGND VPWR VPWR hold2858/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 hold2935/X VGND VGND VPWR VPWR hold2936/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 hold2983/X VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6076_ _7511_/Q _6110_/A _6317_/C _6075_/X _7423_/Q VGND VGND VPWR VPWR _6076_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6574__B _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1135 hold3006/X VGND VGND VPWR VPWR hold3007/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1146 hold2954/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5085__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6282__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1157 hold2850/X VGND VGND VPWR VPWR hold2851/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5027_ _5183_/A _5295_/C _5038_/B _5339_/C VGND VGND VPWR VPWR _5028_/B sky130_fd_sc_hd__nand4_1
Xhold1168 hold1168/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
Xhold1179 hold2863/X VGND VGND VPWR VPWR hold1179/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3635__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6585__A1 _7316_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6978_ _7636_/CLK _6978_/D VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3938__A3 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5929_ _5929_/A _5992_/D VGND VGND VPWR VPWR _5937_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6337__B2 _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4899__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6468__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input161_A wb_dat_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold980 hold980/A VGND VGND VPWR VPWR _7420_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold991 hold991/A VGND VGND VPWR VPWR hold991/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3060 hold3060/A VGND VGND VPWR VPWR _4235_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3874__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3071 _7248_/Q VGND VGND VPWR VPWR hold3071/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3082 _7527_/Q VGND VGND VPWR VPWR hold3082/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3093 _7487_/Q VGND VGND VPWR VPWR hold3093/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2370 hold929/X VGND VGND VPWR VPWR _5953_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input22_A mask_rev_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2381 _7380_/Q VGND VGND VPWR VPWR hold995/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2392 hold915/X VGND VGND VPWR VPWR _4344_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4285__A _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3626__A2 _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1680 _7436_/Q VGND VGND VPWR VPWR hold251/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1691 _4438_/X VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5379__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_168_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6733__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4260_ _4260_/A0 _5948_/A1 _4264_/S VGND VGND VPWR VPWR _4260_/X sky130_fd_sc_hd__mux2_1
X_4191_ _5619_/A _5947_/A _5640_/D VGND VGND VPWR VPWR _4202_/S sky130_fd_sc_hd__and3_4
XFILLER_0_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6264__B1 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3530__C _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6901_ _4150_/A1 _6901_/D _6851_/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6832_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6832_/X sky130_fd_sc_hd__and2_1
XFILLER_0_187_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6567__A1 _7499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6567__B2 _7459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3975_ _7407_/Q _3493_/X _4322_/A _7001_/Q _3974_/X VGND VGND VPWR VPWR _3975_/X
+ sky130_fd_sc_hd__a221o_1
X_6763_ _7151_/Q _6408_/A _6435_/X _7050_/Q _6762_/X VGND VGND VPWR VPWR _6763_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5714_ _5714_/A0 _5714_/A1 _5721_/S VGND VGND VPWR VPWR _5714_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6319__A1 _7183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6694_ _7047_/Q _6435_/X _6452_/X _7022_/Q _6693_/X VGND VGND VPWR VPWR _6697_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5645_ _5805_/A1 _5645_/A1 _5649_/S VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5576_ _5543_/X _5575_/Y _5550_/Y _5572_/X VGND VGND VPWR VPWR _5576_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5542__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold210 hold210/A VGND VGND VPWR VPWR _7564_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold221 hold221/A VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7315_ _7478_/CLK _7315_/D fanout583/X VGND VGND VPWR VPWR _7315_/Q sky130_fd_sc_hd__dfrtp_4
X_4527_ hold56/X _5619_/B _5640_/D VGND VGND VPWR VPWR _4532_/S sky130_fd_sc_hd__and3_4
XFILLER_0_130_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold232 _5888_/X VGND VGND VPWR VPWR _7482_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold243 hold243/A VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold254 hold254/A VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold265 hold265/A VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6098__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4458_ _4458_/A0 _5914_/A1 _4460_/S VGND VGND VPWR VPWR _4458_/X sky130_fd_sc_hd__mux2_1
Xhold276 hold276/A VGND VGND VPWR VPWR _7497_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7246_ _7366_/CLK _7246_/D fanout579/X VGND VGND VPWR VPWR _7246_/Q sky130_fd_sc_hd__dfrtp_4
Xhold287 hold287/A VGND VGND VPWR VPWR _7274_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold298 hold298/A VGND VGND VPWR VPWR hold298/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4502__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3409_ _7256_/Q VGND VGND VPWR VPWR _3409_/Y sky130_fd_sc_hd__inv_2
X_7177_ _7268_/CLK _7177_/D _6871_/A VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_4
X_4389_ _5714_/A0 _4389_/A1 _4393_/S VGND VGND VPWR VPWR _4389_/X sky130_fd_sc_hd__mux2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _7424_/Q _6075_/X _6121_/X _7304_/Q _6127_/X VGND VGND VPWR VPWR _6128_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6255__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6050_/Y _7598_/Q _6427_/A _6058_/X VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_4_8__f_wb_clk_i clkbuf_3_4_0_wb_clk_i/X VGND VGND VPWR VPWR _7633_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5929__A _5929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6558__A1 _7443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3847__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5830__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6246__B1 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4219__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6797__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6797__B2 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6214__A2_N _6212_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5839__A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4743__A _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3760_ _6991_/Q _4346_/C _5623_/B _3667_/X _7024_/Q VGND VGND VPWR VPWR _3760_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_172_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3691_ _7299_/Q hold12/A _3669_/C _5794_/A _7403_/Q VGND VGND VPWR VPWR _3691_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_171_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5430_ _5429_/X _5216_/X _5339_/A VGND VGND VPWR VPWR _5554_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput304 _4167_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
X_5361_ _5361_/A _5361_/B _5573_/B _5444_/A VGND VGND VPWR VPWR _5363_/B sky130_fd_sc_hd__and4_1
Xoutput315 hold1205/X VGND VGND VPWR VPWR hold1206/A sky130_fd_sc_hd__buf_6
XFILLER_0_112_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput326 hold2764/X VGND VGND VPWR VPWR hold1154/A sky130_fd_sc_hd__buf_6
Xoutput337 hold2851/X VGND VGND VPWR VPWR hold1158/A sky130_fd_sc_hd__buf_6
X_7100_ _7521_/CLK _7100_/D fanout600/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_1
X_4312_ _3922_/Y _4312_/A1 _4321_/S VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3525__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5292_ _4969_/Y _5506_/B _5288_/Y _4428_/Y _5290_/X VGND VGND VPWR VPWR _5292_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_10_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7031_ _7112_/CLK _7031_/D fanout589/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_4
X_4243_ _4243_/A0 _4242_/X _4249_/S VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3838__A2 _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4174_ _4174_/A _4174_/B VGND VGND VPWR VPWR _4174_/X sky130_fd_sc_hd__and2_1
XANTENNA__4637__B _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6237__B1 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3541__B _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5749__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6815_ _7110_/Q _6815_/A2 _6815_/B1 wire463/A _6814_/X VGND VGND VPWR VPWR _6815_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6746_ _7039_/Q _6459_/B _6651_/C _6463_/X _7165_/Q VGND VGND VPWR VPWR _6746_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_175_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3958_ _7519_/Q _5785_/B _3496_/Y _3957_/X VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4971__B1 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3889_ _7245_/Q _5947_/A _3519_/B _5713_/A _7328_/Q VGND VGND VPWR VPWR _3889_/X
+ sky130_fd_sc_hd__a32o_4
X_6677_ _7178_/Q _6058_/X _6409_/X _7133_/Q VGND VGND VPWR VPWR _6677_/X sky130_fd_sc_hd__a22o_1
X_5628_ _5628_/A0 _5954_/A1 _5629_/S VGND VGND VPWR VPWR _5628_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6173__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6712__B2 _7119_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5559_ _5559_/A _5559_/B _5559_/C _5559_/D VGND VGND VPWR VPWR _5560_/C sky130_fd_sc_hd__nor4_1
XFILLER_0_130_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7229_ _7255_/CLK _7229_/D _4128_/B VGND VGND VPWR VPWR _7229_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout520 _7591_/Q VGND VGND VPWR VPWR _6119_/A sky130_fd_sc_hd__buf_12
XANTENNA__4828__A _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout531 _4940_/C VGND VGND VPWR VPWR _5260_/D sky130_fd_sc_hd__buf_12
XANTENNA__3829__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout542 fanout542/A VGND VGND VPWR VPWR _5260_/C sky130_fd_sc_hd__buf_12
Xfanout564 fanout569/X VGND VGND VPWR VPWR _4128_/B sky130_fd_sc_hd__clkbuf_16
Xfanout575 fanout587/X VGND VGND VPWR VPWR fanout575/X sky130_fd_sc_hd__buf_12
Xfanout586 fanout587/X VGND VGND VPWR VPWR fanout586/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__6228__B1 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout597 fanout606/X VGND VGND VPWR VPWR fanout597/X sky130_fd_sc_hd__buf_12
XANTENNA_input124_A wb_adr_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__A1 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5659__A _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6093__B_N _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6400__B1 _6398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6703__A1 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3517__A1 _7242_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4190__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7579__RESET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6219__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7161__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5442__A1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4473__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4930_ _4930_/A _4930_/B _4930_/C VGND VGND VPWR VPWR _4934_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_47_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4861_ _4861_/A _4861_/B _4974_/C _4974_/D VGND VGND VPWR VPWR _4861_/X sky130_fd_sc_hd__and4_4
XFILLER_0_129_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6600_ _7501_/Q _6600_/B _6651_/C VGND VGND VPWR VPWR _6600_/X sky130_fd_sc_hd__and3_1
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3812_ _7489_/Q _3569_/X _3669_/X _6969_/Q _3811_/X VGND VGND VPWR VPWR _3812_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_16 _6594_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7580_ _7580_/CLK _7580_/D fanout596/X VGND VGND VPWR VPWR _7580_/Q sky130_fd_sc_hd__dfrtp_2
X_4792_ _4700_/Y _4789_/Y _4791_/Y VGND VGND VPWR VPWR _4800_/C sky130_fd_sc_hd__o21ai_1
XANTENNA_27 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3756__A1 _7554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ _7434_/Q _6747_/B _6747_/C _6447_/X _7442_/Q VGND VGND VPWR VPWR _6531_/X
+ sky130_fd_sc_hd__a32o_1
X_3743_ _7562_/Q hold72/A _4231_/S input38/X _3742_/X VGND VGND VPWR VPWR _3743_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3756__B2 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4412__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6462_ _6435_/B _6463_/A _6651_/B _6462_/D VGND VGND VPWR VPWR _6462_/X sky130_fd_sc_hd__and4b_4
X_3674_ _4449_/B _5612_/C hold56/A VGND VGND VPWR VPWR _5581_/A sky130_fd_sc_hd__and3_4
XFILLER_0_113_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5413_ _5538_/B _5569_/A _5568_/A _5488_/B VGND VGND VPWR VPWR _5416_/B sky130_fd_sc_hd__and4_1
X_6393_ _7213_/Q _6110_/A _6089_/X _6092_/X _7181_/Q VGND VGND VPWR VPWR _6393_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6170__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5344_ _4743_/A _5073_/A _4846_/Y _5204_/X VGND VGND VPWR VPWR _5506_/C sky130_fd_sc_hd__o31a_1
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6458__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput178 _3433_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 _3423_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_5275_ _5563_/A1 _4806_/Y _5255_/X _5274_/X VGND VGND VPWR VPWR _5278_/C sky130_fd_sc_hd__o31a_1
Xhold2903 hold2903/A VGND VGND VPWR VPWR _4462_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3552__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2914 hold2914/A VGND VGND VPWR VPWR hold2914/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2925 hold2925/A VGND VGND VPWR VPWR hold2925/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2936 hold2936/A VGND VGND VPWR VPWR _5583_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7014_ _7070_/CLK _7014_/D fanout590/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfrtp_4
X_4226_ _4226_/A0 _4225_/X _4232_/S VGND VGND VPWR VPWR _4226_/X sky130_fd_sc_hd__mux2_1
Xhold2947 _7496_/Q VGND VGND VPWR VPWR hold2947/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2958 hold2958/A VGND VGND VPWR VPWR _5921_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5681__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2969 _4226_/X VGND VGND VPWR VPWR hold990/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4157_ _7257_/Q _7306_/Q _4168_/D _7290_/Q VGND VGND VPWR VPWR _4157_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_0_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6225__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4088_ _4825_/A _5071_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _4088_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_0_167_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_179_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4814__C _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3747__A1 _7185_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_163_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6729_ _7014_/Q _4105_/B _6459_/B _6422_/X _6965_/Q VGND VGND VPWR VPWR _6729_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7278_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6161__A2 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1823_A _7538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold586_A _7336_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6449__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7409_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout361 _4725_/X VGND VGND VPWR VPWR _5453_/A sky130_fd_sc_hd__buf_6
XANTENNA__4277__B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7601__RESET_B fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout372 _5659_/B VGND VGND VPWR VPWR _5640_/C sky130_fd_sc_hd__buf_12
Xfanout383 _3492_/X VGND VGND VPWR VPWR _5947_/A sky130_fd_sc_hd__buf_12
Xfanout394 _4933_/A VGND VGND VPWR VPWR _4929_/A sky130_fd_sc_hd__buf_12
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6216__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5424__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_62_csclk_A _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__B2 _7463_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3637__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _4175_/A sky130_fd_sc_hd__buf_8
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_4
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _4076_/B sky130_fd_sc_hd__buf_12
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_2
Xhold809 hold809/A VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_122_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap539 _4717_/B VGND VGND VPWR VPWR _4765_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6152__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5060_ _5060_/A _5060_/B _5060_/C VGND VGND VPWR VPWR _5064_/A sky130_fd_sc_hd__nor3_1
Xhold1509 _7526_/Q VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5998__S hold37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5663__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4011_ _6910_/Q _6909_/Q _6908_/Q _7073_/Q VGND VGND VPWR VPWR _4011_/X sky130_fd_sc_hd__and4_2
XANTENNA__4915__B _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5415__B2 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5962_ _5962_/A0 _5998_/A1 _5964_/S VGND VGND VPWR VPWR _5962_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_176_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4913_ _4913_/A _4913_/B _4913_/C VGND VGND VPWR VPWR _4916_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5893_ _5893_/A _5902_/B VGND VGND VPWR VPWR _5893_/Y sky130_fd_sc_hd__nand2_8
X_7632_ _7636_/CLK _7632_/D VGND VGND VPWR VPWR _7632_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4931__A _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4844_ _4887_/B _4879_/C _5091_/A VGND VGND VPWR VPWR _4844_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__6376__C1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7563_ _7563_/CLK _7563_/D fanout602/X VGND VGND VPWR VPWR _7563_/Q sky130_fd_sc_hd__dfrtp_4
X_4775_ _5387_/C _4790_/B _4775_/C VGND VGND VPWR VPWR _4776_/A sky130_fd_sc_hd__and3_1
XFILLER_0_133_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6514_ _7441_/Q _6424_/C _6771_/A3 _6513_/X VGND VGND VPWR VPWR _6514_/X sky130_fd_sc_hd__a31o_1
X_3726_ _7307_/Q _5686_/A _3667_/X _7025_/Q _3725_/X VGND VGND VPWR VPWR _3726_/X
+ sky130_fd_sc_hd__a221o_1
X_7494_ _7580_/CLK _7494_/D fanout594/X VGND VGND VPWR VPWR _7494_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6679__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6445_ _7535_/Q _6408_/D _6420_/A _7295_/Q _6444_/X VGND VGND VPWR VPWR _6445_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3657_ _5640_/B _5612_/C _5659_/B VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__and3_4
XFILLER_0_30_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4154__A1 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5351__B1 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6376_ _6960_/Q _6036_/Y _6362_/Y _6375_/X _6775_/B1 VGND VGND VPWR VPWR _6376_/Y
+ sky130_fd_sc_hd__o221ai_4
X_3588_ _7541_/Q _3590_/C _5947_/B _3544_/X _7421_/Q VGND VGND VPWR VPWR _3588_/X
+ sky130_fd_sc_hd__a32o_1
X_5327_ _4743_/A _5072_/B _5295_/C _5260_/D VGND VGND VPWR VPWR _5339_/B sky130_fd_sc_hd__a211o_4
XANTENNA_fanout491_A _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2700 hold708/X VGND VGND VPWR VPWR _4393_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout589_A fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2711 hold833/X VGND VGND VPWR VPWR _4514_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2722 _4556_/X VGND VGND VPWR VPWR hold824/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5258_ _5260_/C _5387_/D _4755_/C _5257_/X VGND VGND VPWR VPWR _5266_/A sky130_fd_sc_hd__a31o_1
Xhold2733 _4270_/X VGND VGND VPWR VPWR hold849/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2744 hold2744/A VGND VGND VPWR VPWR _5750_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2755 _4245_/X VGND VGND VPWR VPWR hold2755/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4209_ _4209_/A0 _5863_/A0 _4211_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
Xhold2766 hold856/X VGND VGND VPWR VPWR _4381_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2777 _7141_/Q VGND VGND VPWR VPWR hold860/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5189_ _4929_/A _5180_/B _5034_/C _5031_/B VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__a31o_1
Xhold2788 hold2788/A VGND VGND VPWR VPWR hold2788/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2799 hold2799/A VGND VGND VPWR VPWR _4450_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5406__A1 _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6603__B1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3968__A1 _7279_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1773_A _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6382__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6134__A2 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4145__A1 _7562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input52_A mgmt_gpio_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4227__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3959__A1 _7503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5176__A3 _4971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6373__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4560_ _4825_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _5089_/C sky130_fd_sc_hd__nor3_4
XFILLER_0_182_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2087_A _7242_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3511_ _3511_/A _3557_/B _3511_/C VGND VGND VPWR VPWR _3511_/X sky130_fd_sc_hd__and3_2
Xhold606 hold606/A VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4491_ _4491_/A _4491_/B _4491_/C _4551_/D VGND VGND VPWR VPWR _4496_/S sky130_fd_sc_hd__and4_4
XFILLER_0_100_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold617 _4372_/X VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold628 hold628/A VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3442_ _7298_/Q VGND VGND VPWR VPWR _3442_/Y sky130_fd_sc_hd__inv_2
X_6230_ _7476_/Q _6032_/Y _6081_/X _7452_/Q _6229_/X VGND VGND VPWR VPWR _6230_/X
+ sky130_fd_sc_hd__a221o_1
Xhold639 hold639/A VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _7361_/Q _6332_/C _6158_/X _6160_/X VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a211o_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _7237_/Q VGND VGND VPWR VPWR hold574/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_110_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2018 _7044_/Q VGND VGND VPWR VPWR hold438/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2519_A _7143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _4828_/Y _5528_/A3 _5200_/C _4747_/B _5111_/Y VGND VGND VPWR VPWR _5112_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 hold609/X VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6092_ _6112_/C _6119_/A _6119_/B _6121_/A VGND VGND VPWR VPWR _6092_/X sky130_fd_sc_hd__and4_4
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 hold3132/X VGND VGND VPWR VPWR _5631_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 hold3071/X VGND VGND VPWR VPWR hold3072/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _4984_/B _4984_/A _4672_/X _4660_/Y _4759_/Y VGND VGND VPWR VPWR _5044_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 _4347_/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1339 _4320_/A1 VGND VGND VPWR VPWR hold2768/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4926__A _4932_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_wbbd_sck _7645_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__4364__C _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6994_ _6999_/CLK _6994_/D VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5945_ _5945_/A0 hold61/X hold23/X VGND VGND VPWR VPWR _5945_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5876_ _5876_/A0 _5993_/A1 _5883_/S VGND VGND VPWR VPWR _5876_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7615_ _7621_/CLK _7615_/D fanout576/X VGND VGND VPWR VPWR _7615_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4827_ _5115_/A _5115_/B _5399_/C VGND VGND VPWR VPWR _4827_/X sky130_fd_sc_hd__and3_1
XFILLER_0_8_776 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6364__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4811__D _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7546_ _7580_/CLK _7546_/D fanout594/X VGND VGND VPWR VPWR _7546_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout504_A hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4758_ _5158_/A _4758_/B _5328_/B VGND VGND VPWR VPWR _4758_/X sky130_fd_sc_hd__and3_4
XFILLER_0_16_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3709_ _7151_/Q _3652_/X _3654_/X _7121_/Q _3655_/X VGND VGND VPWR VPWR _3709_/X
+ sky130_fd_sc_hd__a221o_1
X_7477_ _7478_/CLK _7477_/D fanout585/X VGND VGND VPWR VPWR _7477_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4689_ _4679_/C _4679_/A _5328_/B VGND VGND VPWR VPWR _4997_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_120_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4127__A1 _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6428_ _7594_/Q _6435_/B _6462_/D _7593_/Q VGND VGND VPWR VPWR _6459_/C sky130_fd_sc_hd__and4bb_4
XANTENNA__6667__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6100__B _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6359_ _7155_/Q _6072_/X _6099_/X _7029_/Q _6358_/X VGND VGND VPWR VPWR _6362_/B
+ sky130_fd_sc_hd__a221oi_4
Xhold3220 _7607_/Q VGND VGND VPWR VPWR _6260_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3231 _4115_/Y VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1619_A _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3242 _7608_/Q VGND VGND VPWR VPWR _6261_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3253 _7583_/Q VGND VGND VPWR VPWR _6002_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3264 _6897_/Q VGND VGND VPWR VPWR _4050_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold284_A _4078_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2530 _7230_/Q VGND VGND VPWR VPWR hold674/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3275 _7074_/Q VGND VGND VPWR VPWR _4005_/C sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5627__A1 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2541 _7405_/Q VGND VGND VPWR VPWR hold795/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2552 hold827/X VGND VGND VPWR VPWR _5999_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2563 _5642_/X VGND VGND VPWR VPWR hold703/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2574 hold839/X VGND VGND VPWR VPWR _5666_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3638__B1 _7452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1840 _7521_/Q VGND VGND VPWR VPWR hold362/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2585 hold967/X VGND VGND VPWR VPWR _4207_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2596 hold769/X VGND VGND VPWR VPWR _5814_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1851 hold507/X VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1862 _5663_/X VGND VGND VPWR VPWR hold347/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1873 _5846_/X VGND VGND VPWR VPWR hold123/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1884 hold310/X VGND VGND VPWR VPWR _5851_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1895 hold328/X VGND VGND VPWR VPWR _5771_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5089__D _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4571__A _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3810__B1 _3800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4290__B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6355__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4366__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6107__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6658__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output256_A _7233_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3877__B1 _3543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5618__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4168__D _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3892__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3629__B1 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3650__A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_178_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_187_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6594__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3991_ _7375_/Q _5785_/A _5911_/A _3658_/X _7112_/Q VGND VGND VPWR VPWR _3991_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5730_ _5730_/A0 _5991_/A1 _5730_/S VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3801__B1 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5661_ _5661_/A0 _5967_/A1 _5667_/S VGND VGND VPWR VPWR _5661_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6346__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5149__A3 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2371_A _7198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7400_ _7476_/CLK _7400_/D fanout578/X VGND VGND VPWR VPWR _7400_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__4357__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4612_ _4571_/Y _5387_/B _4814_/C VGND VGND VPWR VPWR _4909_/C sky130_fd_sc_hd__o21ai_4
XANTENNA_hold2469_A _7288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5592_ _5592_/A0 _5805_/A1 _5595_/S VGND VGND VPWR VPWR _5592_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7331_ _7363_/CLK _7331_/D fanout575/X VGND VGND VPWR VPWR _7331_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4543_ _4543_/A0 _5647_/A0 hold57/X VGND VGND VPWR VPWR _4543_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold403 hold403/A VGND VGND VPWR VPWR _7401_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold414 hold414/A VGND VGND VPWR VPWR hold414/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4109__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4420__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold425 hold425/A VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3580__A2 _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold436 hold436/A VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7262_ _7578_/CLK _7262_/D fanout604/X VGND VGND VPWR VPWR _7262_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4474_ _4474_/A0 _5840_/A1 _4478_/S VGND VGND VPWR VPWR _4474_/X sky130_fd_sc_hd__mux2_1
Xhold447 hold447/A VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold458 hold458/A VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3544__B _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6213_ _7283_/Q _6036_/Y _6775_/B1 VGND VGND VPWR VPWR _6213_/Y sky130_fd_sc_hd__o21ai_1
Xhold469 hold469/A VGND VGND VPWR VPWR _7262_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3425_ _7442_/Q VGND VGND VPWR VPWR _3425_/Y sky130_fd_sc_hd__inv_2
X_7193_ _7213_/CLK _7193_/D fanout590/X VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3868__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2803_A _7137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6144_/A _6144_/B _6144_/C VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__and3_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5609__A1 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 hold2859/X VGND VGND VPWR VPWR _7415_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3883__A3 _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1114 _5583_/X VGND VGND VPWR VPWR _7210_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6112_/C _6136_/B _6136_/C VGND VGND VPWR VPWR _6075_/X sky130_fd_sc_hd__and3_4
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_7__f_wb_clk_i clkbuf_3_3_0_wb_clk_i/X VGND VGND VPWR VPWR _7627_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1125 hold2715/X VGND VGND VPWR VPWR hold2716/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5085__A2 _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6574__C _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1136 _4336_/X VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1147 hold2984/X VGND VGND VPWR VPWR hold2985/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1158 hold1158/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
X_5026_ _5026_/A _5026_/B _5026_/C VGND VGND VPWR VPWR _5028_/A sky130_fd_sc_hd__nor3_1
XANTENNA__4293__A0 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1169 hold2782/X VGND VGND VPWR VPWR hold2783/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3635__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6871__A _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6034__A1 _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7636_/CLK _6977_/D VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6585__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6894__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5928_ _5991_/A1 _5928_/A1 _5928_/S VGND VGND VPWR VPWR _5928_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3938__A4 _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4822__C _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6337__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5859_ hold43/X _5859_/A1 _5865_/S VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4348__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7445__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7529_ _7563_/CLK _7529_/D fanout599/X VGND VGND VPWR VPWR _7529_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_160_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold970 _5615_/X VGND VGND VPWR VPWR _7244_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold981 hold981/A VGND VGND VPWR VPWR hold981/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold992 _4476_/X VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input154_A wb_dat_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4520__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3050 _7229_/Q VGND VGND VPWR VPWR hold3050/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3061 _4235_/X VGND VGND VPWR VPWR hold3061/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3874__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3072 hold3072/A VGND VGND VPWR VPWR _5620_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3083 hold3083/A VGND VGND VPWR VPWR _5939_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3094 hold3094/A VGND VGND VPWR VPWR _5894_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2360 hold106/X VGND VGND VPWR VPWR _5727_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2371 _7198_/Q VGND VGND VPWR VPWR hold624/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2382 hold995/X VGND VGND VPWR VPWR _5773_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2393 _7174_/Q VGND VGND VPWR VPWR hold911/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input15_A mask_rev_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1670 _4209_/X VGND VGND VPWR VPWR hold283/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3626__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1681 hold251/X VGND VGND VPWR VPWR _5836_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1692 _7340_/Q VGND VGND VPWR VPWR hold358/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6781__A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6025__A1 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6576__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5784__A0 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4339__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4240__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6500__A2 _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4511__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4190_ _4190_/A0 _5979_/A0 _4190_/S VGND VGND VPWR VPWR _4190_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6264__A1 _7294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4907__C _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6264__B2 _7302_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6900_ _7075_/CLK _6900_/D _6850_/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6831_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6831_/X sky130_fd_sc_hd__and2_1
XFILLER_0_159_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6567__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4415__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6762_ _7186_/Q _6574_/B _6771_/A3 _6468_/X _7146_/Q VGND VGND VPWR VPWR _6762_/X
+ sky130_fd_sc_hd__a32o_1
X_3974_ _6957_/Q _3657_/X _4485_/A _7142_/Q VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_174_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5100__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5713_ _5713_/A hold47/X VGND VGND VPWR VPWR _5721_/S sky130_fd_sc_hd__nand2_8
X_6693_ _7067_/Q _6463_/A _6441_/X _6466_/X _7210_/Q VGND VGND VPWR VPWR _6693_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6319__A2 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5644_ _5948_/A1 _5644_/A1 _5649_/S VGND VGND VPWR VPWR _5644_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5575_ _5575_/A _5575_/B _5575_/C VGND VGND VPWR VPWR _5575_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_170_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5542__A3 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold200 hold200/A VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3555__A _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7314_ _7412_/CLK _7314_/D fanout580/X VGND VGND VPWR VPWR _7314_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4150__S _6898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold211 hold211/A VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4526_ _4526_/A0 _5586_/A0 _4526_/S VGND VGND VPWR VPWR _4526_/X sky130_fd_sc_hd__mux2_1
Xhold222 hold222/A VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold233 hold233/A VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold244 hold244/A VGND VGND VPWR VPWR _7330_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold255 hold255/A VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7245_ _7366_/CLK _7245_/D fanout582/X VGND VGND VPWR VPWR _7245_/Q sky130_fd_sc_hd__dfrtp_4
X_4457_ _4457_/A0 _5583_/A0 _4460_/S VGND VGND VPWR VPWR _4457_/X sky130_fd_sc_hd__mux2_1
Xhold266 hold266/A VGND VGND VPWR VPWR _7313_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold277 hold277/A VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold288 hold288/A VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold299 hold299/A VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3408_ _6751_/S VGND VGND VPWR VPWR _6067_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7176_ _7176_/CLK _7176_/D fanout590/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_4
X_4388_ hold56/X _4388_/B _5596_/B _5640_/D VGND VGND VPWR VPWR _4393_/S sky130_fd_sc_hd__nand4_4
XANTENNA_input7_A mask_rev_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _7496_/Q _6094_/A _6084_/X _6120_/X _7336_/Q VGND VGND VPWR VPWR _6127_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout571_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6462_/D _6435_/B _6747_/B VGND VGND VPWR VPWR _6058_/X sky130_fd_sc_hd__and3_4
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4596__A_N _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _5024_/A1 _4669_/X _4996_/A _4974_/B VGND VGND VPWR VPWR _5013_/C sky130_fd_sc_hd__o211a_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6558__A2 _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1686_A _7234_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5766__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6106__A _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5230__A2 _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7072__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7626__RESET_B fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4271__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6191__B1 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6730__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6479__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3847__A3 _3519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4296__A _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6246__A1 _7517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2190 _7374_/Q VGND VGND VPWR VPWR hold496/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_59_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5839__B _5911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4743__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6549__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4235__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3783__A2 _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3690_ _7331_/Q _3933_/A _3669_/C _3666_/X _7015_/Q VGND VGND VPWR VPWR _3690_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6182__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6721__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2167_A _6925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput305 _4166_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
X_5360_ _5213_/A _4929_/A _5346_/X _5231_/C VGND VGND VPWR VPWR _5444_/A sky130_fd_sc_hd__a31oi_2
XFILLER_0_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput316 hold1187/X VGND VGND VPWR VPWR hold1188/A sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_57_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput327 hold2810/X VGND VGND VPWR VPWR hold1152/A sky130_fd_sc_hd__buf_6
X_4311_ _4321_/S _3996_/B _4310_/Y VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__o21ai_1
Xoutput338 hold1195/X VGND VGND VPWR VPWR hold1196/A sky130_fd_sc_hd__buf_6
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5291_ _4821_/Y _4858_/Y _4672_/X _4873_/X _4679_/Y VGND VGND VPWR VPWR _5506_/B
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5590__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6485__A1 _7480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7030_ _7196_/CLK _7030_/D fanout590/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfrtp_4
X_4242_ _5655_/A1 hold84/X _4248_/S VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4918__B _4932_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3838__A3 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4173_ _4173_/A _4173_/B VGND VGND VPWR VPWR _4173_/X sky130_fd_sc_hd__and2_1
XANTENNA__6625__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5460__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5749__B hold12/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6814_ _7111_/Q _6814_/A2 _6814_/B1 _7109_/Q VGND VGND VPWR VPWR _6814_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6745_ _7212_/Q _6466_/X _6467_/X _7155_/Q _6744_/X VGND VGND VPWR VPWR _6745_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3957_ _7479_/Q _3535_/X _3673_/X _7197_/Q _3956_/X VGND VGND VPWR VPWR _3957_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4971__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3774__A2 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout417_A hold21/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6676_ _6675_/X _6676_/A1 _6777_/S VGND VGND VPWR VPWR _7623_/D sky130_fd_sc_hd__mux2_1
X_3888_ _7512_/Q _5920_/A _3881_/X _3884_/X _3887_/X VGND VGND VPWR VPWR _3888_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_5627_ _5627_/A0 _5863_/A0 _5629_/S VGND VGND VPWR VPWR _5627_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6173__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6712__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5558_ _5061_/B _4827_/X _5115_/X _4645_/D _5324_/A VGND VGND VPWR VPWR _5559_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4509_ _4509_/A _5612_/C _5596_/B _5902_/B VGND VGND VPWR VPWR _4514_/S sky130_fd_sc_hd__and4_4
X_5489_ _5038_/A _5127_/A _5118_/C _5164_/A VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__a31o_1
X_7228_ _7231_/CLK _7228_/D _4128_/B VGND VGND VPWR VPWR _7228_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6476__B2 _7440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4487__A0 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout510 _6116_/B VGND VGND VPWR VPWR _6121_/C sky130_fd_sc_hd__buf_12
XANTENNA_hold197_A _7289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout521 _7591_/Q VGND VGND VPWR VPWR _6112_/D sky130_fd_sc_hd__clkbuf_8
Xfanout532 _4937_/C VGND VGND VPWR VPWR _5180_/B sky130_fd_sc_hd__buf_12
Xfanout543 _4704_/Y VGND VGND VPWR VPWR _5387_/C sky130_fd_sc_hd__buf_12
X_7159_ _7268_/CLK _7159_/D _6871_/A VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfstp_2
Xfanout565 fanout569/X VGND VGND VPWR VPWR fanout565/X sky130_fd_sc_hd__buf_12
Xfanout576 fanout587/X VGND VGND VPWR VPWR fanout576/X sky130_fd_sc_hd__clkbuf_16
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout587 fanout606/X VGND VGND VPWR VPWR fanout587/X sky130_fd_sc_hd__buf_12
Xfanout598 fanout602/X VGND VGND VPWR VPWR fanout598/X sky130_fd_sc_hd__buf_12
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5659__B _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A wb_adr_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6400__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3765__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input82_A spi_sdoenb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6164__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6703__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3517__A2 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6219__A1 _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5978__A0 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5442__A2 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7548__RESET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4473__B _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4860_ _4860_/A _4860_/B VGND VGND VPWR VPWR _4933_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_87_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ _7289_/Q _4212_/A _4346_/C _3666_/X _7013_/Q VGND VGND VPWR VPWR _3811_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4791_ _4791_/A _4791_/B VGND VGND VPWR VPWR _4791_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_17 _6631_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _7554_/Q _6408_/A _6463_/X _7426_/Q VGND VGND VPWR VPWR _6530_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3742_ _7140_/Q _5965_/A _4521_/B _3531_/X _7338_/Q VGND VGND VPWR VPWR _3742_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3756__A2 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4920__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6155__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6461_ _7383_/Q _6460_/X _6459_/X _6458_/X _6456_/X VGND VGND VPWR VPWR _6471_/B
+ sky130_fd_sc_hd__a2111o_2
XFILLER_0_179_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3673_ _4551_/A _5866_/B _4551_/C VGND VGND VPWR VPWR _3673_/X sky130_fd_sc_hd__and3_2
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5412_ _5406_/Y _4783_/Y _5150_/A _5311_/B VGND VGND VPWR VPWR _5488_/B sky130_fd_sc_hd__o211a_1
X_6392_ _7186_/Q _6097_/X _6110_/X _7176_/Q _6391_/X VGND VGND VPWR VPWR _6397_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5343_ _5343_/A _5343_/B _5343_/C VGND VGND VPWR VPWR _5343_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4929__A _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput179 _3432_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4469__A0 _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5274_ _5255_/X _4798_/Y _5476_/A _5272_/X VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__o211a_1
Xhold2904 _7544_/Q VGND VGND VPWR VPWR hold2904/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3552__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7013_ _7189_/CLK _7013_/D fanout572/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfstp_2
Xhold2915 _7629_/Q VGND VGND VPWR VPWR _6781_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2926 _7052_/Q VGND VGND VPWR VPWR hold2926/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4225_ _4255_/A0 _5997_/A1 _4231_/S VGND VGND VPWR VPWR _4225_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5130__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2937 _7020_/Q VGND VGND VPWR VPWR hold698/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5130__B2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2948 hold2948/A VGND VGND VPWR VPWR _5904_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2959 _5921_/X VGND VGND VPWR VPWR _7511_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4156_ _6941_/Q input3/X input1/X VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_4
X_4087_ _5071_/B _5071_/C VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6394__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4989_ _5138_/D _5038_/B _5038_/C VGND VGND VPWR VPWR _5039_/A sky130_fd_sc_hd__and3_1
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6728_ _7593_/Q _7120_/Q _6408_/C _6409_/X _7135_/Q VGND VGND VPWR VPWR _6728_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6146__B1 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6659_ _7011_/Q _6423_/X _6462_/X _7031_/Q _6658_/X VGND VGND VPWR VPWR _6659_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6449__A1 _7311_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5121__A1 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout373 _3557_/X VGND VGND VPWR VPWR _5659_/B sky130_fd_sc_hd__buf_12
Xfanout384 _3492_/X VGND VGND VPWR VPWR _3590_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6621__A1 _7469_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5188__A1 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6385__B1 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4740__C _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_2
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3637__B _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6137__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_2
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3653__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3910__A2 _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5112__B2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4010_ _6910_/Q _6909_/Q _6908_/Q VGND VGND VPWR VPWR _4010_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__6612__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5961_ _5961_/A0 _5997_/A1 _5964_/S VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__mux2_1
X_4912_ _4943_/B _4915_/C VGND VGND VPWR VPWR _4913_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3977__A2 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5892_ _5892_/A0 _5991_/A1 _5892_/S VGND VGND VPWR VPWR _5892_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7631_ _7636_/CLK _7631_/D VGND VGND VPWR VPWR _7631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4843_ _4843_/A _5073_/B VGND VGND VPWR VPWR _5453_/C sky130_fd_sc_hd__nor2_8
XFILLER_0_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4423__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3729__A2 _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7562_ _7566_/CLK _7562_/D fanout599/X VGND VGND VPWR VPWR _7562_/Q sky130_fd_sc_hd__dfrtp_4
X_4774_ _5387_/C _4775_/C VGND VGND VPWR VPWR _4774_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_28_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6391__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6513_ _7465_/Q _6434_/B _6771_/A3 _6466_/X _7505_/Q VGND VGND VPWR VPWR _6513_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6128__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3725_ _7259_/Q _5619_/B _5659_/B _4497_/A _7156_/Q VGND VGND VPWR VPWR _3725_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_15_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7493_ _7581_/CLK _7493_/D fanout585/X VGND VGND VPWR VPWR _7493_/Q sky130_fd_sc_hd__dfrtp_2
X_6444_ _7447_/Q _6467_/A _6771_/A3 _6423_/X _7327_/Q VGND VGND VPWR VPWR _6444_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3656_ _4473_/A _5830_/C _4551_/C VGND VGND VPWR VPWR _4370_/A sky130_fd_sc_hd__and3_4
XFILLER_0_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5351__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6375_ _6110_/A _6365_/X _6370_/X _6374_/X VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__a211o_2
X_3587_ _3587_/A _3587_/B _3587_/C _3587_/D VGND VGND VPWR VPWR _3607_/B sky130_fd_sc_hd__nor4_2
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3563__A _7302_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5326_ _4672_/X _4980_/X _5174_/Y _5325_/X VGND VGND VPWR VPWR _5423_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3901__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2701 _7136_/Q VGND VGND VPWR VPWR hold797/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2712 _4514_/X VGND VGND VPWR VPWR hold834/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5257_ _5255_/X _5077_/Y _4765_/B _4803_/A VGND VGND VPWR VPWR _5257_/X sky130_fd_sc_hd__a2bb2o_1
Xhold2723 _7055_/Q VGND VGND VPWR VPWR hold811/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout484_A _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2734 _7279_/Q VGND VGND VPWR VPWR hold2734/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2745 _7176_/Q VGND VGND VPWR VPWR hold815/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2756 _7295_/Q VGND VGND VPWR VPWR hold2756/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4208_ _4208_/A0 _5754_/A1 _4211_/S VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__mux2_1
Xhold2767 _6999_/Q VGND VGND VPWR VPWR _4320_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2778 hold860/X VGND VGND VPWR VPWR _4484_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5188_ _5295_/C _5183_/C _4861_/X VGND VGND VPWR VPWR _5188_/X sky130_fd_sc_hd__o21a_1
Xhold2789 _6974_/Q VGND VGND VPWR VPWR _4281_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_4139_ _7269_/Q input89/X _4142_/A VGND VGND VPWR VPWR _4139_/X sky130_fd_sc_hd__mux2_2
XANTENNA__4394__A _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6603__B2 _7533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3968__A2 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6367__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_190_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4569__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3473__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4719__D _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input45_A mgmt_gpio_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6784__A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3959__A2 _5911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4081__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6358__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4243__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4908__A1 wire533/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3510_ _7582_/Q _3501_/X _3503_/X input33/X _3509_/X VGND VGND VPWR VPWR _3524_/B
+ sky130_fd_sc_hd__a221o_1
Xwire560 _5089_/C VGND VGND VPWR VPWR _4823_/C sky130_fd_sc_hd__clkbuf_4
X_4490_ _5754_/A1 _4490_/A1 _4490_/S VGND VGND VPWR VPWR _4490_/X sky130_fd_sc_hd__mux2_1
Xhold607 hold607/A VGND VGND VPWR VPWR _7478_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold618 hold618/A VGND VGND VPWR VPWR hold618/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_122_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold629 hold629/A VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3441_ _7314_/Q VGND VGND VPWR VPWR _3441_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6530__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4479__A _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6160_ _7297_/Q _6074_/X _6079_/X _7329_/Q _6159_/X VGND VGND VPWR VPWR _6160_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5111_/A _5111_/B _5111_/C VGND VGND VPWR VPWR _5111_/Y sky130_fd_sc_hd__nor3_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 hold574/X VGND VGND VPWR VPWR _5606_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2019 hold438/X VGND VGND VPWR VPWR _4374_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6112_/D _6119_/B _6121_/A VGND VGND VPWR VPWR _6091_/X sky130_fd_sc_hd__and3_4
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5802__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1307 hold2944/X VGND VGND VPWR VPWR hold2945/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6__f_wb_clk_i clkbuf_3_3_0_wb_clk_i/X VGND VGND VPWR VPWR _7610_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__7563__RESET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1318 hold3073/X VGND VGND VPWR VPWR _7248_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5042_ _5042_/A _5042_/B VGND VGND VPWR VPWR _5044_/A sky130_fd_sc_hd__nor2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1329 hold3172/X VGND VGND VPWR VPWR hold3173/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_109_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4418__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6993_ _6999_/CLK _6993_/D VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_51_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7412_/CLK sky130_fd_sc_hd__clkbuf_16
X_5944_ _5944_/A0 _5998_/A1 hold23/X VGND VGND VPWR VPWR _5944_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_164_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6349__B1 _6090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5875_ _5875_/A _5947_/A _5902_/B VGND VGND VPWR VPWR _5883_/S sky130_fd_sc_hd__and3_4
XFILLER_0_118_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3558__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4153__S _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7614_ _7627_/CLK _7614_/D fanout566/X VGND VGND VPWR VPWR _7614_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4826_ _5115_/A _5115_/B VGND VGND VPWR VPWR _4826_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_csclk _7496_/CLK VGND VGND VPWR VPWR _7417_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_788 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7545_ _7580_/CLK _7545_/D fanout594/X VGND VGND VPWR VPWR _7545_/Q sky130_fd_sc_hd__dfrtp_4
X_4757_ _4692_/Y _4730_/Y _4741_/Y _4755_/Y VGND VGND VPWR VPWR _4760_/C sky130_fd_sc_hd__o22a_1
XFILLER_0_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3583__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3708_ input7/X _5983_/A _3485_/X _3532_/X input56/X VGND VGND VPWR VPWR _3708_/X
+ sky130_fd_sc_hd__a32o_1
X_7476_ _7476_/CLK _7476_/D fanout581/X VGND VGND VPWR VPWR _7476_/Q sky130_fd_sc_hd__dfrtp_2
X_4688_ _4088_/Y _4558_/X _4591_/Y VGND VGND VPWR VPWR _5328_/B sky130_fd_sc_hd__o21a_4
X_6427_ _6427_/A _6455_/B _6467_/A VGND VGND VPWR VPWR _6427_/X sky130_fd_sc_hd__and3_4
XANTENNA__6521__B1 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3639_ _7580_/Q _3501_/X _5643_/A _7673_/A _3638_/X VGND VGND VPWR VPWR _3642_/C
+ sky130_fd_sc_hd__a221o_4
X_6358_ _7200_/Q _6110_/A _6079_/X _6120_/X _7019_/Q VGND VGND VPWR VPWR _6358_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3886__A1 _7480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3210 _7107_/Q VGND VGND VPWR VPWR _4171_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3221 _7638_/Q VGND VGND VPWR VPWR _6804_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6100__C _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3232 _7207_/Q VGND VGND VPWR VPWR _5566_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3886__B2 _7198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4539__D _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5309_ _4698_/Y _4755_/Y _4777_/X _4692_/Y _5150_/C VGND VGND VPWR VPWR _5311_/B
+ sky130_fd_sc_hd__o221a_1
Xhold3243 _7640_/Q VGND VGND VPWR VPWR _6810_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3254 _6890_/Q VGND VGND VPWR VPWR _4098_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6289_ _7041_/Q _6089_/X _6285_/X _6286_/X _6288_/X VGND VGND VPWR VPWR _6289_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold2520 hold694/X VGND VGND VPWR VPWR _4487_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3265 _7585_/Q VGND VGND VPWR VPWR _6012_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3276 _7597_/Q VGND VGND VPWR VPWR _6055_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2531 hold674/X VGND VGND VPWR VPWR _5598_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2542 hold795/X VGND VGND VPWR VPWR _5801_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2553 _7309_/Q VGND VGND VPWR VPWR hold791/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2564 _7333_/Q VGND VGND VPWR VPWR hold821/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3638__B2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2575 _5666_/X VGND VGND VPWR VPWR hold840/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1830 _3669_/C VGND VGND VPWR VPWR _4352_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1841 hold362/X VGND VGND VPWR VPWR _5932_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2586 _7317_/Q VGND VGND VPWR VPWR hold864/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2597 _5814_/X VGND VGND VPWR VPWR hold770/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1852 _6964_/Q VGND VGND VPWR VPWR hold456/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1863 hold347/X VGND VGND VPWR VPWR _7282_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1874 _7456_/Q VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5013__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1885 _5851_/X VGND VGND VPWR VPWR hold311/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1896 _5771_/X VGND VGND VPWR VPWR hold329/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6588__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7156_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold1883_A _7449_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6052__A2 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4571__B _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_164_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6760__B1 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold3264_A _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3574__B1 hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6107__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4118__A2 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5315__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6512__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3877__A1 _7027_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3877__B2 _7288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6815__A1 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3650__B _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4238__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6291__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6579__B1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3990_ input11/X _3490_/X _5686_/A _7303_/Q _3989_/X VGND VGND VPWR VPWR _3990_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_159_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3801__A1 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5660_ _5660_/A0 _5903_/A0 _5667_/S VGND VGND VPWR VPWR _5660_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4611_ _4814_/C _4608_/Y _4772_/A VGND VGND VPWR VPWR _4657_/C sky130_fd_sc_hd__o21bai_4
XFILLER_0_154_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5591_ _5591_/A0 _5948_/A1 _5595_/S VGND VGND VPWR VPWR _5591_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2364_A _7199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7330_ _7366_/CLK _7330_/D fanout582/X VGND VGND VPWR VPWR _7330_/Q sky130_fd_sc_hd__dfrtp_4
X_4542_ _4542_/A0 _5815_/A1 hold57/X VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold404 hold404/A VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold415 hold415/A VGND VGND VPWR VPWR _7369_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7261_ _7522_/CLK _7261_/D fanout603/X VGND VGND VPWR VPWR _7261_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6503__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold426 hold426/A VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4473_ _4473_/A _5619_/B _4551_/D VGND VGND VPWR VPWR _4478_/S sky130_fd_sc_hd__and3_2
Xhold437 hold437/A VGND VGND VPWR VPWR _7278_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold448 hold448/A VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold459 hold459/A VGND VGND VPWR VPWR _7302_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6212_ _6212_/A _6212_/B _6212_/C VGND VGND VPWR VPWR _6212_/Y sky130_fd_sc_hd__nor3_4
X_3424_ _7450_/Q VGND VGND VPWR VPWR _3424_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3544__C _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7192_ _7212_/CLK _7192_/D fanout574/X VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6143_ _6116_/B _6138_/X _6140_/X _6142_/X VGND VGND VPWR VPWR _6143_/X sky130_fd_sc_hd__a211o_2
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6806__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 hold2880/X VGND VGND VPWR VPWR hold2881/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6074_ _7588_/Q _6136_/C _7589_/Q VGND VGND VPWR VPWR _6074_/X sky130_fd_sc_hd__and3b_4
XANTENNA__3883__A4 _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1115 hold3003/X VGND VGND VPWR VPWR hold3004/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _4390_/X VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1137 hold2970/X VGND VGND VPWR VPWR hold2971/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6282__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5025_ _5025_/A _5185_/B _5025_/C _5025_/D VGND VGND VPWR VPWR _5026_/C sky130_fd_sc_hd__nand4_2
XANTENNA_hold2998_A _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1148 hold2986/X VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1159 hold2796/X VGND VGND VPWR VPWR hold2797/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_A _6072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6976_ _7206_/CLK _6976_/D VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5388__A4 _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5927_ hold61/X _5927_/A1 _5928_/S VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5793__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5858_ _5993_/A1 _5858_/A1 _5865_/S VGND VGND VPWR VPWR _5858_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6337__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4809_ _4809_/A _4809_/B _4809_/C VGND VGND VPWR VPWR _4812_/A sky130_fd_sc_hd__nor3_1
XANTENNA__6742__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5789_ _5789_/A0 _5987_/A1 _5793_/S VGND VGND VPWR VPWR _5789_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7528_ _7560_/CLK _7528_/D fanout599/X VGND VGND VPWR VPWR _7528_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7459_ _7487_/CLK _7459_/D fanout593/X VGND VGND VPWR VPWR _7459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_160_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold960 _4195_/X VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold971 hold971/A VGND VGND VPWR VPWR hold971/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold982 _4373_/X VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold993 hold993/A VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3040 _6961_/Q VGND VGND VPWR VPWR hold759/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4847__A _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3051 hold3051/A VGND VGND VPWR VPWR _5597_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3062 _7265_/Q VGND VGND VPWR VPWR hold3062/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3073 _5620_/X VGND VGND VPWR VPWR hold3073/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input147_A wb_dat_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3084 _7567_/Q VGND VGND VPWR VPWR hold3084/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4566__B _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2350 _7283_/Q VGND VGND VPWR VPWR hold100/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3095 _7543_/Q VGND VGND VPWR VPWR hold3095/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2361 _5727_/X VGND VGND VPWR VPWR hold107/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2372 hold624/X VGND VGND VPWR VPWR _4553_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2383 _7308_/Q VGND VGND VPWR VPWR hold921/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4284__A1 _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2394 hold911/X VGND VGND VPWR VPWR _4524_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1660 hold59/X VGND VGND VPWR VPWR _4199_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1671 _7204_/Q VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1682 _5836_/X VGND VGND VPWR VPWR hold252/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1693 hold358/X VGND VGND VPWR VPWR _5728_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6025__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4582__A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5233__B1 _5102_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_171_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5536__A1 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3547__B1 _3543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6500__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3661__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6264__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4275__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6830_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6830_/X sky130_fd_sc_hd__and2_1
XFILLER_0_82_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_53_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4923__C _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6567__A3 _6429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6761_ _7191_/Q _6446_/X _6452_/X _7025_/Q _6760_/X VGND VGND VPWR VPWR _6761_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5775__A1 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3973_ _7535_/Q _5947_/A _5947_/B _3972_/X VGND VGND VPWR VPWR _3973_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_119_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4642__D _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5712_ _5955_/A1 _5712_/A1 _5712_/S VGND VGND VPWR VPWR _5712_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_174_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6692_ _7123_/Q _6420_/C _6419_/A _7158_/Q _6691_/X VGND VGND VPWR VPWR _6697_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5643_ _5643_/A _5992_/D VGND VGND VPWR VPWR _5649_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_72_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5574_ _5574_/A _5574_/B VGND VGND VPWR VPWR _5575_/C sky130_fd_sc_hd__and2_1
XFILLER_0_115_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7313_ _7577_/CLK _7313_/D fanout583/X VGND VGND VPWR VPWR _7313_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3555__B _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold201 hold201/A VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4525_ _4525_/A0 _5852_/A0 _4526_/S VGND VGND VPWR VPWR _4525_/X sky130_fd_sc_hd__mux2_1
Xhold212 hold212/A VGND VGND VPWR VPWR hold212/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold223 hold223/A VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold234 hold234/A VGND VGND VPWR VPWR _7572_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold245 hold245/A VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7244_ _7366_/CLK _7244_/D fanout579/X VGND VGND VPWR VPWR _7244_/Q sky130_fd_sc_hd__dfrtp_4
Xhold256 hold256/A VGND VGND VPWR VPWR _7556_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4456_ _4456_/A0 _5840_/A1 _4460_/S VGND VGND VPWR VPWR _4456_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold267 hold267/A VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold278 hold278/A VGND VGND VPWR VPWR _7578_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3407_ _6932_/Q VGND VGND VPWR VPWR _6065_/C sky130_fd_sc_hd__inv_2
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold289 hold289/A VGND VGND VPWR VPWR _7370_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4667__A _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7175_ _7176_/CLK _7175_/D fanout588/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_4
X_4387_ _5586_/A0 _4387_/A1 _4387_/S VGND VGND VPWR VPWR _4387_/X sky130_fd_sc_hd__mux2_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _7528_/Q _6092_/X _6112_/X _7480_/Q _6125_/X VGND VGND VPWR VPWR _6126_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3710__B1 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6255__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6057_ _7594_/Q _7593_/Q _6600_/B VGND VGND VPWR VPWR _6747_/B sky130_fd_sc_hd__and3_4
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout564_A fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4266__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5008_ _5113_/A _5180_/B _5260_/D _5107_/A VGND VGND VPWR VPWR _5008_/X sky130_fd_sc_hd__o31a_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6007__A2 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6558__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4833__C _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6959_ _7024_/CLK _6959_/D fanout567/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6106__B _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4577__A _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold790 _5864_/X VGND VGND VPWR VPWR _7461_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3481__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3701__B1 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6246__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2180 _7292_/Q VGND VGND VPWR VPWR hold889/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5900__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4257__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2191 hold496/X VGND VGND VPWR VPWR _5766_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_188_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1490 _3496_/Y VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5757__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _4127_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5509__A1 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3783__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6706__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3656__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6032__A _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6721__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput306 _4174_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput317 hold1185/X VGND VGND VPWR VPWR hold1186/A sky130_fd_sc_hd__buf_6
X_4310_ _4321_/S _4310_/B VGND VGND VPWR VPWR _4310_/Y sky130_fd_sc_hd__nand2_1
Xoutput328 hold1197/X VGND VGND VPWR VPWR hold1198/A sky130_fd_sc_hd__buf_6
XFILLER_0_140_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3940__B1 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput339 hold2807/X VGND VGND VPWR VPWR hold1164/A sky130_fd_sc_hd__buf_6
X_5290_ _5252_/Y _5461_/B _4854_/X VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5590__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_wire365_A _4145_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4241_ _4241_/A0 _4240_/X _4249_/S VGND VGND VPWR VPWR _4241_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6485__A2 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5693__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4496__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4918__C _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4172_ _4178_/A _7110_/Q VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__and2_1
XANTENNA__4248__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5810__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5996__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5749__C _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6813_ _6812_/X _6813_/A1 _6822_/S VGND VGND VPWR VPWR _7641_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5748__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5212__A3 _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6744_ _7200_/Q _6463_/A _6771_/A3 _6419_/C _7140_/Q VGND VGND VPWR VPWR _6744_/X
+ sky130_fd_sc_hd__a32o_1
X_3956_ input98/X _5785_/B _5659_/B _4370_/A _7041_/Q VGND VGND VPWR VPWR _3956_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4420__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6675_ _6649_/S _6675_/A2 _6673_/X _6674_/X VGND VGND VPWR VPWR _6675_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_190_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3774__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3887_ _7133_/Q _3670_/X _4497_/A _7153_/Q _3886_/X VGND VGND VPWR VPWR _3887_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4161__S _7260_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5626_ _5626_/A0 _5950_/A1 _5629_/S VGND VGND VPWR VPWR _5626_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6173__A1 _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7077__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5557_ _5543_/X _5548_/Y _5556_/Y VGND VGND VPWR VPWR _5557_/X sky130_fd_sc_hd__a21o_1
X_4508_ _4508_/A0 _5754_/A1 _4508_/S VGND VGND VPWR VPWR _4508_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5488_ _5488_/A _5488_/B _5488_/C VGND VGND VPWR VPWR _5488_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__6476__A2 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7227_ _7231_/CLK _7227_/D fanout565/X VGND VGND VPWR VPWR _7227_/Q sky130_fd_sc_hd__dfrtp_4
X_4439_ _4439_/A0 _5991_/A1 _4439_/S VGND VGND VPWR VPWR _4439_/X sky130_fd_sc_hd__mux2_1
Xfanout500 hold2039/X VGND VGND VPWR VPWR hold2040/A sky130_fd_sc_hd__buf_6
Xfanout511 _6116_/B VGND VGND VPWR VPWR _6144_/C sky130_fd_sc_hd__clkbuf_16
Xfanout522 _7590_/Q VGND VGND VPWR VPWR _6106_/B sky130_fd_sc_hd__buf_12
X_7158_ _7191_/CLK _7158_/D _6871_/A VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout566 fanout569/X VGND VGND VPWR VPWR fanout566/X sky130_fd_sc_hd__buf_12
Xfanout577 fanout587/X VGND VGND VPWR VPWR fanout577/X sky130_fd_sc_hd__buf_12
XANTENNA__6228__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6109_ _6112_/D _6119_/B _6144_/A _6144_/C VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__and4_1
Xfanout588 fanout589/X VGND VGND VPWR VPWR fanout588/X sky130_fd_sc_hd__buf_12
X_7089_ _7530_/CLK hold95/X fanout600/X VGND VGND VPWR VPWR _7668_/A sky130_fd_sc_hd__dfrtp_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout599 fanout602/X VGND VGND VPWR VPWR fanout599/X sky130_fd_sc_hd__buf_12
XANTENNA__5987__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4844__B _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__A3 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5659__C _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5739__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5956__A _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3765__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6164__A1 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6164__B2 _7441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6703__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input75_A porb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5675__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4478__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6219__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6726__S _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4246__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5442__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4473__C _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _7553_/Q _3508_/X _3800_/X _3802_/X _3809_/X VGND VGND VPWR VPWR _3855_/A
+ sky130_fd_sc_hd__a2111oi_2
XANTENNA__4770__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4790_ _5387_/C _4790_/B _4790_/C VGND VGND VPWR VPWR _4791_/A sky130_fd_sc_hd__and3_1
XFILLER_0_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4402__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 _6712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7517__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _7120_/Q _5830_/C _5992_/C _3502_/X _3740_/X VGND VGND VPWR VPWR _3741_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4920__D _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6460_ _7596_/Q _7595_/Q _6467_/A _6651_/B VGND VGND VPWR VPWR _6460_/X sky130_fd_sc_hd__and4_4
XFILLER_0_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3672_ _4473_/A _5938_/B _4388_/B VGND VGND VPWR VPWR _4497_/A sky130_fd_sc_hd__and3_4
XFILLER_0_113_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5411_ _5408_/Y _4769_/Y _5145_/A _5306_/B VGND VGND VPWR VPWR _5568_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_3_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6391_ _7070_/Q _6110_/A _6332_/C _6075_/X _7166_/Q VGND VGND VPWR VPWR _6391_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5805__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5342_ _5342_/A _5342_/B _5342_/C VGND VGND VPWR VPWR _5343_/A sky130_fd_sc_hd__and3_2
XANTENNA__4929__B _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6458__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5273_ _5563_/A1 _4709_/Y _4806_/Y _4946_/Y _4798_/Y VGND VGND VPWR VPWR _5476_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2905 hold2905/A VGND VGND VPWR VPWR _5958_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7012_ _7112_/CLK _7012_/D fanout589/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3552__C _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2916 hold2916/A VGND VGND VPWR VPWR hold2916/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4224_ _4224_/A0 _4223_/X _4232_/S VGND VGND VPWR VPWR _4224_/X sky130_fd_sc_hd__mux2_1
Xhold2927 hold2927/A VGND VGND VPWR VPWR _4384_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2938 hold698/X VGND VGND VPWR VPWR _4345_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2949 _7463_/Q VGND VGND VPWR VPWR hold2949/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4155_ _4154_/X _4135_/B _6896_/Q VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_2
XANTENNA__4945__A _4945_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3692__A2 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4086_ _4825_/A _5071_/A VGND VGND VPWR VPWR _4086_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_179_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5969__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4156__S input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6630__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_176_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5776__A _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4680__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5197__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4988_ _5339_/D _5183_/A _5295_/C _5339_/C VGND VGND VPWR VPWR _5041_/D sky130_fd_sc_hd__nand4_1
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6727_ _6726_/X _6751_/A1 _6777_/S VGND VGND VPWR VPWR _7625_/D sky130_fd_sc_hd__mux2_1
X_3939_ _7137_/Q _4491_/B _4521_/B _4467_/A _7127_/Q VGND VGND VPWR VPWR _3939_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6658_ _7026_/Q _6651_/B _6459_/C _6408_/B _7041_/Q VGND VGND VPWR VPWR _6658_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4157__B1 _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5609_ _5609_/A0 _5863_/A0 _5611_/S VGND VGND VPWR VPWR _5609_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6589_ _7500_/Q _6600_/B _6651_/C _6468_/X _7412_/Q VGND VGND VPWR VPWR _6589_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6449__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5657__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout374 _3548_/X VGND VGND VPWR VPWR _5619_/B sky130_fd_sc_hd__buf_12
Xfanout385 _5587_/C VGND VGND VPWR VPWR _5612_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__3683__A2 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4574__B _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6621__A2 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4632__A1 _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5686__A _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5188__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4396__A0 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4740__D _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__6137__A1 _7288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6137__B2 _7328_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_4
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_4
XANTENNA__6688__A2 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5896__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5360__A2 _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3653__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5648__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5__f_wb_clk_i clkbuf_3_2_0_wb_clk_i/X VGND VGND VPWR VPWR _7621_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5112__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4320__A0 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5960_ _5960_/A0 _5987_/A1 _5964_/S VGND VGND VPWR VPWR _5960_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_149_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4911_ _5213_/B _4929_/A _5180_/B _4940_/D VGND VGND VPWR VPWR _4913_/B sky130_fd_sc_hd__nand4_4
X_5891_ _5891_/A0 hold61/X _5892_/S VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__mux2_1
XANTENNA__3977__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5596__A _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7630_ _7630_/CLK _7630_/D VGND VGND VPWR VPWR _7630_/Q sky130_fd_sc_hd__dfxtp_1
X_4842_ _4887_/B _5091_/A VGND VGND VPWR VPWR _4960_/A sky130_fd_sc_hd__nand2b_4
XFILLER_0_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4387__A0 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4773_ _5100_/A _4797_/B _5260_/C VGND VGND VPWR VPWR _5086_/B sky130_fd_sc_hd__and3_2
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3729__A3 _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7561_ _7563_/CLK _7561_/D fanout598/X VGND VGND VPWR VPWR _7561_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3724_ _6923_/Q _3542_/X _5704_/A _7323_/Q VGND VGND VPWR VPWR _3724_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_7_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6512_ _7513_/Q _6435_/X _6446_/X _7521_/Q VGND VGND VPWR VPWR _6512_/X sky130_fd_sc_hd__a22o_1
X_7492_ _7580_/CLK _7492_/D fanout594/X VGND VGND VPWR VPWR _7492_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6679__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6443_ _6455_/B _6467_/A _6447_/C VGND VGND VPWR VPWR _6443_/X sky130_fd_sc_hd__and3_4
X_3655_ _7672_/A hold36/A _4491_/A _4491_/B VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__and4_1
XFILLER_0_113_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6374_ _6877_/Q _6112_/X _6371_/X _6373_/X _6372_/X VGND VGND VPWR VPWR _6374_/X
+ sky130_fd_sc_hd__a2111o_1
X_3586_ _7357_/Q _3506_/X _5758_/A _7373_/Q _3585_/X VGND VGND VPWR VPWR _3587_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4659__B _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3563__B hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5325_ _5295_/B _4977_/X _5046_/A _5007_/Y VGND VGND VPWR VPWR _5325_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5639__A0 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5256_ _4601_/Y _4744_/Y _4716_/Y _5451_/A1 VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__a211o_1
Xhold2702 hold797/X VGND VGND VPWR VPWR _4478_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2713 _7171_/Q VGND VGND VPWR VPWR hold829/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_139_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2724 hold811/X VGND VGND VPWR VPWR _4387_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2735 hold2735/A VGND VGND VPWR VPWR _5660_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4207_ _4207_/A0 _5647_/A0 _4211_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
Xhold2746 hold815/X VGND VGND VPWR VPWR _4526_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2757 hold2757/A VGND VGND VPWR VPWR _5678_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5187_ _5178_/X _5038_/C _5186_/X _5185_/Y VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6793__B1_N _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_A _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2768 hold2768/A VGND VGND VPWR VPWR hold2768/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2779 _7026_/Q VGND VGND VPWR VPWR hold2779/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4138_ _7270_/Q input91/X _4142_/A VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_2
XANTENNA__4394__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6603__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4069_ hold15/A hold59/A _4075_/S VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_78_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6367__B2 _7034_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5024__D1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_834 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3738__B _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5327__C1 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1926_A _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4550__A0 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3473__B _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4302__A0 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input38_A mgmt_gpio_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5802__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3959__A3 _3496_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6358__A1 _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_826 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3664__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold608 hold608/A VGND VGND VPWR VPWR hold608/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6040__A _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3440_ _7322_/Q VGND VGND VPWR VPWR _3440_/Y sky130_fd_sc_hd__inv_2
Xhold619 hold619/A VGND VGND VPWR VPWR _7552_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6530__A1 _7554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4479__B _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3895__A2 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5110_ _5282_/B _5453_/B _5113_/B VGND VGND VPWR VPWR _5110_/X sky130_fd_sc_hd__and3_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2009 _5606_/X VGND VGND VPWR VPWR hold575/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6090_ _6119_/A _6119_/B _6116_/C _6121_/C VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__and4_4
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__B1 _6988_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A _5041_/B _5041_/C _5041_/D VGND VGND VPWR VPWR _5042_/B sky130_fd_sc_hd__nand4_1
Xhold1308 hold2946/X VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1319 hold3166/X VGND VGND VPWR VPWR hold3167/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4926__C _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_192_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4645__D _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_6992_ _7024_/CLK _6992_/D fanout568/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5943_ _5943_/A0 _5979_/A0 hold23/X VGND VGND VPWR VPWR _5943_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4942__B _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6349__B2 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5874_ _5874_/A0 _5991_/A1 _5874_/S VGND VGND VPWR VPWR _5874_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_164_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_192_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3558__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7613_ _7627_/CLK _7613_/D fanout566/X VGND VGND VPWR VPWR _7613_/Q sky130_fd_sc_hd__dfrtp_1
X_4825_ _4825_/A _5071_/B _5071_/C _5089_/B VGND VGND VPWR VPWR _4825_/Y sky130_fd_sc_hd__nor4_2
XFILLER_0_8_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7544_ _7580_/CLK _7544_/D fanout594/X VGND VGND VPWR VPWR _7544_/Q sky130_fd_sc_hd__dfstp_2
X_4756_ _5038_/A _5134_/A _5260_/C VGND VGND VPWR VPWR _4756_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3707_ _7547_/Q _5965_/A _4212_/A _3508_/X _7555_/Q VGND VGND VPWR VPWR _3707_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4687_ _5138_/B _4687_/B _4687_/C VGND VGND VPWR VPWR _4687_/Y sky130_fd_sc_hd__nand3_4
X_7475_ _7563_/CLK _7475_/D fanout599/X VGND VGND VPWR VPWR _7475_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_160_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6426_ _6462_/D _6435_/B _6467_/A VGND VGND VPWR VPWR _6426_/X sky130_fd_sc_hd__and3_4
X_3638_ _7572_/Q _5983_/A _5992_/C _7452_/Q _5848_/A VGND VGND VPWR VPWR _3638_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_48_csclk_A _7496_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3200 _6215_/X VGND VGND VPWR VPWR _7606_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3569_ _3569_/A _5947_/B _4491_/C VGND VGND VPWR VPWR _3569_/X sky130_fd_sc_hd__and3_4
X_6357_ _7059_/Q _6085_/X _6119_/X _7135_/Q _6356_/X VGND VGND VPWR VPWR _6357_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout594_A fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3211 _7621_/Q VGND VGND VPWR VPWR _6649_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6100__D _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3222 _6880_/Q VGND VGND VPWR VPWR _4121_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3233 _7642_/Q VGND VGND VPWR VPWR _6816_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5308_ _5308_/A _5308_/B _5308_/C VGND VGND VPWR VPWR _5311_/A sky130_fd_sc_hd__nor3_1
Xhold3244 _7609_/Q VGND VGND VPWR VPWR _6284_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6288_ _7112_/Q _6317_/C _6074_/X _6967_/Q _6287_/X VGND VGND VPWR VPWR _6288_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5088__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2510 _5594_/X VGND VGND VPWR VPWR hold956/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3255 _4066_/Y VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3266 _6909_/Q VGND VGND VPWR VPWR _4004_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2521 _7360_/Q VGND VGND VPWR VPWR hold686/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3277 _7588_/Q VGND VGND VPWR VPWR _6020_/S sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2532 _5598_/X VGND VGND VPWR VPWR hold675/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2543 _6912_/Q VGND VGND VPWR VPWR hold660/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5239_ _5222_/A _5453_/A _5453_/B _4934_/B _5237_/Y VGND VGND VPWR VPWR _5239_/X
+ sky130_fd_sc_hd__a311o_1
Xhold2554 hold791/X VGND VGND VPWR VPWR _5693_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_166_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2565 hold821/X VGND VGND VPWR VPWR _5720_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1820 _7569_/Q VGND VGND VPWR VPWR hold304/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3638__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4835__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1831 _4337_/X VGND VGND VPWR VPWR hold471/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4835__B2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2576 _7557_/Q VGND VGND VPWR VPWR hold803/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2587 hold864/X VGND VGND VPWR VPWR _5702_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1842 _7458_/Q VGND VGND VPWR VPWR hold300/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2598 _7512_/Q VGND VGND VPWR VPWR hold2598/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1853 hold456/X VGND VGND VPWR VPWR _4268_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1864 _7522_/Q VGND VGND VPWR VPWR hold350/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1875 hold63/X VGND VGND VPWR VPWR _5859_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1886 _6990_/Q VGND VGND VPWR VPWR hold512/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1897 hold329/X VGND VGND VPWR VPWR _7378_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7202__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3810__A2 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5563__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3574__B2 _7565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6512__A1 _7513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6512__B2 _7521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5903__S _5910_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3877__A2 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3931__B _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6276__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__buf_12
XANTENNA__3650__C _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output311_A _7628_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6579__B2 _7532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3659__A _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6035__A _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3801__A2 _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6200__B1 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4610_ _5100_/A _4645_/D VGND VGND VPWR VPWR _4657_/D sky130_fd_sc_hd__nand2_2
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5590_ _5590_/A _5596_/B _5640_/C _5640_/D VGND VGND VPWR VPWR _5595_/S sky130_fd_sc_hd__and4_4
X_4541_ _4541_/A0 hold43/X hold57/X VGND VGND VPWR VPWR _4541_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2357_A _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold405 hold405/A VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold416 hold416/A VGND VGND VPWR VPWR hold416/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4472_ _5979_/A0 _4472_/A1 _4472_/S VGND VGND VPWR VPWR _4472_/X sky130_fd_sc_hd__mux2_1
X_7260_ _7578_/CLK _7260_/D fanout604/X VGND VGND VPWR VPWR _7260_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold427 _5896_/X VGND VGND VPWR VPWR _7489_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6503__B2 _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold438 hold438/A VGND VGND VPWR VPWR hold438/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3423_ _7458_/Q VGND VGND VPWR VPWR _3423_/Y sky130_fd_sc_hd__inv_2
Xhold449 hold449/A VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6211_ _6094_/A _6202_/X _6207_/X _6210_/X VGND VGND VPWR VPWR _6212_/C sky130_fd_sc_hd__a211o_1
X_7191_ _7191_/CLK _7191_/D fanout573/X VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5813__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3868__A2 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _7456_/Q _6080_/X _6090_/X _7376_/Q _6141_/X VGND VGND VPWR VPWR _6142_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6267__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6119_/A _6106_/B _6144_/A VGND VGND VPWR VPWR _6073_/X sky130_fd_sc_hd__and3_4
Xhold1105 _5903_/X VGND VGND VPWR VPWR _7495_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 hold3005/X VGND VGND VPWR VPWR _7440_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5024_/A1 _4669_/X _4974_/B _5180_/A _5038_/A VGND VGND VPWR VPWR _5185_/B
+ sky130_fd_sc_hd__o2111ai_4
Xhold1127 hold2978/X VGND VGND VPWR VPWR hold2979/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1138 hold2972/X VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1149 hold3035/X VGND VGND VPWR VPWR hold3036/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5490__A1 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6078__A_N _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6416__B_N _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6975_ _7630_/CLK _6975_/D VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5242__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3569__A _3569_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4164__S _7259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5926_ _5998_/A1 _5926_/A1 _5928_/S VGND VGND VPWR VPWR _5926_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5857_ _5857_/A hold47/X VGND VGND VPWR VPWR _5865_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_63_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4808_ _5410_/A _5061_/B _5453_/B VGND VGND VPWR VPWR _4809_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout607_A _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5788_ _5788_/A0 _5914_/A1 _5793_/S VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7527_ _7560_/CLK _7527_/D fanout599/X VGND VGND VPWR VPWR _7527_/Q sky130_fd_sc_hd__dfstp_4
X_4739_ _4730_/Y _4732_/Y _4738_/X VGND VGND VPWR VPWR _5139_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7458_ _7566_/CLK _7458_/D fanout593/X VGND VGND VPWR VPWR _7458_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6111__C _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6409_ _6462_/D _6435_/B _6434_/B _6651_/B VGND VGND VPWR VPWR _6409_/X sky130_fd_sc_hd__and4_4
XFILLER_0_101_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold950 _5647_/X VGND VGND VPWR VPWR _7268_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7389_ _7577_/CLK _7389_/D fanout584/X VGND VGND VPWR VPWR _7389_/Q sky130_fd_sc_hd__dfrtp_4
Xhold961 hold961/A VGND VGND VPWR VPWR hold961/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5723__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold972 hold972/A VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold983 hold983/A VGND VGND VPWR VPWR hold983/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold994 _4482_/X VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3030 _5591_/X VGND VGND VPWR VPWR hold3030/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3041 hold759/X VGND VGND VPWR VPWR _4264_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_177_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3052 _5597_/X VGND VGND VPWR VPWR hold3052/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3063 hold3063/A VGND VGND VPWR VPWR _5644_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3074 _7455_/Q VGND VGND VPWR VPWR hold3074/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2340 _5661_/X VGND VGND VPWR VPWR hold593/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3085 hold3085/A VGND VGND VPWR VPWR _5984_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2351 hold100/X VGND VGND VPWR VPWR _5664_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3096 hold3096/A VGND VGND VPWR VPWR _5957_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2362 _7170_/Q VGND VGND VPWR VPWR hold917/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2373 _4553_/X VGND VGND VPWR VPWR hold625/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2384 hold921/X VGND VGND VPWR VPWR _5692_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1650 _7068_/Q VGND VGND VPWR VPWR hold374/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4284__A2 _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2395 _4524_/X VGND VGND VPWR VPWR hold912/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1993_A _7155_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1661 _4199_/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1672 hold33/X VGND VGND VPWR VPWR _3463_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1683 _7460_/Q VGND VGND VPWR VPWR hold338/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1694 _5728_/X VGND VGND VPWR VPWR hold359/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4582__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_754 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5536__A2 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3547__A1 _6926_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3547__B2 _7294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6497__B1 _6495_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_50_csclk _7496_/CLK VGND VGND VPWR VPWR _7478_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6249__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3661__B _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4249__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6264__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4773__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6760_ _7060_/Q _6447_/C _6651_/C _6419_/A _7161_/Q VGND VGND VPWR VPWR _6760_/X
+ sky130_fd_sc_hd__a32o_1
X_3972_ _7177_/Q hold56/A _5619_/B _3647_/X _7167_/Q VGND VGND VPWR VPWR _3972_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_128_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5711_ _5999_/A1 _5711_/A1 _5712_/S VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5100__C _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6691_ _7002_/Q _6419_/D _6421_/X _7007_/Q VGND VGND VPWR VPWR _6691_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5808__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5642_ _5642_/A0 _5805_/A1 _5642_/S VGND VGND VPWR VPWR _5642_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5573_ _5231_/B _5573_/B _5573_/C _5573_/D VGND VGND VPWR VPWR _5574_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7312_ _7582_/CLK _7312_/D fanout584/X VGND VGND VPWR VPWR _7312_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_143_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold202 hold202/A VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4524_ _4524_/A0 _5914_/A1 _4526_/S VGND VGND VPWR VPWR _4524_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3555__C hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold213 _7481_/Q VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6488__B1 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7395_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold224 hold224/A VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold235 hold235/A VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold246 hold246/A VGND VGND VPWR VPWR _7442_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7243_ _7363_/CLK _7243_/D fanout575/X VGND VGND VPWR VPWR _7243_/Q sky130_fd_sc_hd__dfstp_4
X_4455_ _5830_/C _4491_/B _4455_/C hold47/X VGND VGND VPWR VPWR _4455_/X sky130_fd_sc_hd__and4_1
Xhold257 hold257/A VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_1_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold268 hold268/A VGND VGND VPWR VPWR hold268/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold279 _7207_/Q VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3406_ _7585_/Q VGND VGND VPWR VPWR _4099_/D sky130_fd_sc_hd__inv_2
X_4386_ _5951_/A1 _4386_/A1 _4387_/S VGND VGND VPWR VPWR _4386_/X sky130_fd_sc_hd__mux2_1
X_7174_ _7176_/CLK _7174_/D fanout588/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfstp_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _7464_/Q _6094_/A _6086_/X _6099_/X _7352_/Q VGND VGND VPWR VPWR _6125_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3710__B2 _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _7598_/Q _7597_/Q VGND VGND VPWR VPWR _6056_/X sky130_fd_sc_hd__and2b_4
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _5107_/A _5180_/B VGND VGND VPWR VPWR _5007_/Y sky130_fd_sc_hd__nand2_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _7024_/CLK _6958_/D fanout566/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_165_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6106__C _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5909_ _5954_/A1 _5909_/A1 _5910_/S VGND VGND VPWR VPWR _5909_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6889_ _4169_/B2 _6889_/D _6839_/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6403__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6715__A1 _6969_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5151__B1 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold780 _4508_/X VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4577__B _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold791 hold791/A VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3481__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6246__A3 _6073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2170 _7366_/Q VGND VGND VPWR VPWR hold394/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5454__A1 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input20_A mask_rev_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2181 hold889/X VGND VGND VPWR VPWR _5674_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6284__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2192 _5766_/X VGND VGND VPWR VPWR hold497/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1480 _7468_/Q VGND VGND VPWR VPWR hold179/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1491 hold55/X VGND VGND VPWR VPWR hold1491/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3768__A1 _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6706__B2 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3656__B _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6111__B_N _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4193__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput307 _4134_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
Xoutput318 hold1193/X VGND VGND VPWR VPWR hold1194/A sky130_fd_sc_hd__buf_6
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput329 hold1213/X VGND VGND VPWR VPWR hold1214/A sky130_fd_sc_hd__buf_6
XANTENNA__3672__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _5654_/A1 _5951_/A1 _4248_/S VGND VGND VPWR VPWR _4240_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5590__C _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4918__D _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4171_ _4178_/A _4171_/B VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__and2_1
XFILLER_0_184_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5445__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6642__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2591_A _7311_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6812_ _7109_/Q _6812_/A2 _6812_/B1 wire463/A _6811_/X VGND VGND VPWR VPWR _6812_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6743_ _7170_/Q _6408_/D _6421_/X _7009_/Q _6742_/X VGND VGND VPWR VPWR _6749_/C
+ sky130_fd_sc_hd__a221o_1
X_3955_ _7527_/Q _3529_/X _5776_/A _7383_/Q VGND VGND VPWR VPWR _3955_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4442__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6674_ _6957_/Q _6431_/Y _6775_/B1 VGND VGND VPWR VPWR _6674_/X sky130_fd_sc_hd__o21a_1
X_3886_ _7480_/Q _3535_/X _3673_/X _7198_/Q _3885_/X VGND VGND VPWR VPWR _3886_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5625_ _5625_/A0 _5647_/A0 _5629_/S VGND VGND VPWR VPWR _5625_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6173__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4184__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5556_ _5533_/Y _5539_/X _5555_/X VGND VGND VPWR VPWR _5556_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4507_ _4507_/A0 _5647_/A0 _4508_/S VGND VGND VPWR VPWR _4507_/X sky130_fd_sc_hd__mux2_1
X_5487_ _4801_/B _4801_/C _4768_/Y _5408_/Y _5153_/C VGND VGND VPWR VPWR _5488_/C
+ sky130_fd_sc_hd__o41a_1
X_7226_ _7231_/CLK _7226_/D _4128_/B VGND VGND VPWR VPWR _7226_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5133__B1 _4940_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4438_ _4438_/A0 hold61/X _4439_/S VGND VGND VPWR VPWR _4438_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout501 _5902_/B VGND VGND VPWR VPWR _5640_/D sky130_fd_sc_hd__buf_12
XANTENNA__5684__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout512 _3444_/Y VGND VGND VPWR VPWR _6116_/B sky130_fd_sc_hd__buf_12
Xfanout523 _7590_/Q VGND VGND VPWR VPWR _6119_/B sky130_fd_sc_hd__clkbuf_8
X_7157_ _7268_/CLK _7157_/D _6871_/A VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfrtp_4
X_4369_ _4369_/A0 _5754_/A1 _4369_/S VGND VGND VPWR VPWR _4369_/X sky130_fd_sc_hd__mux2_1
Xfanout567 fanout569/X VGND VGND VPWR VPWR fanout567/X sky130_fd_sc_hd__buf_12
X_6108_ _6104_/X _6105_/X _6107_/X _6121_/C VGND VGND VPWR VPWR _6108_/X sky130_fd_sc_hd__o31a_1
Xfanout578 fanout587/X VGND VGND VPWR VPWR fanout578/X sky130_fd_sc_hd__buf_6
XANTENNA__4858__A_N _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7088_ _7513_/CLK _7088_/D fanout600/X VGND VGND VPWR VPWR _7667_/A sky130_fd_sc_hd__dfrtp_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 fanout606/X VGND VGND VPWR VPWR fanout589/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__6633__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6039_ _6121_/C _6038_/X _6037_/X VGND VGND VPWR VPWR _7592_/D sky130_fd_sc_hd__o21ai_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input68_A mgmt_gpio_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_4__f_wb_clk_i clkbuf_3_2_0_wb_clk_i/X VGND VGND VPWR VPWR _7623_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6219__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3989__A1 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5866__B _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4770__B _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3667__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 _6749_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _7570_/Q _5983_/A _5992_/C _5643_/A input64/X VGND VGND VPWR VPWR _3740_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3610__B1 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6155__A2 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3671_ hold36/X _4388_/B _5659_/B VGND VGND VPWR VPWR _5634_/A sky130_fd_sc_hd__and3_4
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5410_ _5410_/A _5410_/B _5410_/C VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6390_ _7020_/Q _6120_/X _6386_/X _6387_/X _6389_/X VGND VGND VPWR VPWR _6397_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_113_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5341_ _5180_/B _5058_/C _5202_/B VGND VGND VPWR VPWR _5343_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_112_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4929__C _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6458__A3 _6645_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5272_ _4709_/Y _4798_/Y _4946_/Y _4789_/Y _5271_/X VGND VGND VPWR VPWR _5272_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5666__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7011_ _7211_/CLK _7011_/D fanout572/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2906 _5958_/X VGND VGND VPWR VPWR hold2906/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4223_ _4254_/A0 _5987_/A1 _4231_/S VGND VGND VPWR VPWR _4223_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2917 _6968_/Q VGND VGND VPWR VPWR hold2917/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2928 _4384_/X VGND VGND VPWR VPWR hold2928/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2939 _7648_/A VGND VGND VPWR VPWR hold2939/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4154_ _4153_/X input38/X _6898_/Q VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3692__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4085_ _6895_/Q _6879_/Q _6839_/B VGND VGND VPWR VPWR _4178_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_176_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5776__B hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3466__B1_N _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4987_ _5339_/D _5183_/A _5138_/D _5339_/C VGND VGND VPWR VPWR _5041_/C sky130_fd_sc_hd__nand4_1
XANTENNA__6394__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3577__A _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6726_ _6725_/X _6726_/A1 _6751_/S VGND VGND VPWR VPWR _6726_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout422_A _6106_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3938_ _7243_/Q _4551_/A _3485_/X _4551_/C _3937_/X VGND VGND VPWR VPWR _3938_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_160_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6657_ _7132_/Q _6409_/X _6420_/B _6988_/Q _6655_/X VGND VGND VPWR VPWR _6657_/X
+ sky130_fd_sc_hd__a221o_1
X_3869_ _7148_/Q _3652_/X _3654_/X _7118_/Q _3859_/X VGND VGND VPWR VPWR _3869_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4157__A1 _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5608_ _5608_/A0 _5754_/A1 _5611_/S VGND VGND VPWR VPWR _5608_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6588_ _7460_/Q _6463_/A _6771_/A3 _6463_/X _7428_/Q VGND VGND VPWR VPWR _6588_/X
+ sky130_fd_sc_hd__a32o_1
X_5539_ _5488_/Y _5539_/B _5568_/B VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_169_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7209_ _7212_/CLK _7209_/D fanout573/X VGND VGND VPWR VPWR _7209_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout353 _6573_/S VGND VGND VPWR VPWR _6777_/S sky130_fd_sc_hd__buf_12
Xfanout375 _5603_/B VGND VGND VPWR VPWR _5632_/B sky130_fd_sc_hd__buf_12
Xfanout386 hold281/X VGND VGND VPWR VPWR _5587_/C sky130_fd_sc_hd__buf_8
XANTENNA__6606__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3683__A3 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout397 _5339_/A VGND VGND VPWR VPWR _5183_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__4574__C _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input122_A wb_adr_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4632__A2 _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5686__B hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6385__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6137__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5906__S _5910_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _4177_/B sky130_fd_sc_hd__buf_6
Xmax_cap509 _3856_/A VGND VGND VPWR VPWR _3923_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3653__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4608__C1 _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2018_A _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6612__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4084__B1 _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5820__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4910_ _4856_/A _5399_/A _4929_/A _5058_/D VGND VGND VPWR VPWR _4928_/B sky130_fd_sc_hd__and4b_2
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5890_ _5890_/A0 _5998_/A1 _5892_/S VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5596__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4841_ _4841_/A _4841_/B _4841_/C VGND VGND VPWR VPWR _4851_/A sky130_fd_sc_hd__nor3_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6376__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5584__A0 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7560_ _7560_/CLK _7560_/D fanout599/X VGND VGND VPWR VPWR _7560_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_184_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4772_ _4772_/A _4786_/C _4797_/B VGND VGND VPWR VPWR _4775_/C sky130_fd_sc_hd__and3_4
XANTENNA__3729__A4 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6511_ _7361_/Q _6462_/X _6502_/X _6506_/X _6510_/X VGND VGND VPWR VPWR _6511_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_hold76_A hold76/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3723_ _6992_/Q _5731_/B _5623_/B _3531_/X _7339_/Q VGND VGND VPWR VPWR _3723_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6128__A2 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7491_ _7560_/CLK _7491_/D fanout599/X VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_132_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5816__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4139__A1 input89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6442_ _7495_/Q _6600_/B _6651_/C _6422_/X _7287_/Q VGND VGND VPWR VPWR _6442_/X
+ sky130_fd_sc_hd__a32o_1
X_3654_ _5830_/C _4491_/B _4388_/B VGND VGND VPWR VPWR _3654_/X sky130_fd_sc_hd__and3_2
XFILLER_0_130_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5887__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6373_ _7145_/Q _6144_/C _6097_/B _6144_/B VGND VGND VPWR VPWR _6373_/X sky130_fd_sc_hd__o211a_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3585_ _7285_/Q _3590_/C _5659_/B _5857_/A _7461_/Q VGND VGND VPWR VPWR _3585_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3563__C _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5324_ _5324_/A _5324_/B VGND VGND VPWR VPWR _5340_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_100_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2703 _7056_/Q VGND VGND VPWR VPWR hold2703/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4956__A _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5255_ _4743_/A _4747_/B _5073_/B _4601_/Y VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__o31a_4
XANTENNA__6300__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2714 hold829/X VGND VGND VPWR VPWR _4520_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5103__A3 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3860__A _7183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2725 _4387_/X VGND VGND VPWR VPWR hold812/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2736 _5660_/X VGND VGND VPWR VPWR hold2736/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4206_ _4206_/A0 _5950_/A1 _4211_/S VGND VGND VPWR VPWR _4206_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4311__A1 _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2747 _4526_/X VGND VGND VPWR VPWR hold816/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5186_ _5038_/B _5180_/B _5030_/C _5026_/A VGND VGND VPWR VPWR _5186_/X sky130_fd_sc_hd__a31o_1
Xhold2758 _7116_/Q VGND VGND VPWR VPWR hold852/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2769 hold2769/A VGND VGND VPWR VPWR hold2769/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4167__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4137_ _7073_/Q _4136_/Y _3996_/A VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__o21a_1
XANTENNA_fanout372_A _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6603__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4068_ _4098_/A1 _4062_/B _4062_/Y _4076_/B _4067_/Y VGND VGND VPWR VPWR _6890_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5811__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4691__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5024__C1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6367__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4378__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_846 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3738__C _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6709_ _7134_/Q _6409_/X _6422_/X _6964_/Q _6708_/X VGND VGND VPWR VPWR _6709_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5726__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5327__B1 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5878__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3889__B1 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4569__C _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3473__C _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4866__A _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3813__B1 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4369__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__C _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output291_A _6925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_838 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire540 _4715_/Y VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3592__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5869__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold609 hold609/A VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3664__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6530__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4479__C _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4541__A1 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__B2 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5040_ _5158_/A _5339_/D _5183_/A _5339_/C VGND VGND VPWR VPWR _5041_/B sky130_fd_sc_hd__nand4_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1309 hold3133/X VGND VGND VPWR VPWR hold3134/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7391__SET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4926__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_192_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6991_ _7024_/CLK _6991_/D fanout566/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6597__A2 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5942_ _5942_/A0 _5996_/A1 hold23/X VGND VGND VPWR VPWR _5942_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3804__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6349__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5873_ _5873_/A0 hold61/X _5874_/S VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7612_ _7627_/CLK _7612_/D fanout566/X VGND VGND VPWR VPWR _7612_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3558__C _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4824_ _4824_/A _5531_/D _4824_/C _5531_/C VGND VGND VPWR VPWR _4830_/C sky130_fd_sc_hd__nand4_1
XFILLER_0_158_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7543_ _7551_/CLK _7543_/D fanout595/X VGND VGND VPWR VPWR _7543_/Q sky130_fd_sc_hd__dfstp_2
X_4755_ _4755_/A _5138_/B _4755_/C _5005_/A VGND VGND VPWR VPWR _4755_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_172_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3706_ _7507_/Q _3526_/X _3535_/X _7483_/Q _3705_/X VGND VGND VPWR VPWR _3706_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__3583__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7474_ _7522_/CLK _7474_/D fanout603/X VGND VGND VPWR VPWR _7474_/Q sky130_fd_sc_hd__dfrtp_4
X_4686_ _5138_/B _4687_/B _4687_/C VGND VGND VPWR VPWR _5410_/A sky130_fd_sc_hd__and3_4
XFILLER_0_31_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6425_ _6455_/B _6434_/B _6459_/B VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and3_4
X_3637_ _4551_/A _4491_/A _5992_/C VGND VGND VPWR VPWR _5643_/A sky130_fd_sc_hd__and3_4
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4532__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6356_ _7069_/Q _6110_/A _6332_/C _6075_/X _7165_/Q VGND VGND VPWR VPWR _6356_/X
+ sky130_fd_sc_hd__a32o_1
X_3568_ _3568_/A _3568_/B _3568_/C _3568_/D VGND VGND VPWR VPWR _3570_/C sky130_fd_sc_hd__nor4_2
Xhold3201 _7625_/Q VGND VGND VPWR VPWR _6751_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3212 _6625_/X VGND VGND VPWR VPWR _7621_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5307_ _5297_/A _5404_/C _5410_/B _5086_/B _4755_/C VGND VGND VPWR VPWR _5308_/C
+ sky130_fd_sc_hd__a32o_1
Xhold3223 _4047_/X VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3234 _7614_/Q VGND VGND VPWR VPWR _6401_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6287_ _6962_/Q _6144_/A _6136_/C _6379_/B1 _7122_/Q VGND VGND VPWR VPWR _6287_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2500 hold971/X VGND VGND VPWR VPWR _4263_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3245 _7601_/Q VGND VGND VPWR VPWR _6066_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout587_A fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3499_ _7502_/Q _5902_/A _3498_/X _7382_/Q _3495_/X VGND VGND VPWR VPWR _3524_/A
+ sky130_fd_sc_hd__a221o_1
Xhold3256 _6892_/Q VGND VGND VPWR VPWR _4064_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2511 _7002_/Q VGND VGND VPWR VPWR hold668/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__A1 _7001_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2522 hold686/X VGND VGND VPWR VPWR _5751_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3267 _6893_/Q VGND VGND VPWR VPWR _4057_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__B2 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2533 _7158_/Q VGND VGND VPWR VPWR hold690/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5238_ _5222_/A _5453_/A _5453_/B _4932_/X VGND VGND VPWR VPWR _5238_/X sky130_fd_sc_hd__a31o_1
Xhold3278 _7073_/Q VGND VGND VPWR VPWR _4124_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2544 hold660/X VGND VGND VPWR VPWR _4193_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2555 _7501_/Q VGND VGND VPWR VPWR hold777/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1810 hold116/X VGND VGND VPWR VPWR _5936_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2566 _7389_/Q VGND VGND VPWR VPWR hold793/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4599__A_N _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1821 hold304/X VGND VGND VPWR VPWR _5986_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4836__D _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1832 hold471/X VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2577 hold803/X VGND VGND VPWR VPWR _5972_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2588 _7424_/Q VGND VGND VPWR VPWR hold712/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5169_ _4672_/X _4956_/B _4980_/X _4692_/Y _4814_/Y VGND VGND VPWR VPWR _5169_/X
+ sky130_fd_sc_hd__o32a_1
Xhold1843 hold300/X VGND VGND VPWR VPWR _5861_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6037__A1 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1854 _4268_/X VGND VGND VPWR VPWR hold457/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2599 hold2599/A VGND VGND VPWR VPWR _5922_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6109__C _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1865 hold350/X VGND VGND VPWR VPWR _5933_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1876 _5859_/X VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1887 hold512/X VGND VGND VPWR VPWR _4306_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1898 _7321_/Q VGND VGND VPWR VPWR hold432/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6588__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5796__A0 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1771_A _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_191_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6760__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3574__A2 _5911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6512__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5720__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4523__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input50_A mgmt_gpio_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3877__A3 _5603_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6276__B2 _7406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3931__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4287__A0 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output304_A _4167_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5251__A2 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6035__B _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3801__A3 _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6200__A1 _7467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6200__B2 _7515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3675__A hold36/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4540_ _4540_/A0 _5714_/A0 hold57/X VGND VGND VPWR VPWR _4540_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold406 hold406/A VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4471_ _5852_/A0 _4471_/A1 _4472_/S VGND VGND VPWR VPWR _4471_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold417 _5585_/X VGND VGND VPWR VPWR _7212_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold428 hold428/A VGND VGND VPWR VPWR hold428/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold439 hold439/A VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6210_ _7419_/Q _6072_/X _6099_/X _7355_/Q _6209_/X VGND VGND VPWR VPWR _6210_/X
+ sky130_fd_sc_hd__a221o_1
X_3422_ _7466_/Q VGND VGND VPWR VPWR _3422_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4514__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7190_ _7190_/CLK _7190_/D fanout587/X VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _7512_/Q _6094_/A _6317_/C _6110_/X _7432_/Q VGND VGND VPWR VPWR _6141_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2517_A _7299_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6110_/A _6072_/B _6144_/B VGND VGND VPWR VPWR _6072_/X sky130_fd_sc_hd__and3_4
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 hold2658/X VGND VGND VPWR VPWR hold2659/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 hold2962/X VGND VGND VPWR VPWR hold2963/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5023_ _5023_/A _5023_/B VGND VGND VPWR VPWR _5025_/A sky130_fd_sc_hd__nor2_1
Xhold1128 hold2980/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1139 hold2703/X VGND VGND VPWR VPWR hold2704/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_178_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5778__A0 hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4445__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6974_ _7630_/CLK _6974_/D VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5242__A2 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3569__B _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5925_ _5997_/A1 _5925_/A1 _5928_/S VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5856_ _5991_/A1 _5856_/A1 _5856_/S VGND VGND VPWR VPWR _5856_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4807_ _5410_/A _4815_/B _5453_/B VGND VGND VPWR VPWR _4809_/A sky130_fd_sc_hd__and3_1
X_5787_ _5787_/A0 _5940_/A1 _5793_/S VGND VGND VPWR VPWR _5787_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6742__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7526_ _7572_/CLK hold26/X fanout596/X VGND VGND VPWR VPWR _7526_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_160_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4738_ _4706_/Y _4712_/Y _4734_/Y _4737_/Y _4723_/Y VGND VGND VPWR VPWR _4738_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout502_A hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7457_ _7457_/CLK _7457_/D fanout586/X VGND VGND VPWR VPWR _7457_/Q sky130_fd_sc_hd__dfrtp_2
X_4669_ _4570_/Y _4667_/B _4740_/D VGND VGND VPWR VPWR _4669_/X sky130_fd_sc_hd__o21a_4
XANTENNA__6111__D _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6408_ _6408_/A _6408_/B _6408_/C _6408_/D VGND VGND VPWR VPWR _6431_/A sky130_fd_sc_hd__nor4_4
XANTENNA__4505__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold940 hold940/A VGND VGND VPWR VPWR _7232_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7388_ _7577_/CLK _7388_/D fanout583/X VGND VGND VPWR VPWR _7388_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold951 hold951/A VGND VGND VPWR VPWR hold951/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold962 _4355_/X VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold973 hold973/A VGND VGND VPWR VPWR hold973/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6339_ _6335_/X _6336_/X _6338_/X _6121_/C VGND VGND VPWR VPWR _6339_/X sky130_fd_sc_hd__o31a_1
Xhold984 _4452_/X VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold995 hold995/A VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3020 hold3020/A VGND VGND VPWR VPWR _4360_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3031 _7239_/Q VGND VGND VPWR VPWR hold787/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3042 _4264_/X VGND VGND VPWR VPWR hold760/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4847__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3053 _6992_/Q VGND VGND VPWR VPWR hold745/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold282_A _5587_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3064 _7162_/Q VGND VGND VPWR VPWR hold3064/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2330 hold965/X VGND VGND VPWR VPWR _5782_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3075 hold3075/A VGND VGND VPWR VPWR _5858_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3086 _7016_/Q VGND VGND VPWR VPWR hold3086/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2341 _7420_/Q VGND VGND VPWR VPWR hold979/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2352 _5664_/X VGND VGND VPWR VPWR hold101/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3097 _5957_/X VGND VGND VPWR VPWR hold3097/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2363 hold917/X VGND VGND VPWR VPWR _4519_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2374 _7033_/Q VGND VGND VPWR VPWR hold907/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1640 _7159_/Q VGND VGND VPWR VPWR hold340/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2385 _7042_/Q VGND VGND VPWR VPWR hold616/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1651 hold374/X VGND VGND VPWR VPWR _4403_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2396 _7396_/Q VGND VGND VPWR VPWR hold985/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1662 hold60/X VGND VGND VPWR VPWR hold1662/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1673 _3463_/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1684 hold338/X VGND VGND VPWR VPWR _5863_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1695 hold359/X VGND VGND VPWR VPWR _7340_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4582__C _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5040__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5233__A2 _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input98_A usr2_vdd_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6194__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6733__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3547__A2 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3661__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4773__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3971_ _7209_/Q _5581_/A _3962_/X _3965_/X _3970_/X VGND VGND VPWR VPWR _3988_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_174_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5710_ _5953_/A1 _5710_/A1 _5712_/S VGND VGND VPWR VPWR _5710_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6690_ _7193_/Q _6443_/X _6468_/X _7143_/Q _6689_/X VGND VGND VPWR VPWR _6697_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5641_ _5641_/A0 _5948_/A1 _5642_/S VGND VGND VPWR VPWR _5641_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6185__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5932__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2467_A _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5572_ _5572_/A _5572_/B _5572_/C VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__and3_1
XFILLER_0_127_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7311_ _7577_/CLK _7311_/D fanout584/X VGND VGND VPWR VPWR _7311_/Q sky130_fd_sc_hd__dfstp_4
X_4523_ _4523_/A0 _5583_/A0 _4526_/S VGND VGND VPWR VPWR _4523_/X sky130_fd_sc_hd__mux2_1
Xhold203 hold203/A VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold214 hold214/A VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5824__S _5829_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7242_ _7363_/CLK _7242_/D fanout575/X VGND VGND VPWR VPWR _7242_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6488__B2 _7328_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold225 hold225/A VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold236 hold236/A VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4454_ _4454_/A0 _5586_/A0 _4454_/S VGND VGND VPWR VPWR _4454_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4499__A0 _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold247 hold247/A VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold258 hold258/A VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold269 hold269/A VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3405_ _7306_/Q VGND VGND VPWR VPWR _3405_/Y sky130_fd_sc_hd__inv_2
X_7173_ _7176_/CLK _7173_/D fanout588/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4385_ _5815_/A1 _4385_/A1 _4387_/S VGND VGND VPWR VPWR _4385_/X sky130_fd_sc_hd__mux2_1
X_6124_ _6124_/A1 _6777_/S _6122_/Y _6123_/X VGND VGND VPWR VPWR _7602_/D sky130_fd_sc_hd__a22o_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3710__A2 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A1 _6051_/Y _6054_/X VGND VGND VPWR VPWR _7597_/D sky130_fd_sc_hd__a21bo_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6660__A1 _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5006_ _4605_/Y _5528_/A3 _5046_/A _4690_/Y VGND VGND VPWR VPWR _5006_/Y sky130_fd_sc_hd__o31ai_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__A2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _7024_/CLK _6957_/D fanout567/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3777__A2 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5908_ _5998_/A1 _5908_/A1 _5910_/S VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__mux2_1
X_6888_ _4169_/B2 _6888_/D _6838_/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6176__B1 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5839_ _5866_/B _5911_/A _5992_/D VGND VGND VPWR VPWR _5847_/S sky130_fd_sc_hd__and3_4
XANTENNA__6403__B _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6715__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5923__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_173_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7509_ _7565_/CLK _7509_/D fanout605/X VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5734__S _5739_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4858__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_3__f_wb_clk_i clkbuf_3_1_0_wb_clk_i/X VGND VGND VPWR VPWR _7586_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold770 hold770/A VGND VGND VPWR VPWR _7416_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold781 hold781/A VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold792 _5693_/X VGND VGND VPWR VPWR _7309_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input152_A wb_dat_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3701__A2 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2160 _4445_/X VGND VGND VPWR VPWR hold170/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2171 hold394/X VGND VGND VPWR VPWR _5757_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2182 _7278_/Q VGND VGND VPWR VPWR hold436/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2193 _7519_/Q VGND VGND VPWR VPWR hold614/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1470 _5670_/S VGND VGND VPWR VPWR _5676_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input13_A mask_rev_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1481 hold179/X VGND VGND VPWR VPWR _5872_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1492 _5884_/X VGND VGND VPWR VPWR _5892_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5909__S _5910_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__A2 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6706__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5509__A3 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3656__C _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6182__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5644__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput308 _4135_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
Xoutput319 hold1203/X VGND VGND VPWR VPWR hold1204/A sky130_fd_sc_hd__buf_6
XFILLER_0_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3940__A2 _5911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3672__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5142__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5590__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2048_A _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4170_ _4178_/A _7109_/Q VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__and2_1
XFILLER_0_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4784__A _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5445__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6811_ _7111_/Q _6811_/A2 _6811_/B1 _7110_/Q VGND VGND VPWR VPWR _6811_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5819__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6742_ _7069_/Q _6463_/A _6441_/X _6443_/X _7195_/Q VGND VGND VPWR VPWR _6742_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3954_ _7511_/Q _5920_/A _4533_/A _7182_/Q _3953_/X VGND VGND VPWR VPWR _3954_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6158__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6673_ _7182_/Q _6574_/B _6771_/A3 _6654_/X _6672_/X VGND VGND VPWR VPWR _6673_/X
+ sky130_fd_sc_hd__a311o_2
XFILLER_0_190_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3885_ _7392_/Q _5785_/A _5785_/B _3526_/X _7504_/Q VGND VGND VPWR VPWR _3885_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_hold2751_A _6923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5905__A0 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5624_ _5624_/A0 _5754_/A1 _5629_/S VGND VGND VPWR VPWR _5624_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_171_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5555_ _5504_/B _5551_/X _5572_/B _5550_/Y VGND VGND VPWR VPWR _5555_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_170_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4506_ _4506_/A0 _5815_/A1 _4508_/S VGND VGND VPWR VPWR _4506_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5486_ _5569_/A _5569_/B VGND VGND VPWR VPWR _5486_/Y sky130_fd_sc_hd__nand2_1
X_7225_ _7231_/CLK _7225_/D _4128_/B VGND VGND VPWR VPWR _7225_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5133__A1 _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4437_ _4437_/A0 _5998_/A1 _4439_/S VGND VGND VPWR VPWR _4437_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6330__B1 _6328_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout502 hold47/X VGND VGND VPWR VPWR _5902_/B sky130_fd_sc_hd__buf_12
Xfanout513 _6067_/A VGND VGND VPWR VPWR _6775_/B1 sky130_fd_sc_hd__buf_12
Xfanout524 hold2311/X VGND VGND VPWR VPWR _4429_/B sky130_fd_sc_hd__buf_12
X_7156_ _7156_/CLK _7156_/D fanout598/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_4
X_4368_ _4368_/A0 _5951_/A1 _4369_/S VGND VGND VPWR VPWR _4368_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3695__A1 _7467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout535 _5404_/D VGND VGND VPWR VPWR _5295_/C sky130_fd_sc_hd__buf_12
XANTENNA_input5_A mask_rev_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6107_ _7295_/Q _6136_/B _6136_/C _6379_/B1 _7391_/Q VGND VGND VPWR VPWR _6107_/X
+ sky130_fd_sc_hd__a32o_1
Xfanout568 fanout569/X VGND VGND VPWR VPWR fanout568/X sky130_fd_sc_hd__buf_6
X_7087_ _7513_/CLK _7087_/D fanout600/X VGND VGND VPWR VPWR _7666_/A sky130_fd_sc_hd__dfrtp_1
Xfanout579 fanout582/X VGND VGND VPWR VPWR fanout579/X sky130_fd_sc_hd__buf_12
X_4299_ _4302_/S _6789_/A2 _4298_/Y VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__o21ai_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _6051_/C _6929_/Q _6116_/C _6136_/C VGND VGND VPWR VPWR _6038_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6633__B2 _7294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5729__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5956__C hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7368__SET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6149__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1949_A _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_64_csclk _7496_/CLK VGND VGND VPWR VPWR _7489_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6164__A3 _7289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_39_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6321__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3686__A1 _7233_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3989__A2 _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7447_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6388__B1 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5866__C _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3667__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_172_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6043__B _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3670_ _4473_/A hold36/A _4388_/B VGND VGND VPWR VPWR _3670_/X sky130_fd_sc_hd__and3_2
XANTENNA__6155__A3 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_180_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5340_ _5340_/A _5340_/B _5423_/B _5340_/D VGND VGND VPWR VPWR _5343_/C sky130_fd_sc_hd__nand4_1
X_5271_ _5255_/X _4789_/Y _5473_/B _5269_/X VGND VGND VPWR VPWR _5271_/X sky130_fd_sc_hd__o211a_1
X_7010_ _7191_/CLK _7010_/D fanout573/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfrtp_4
X_4222_ _4222_/A0 _4221_/X _4232_/S VGND VGND VPWR VPWR _4222_/X sky130_fd_sc_hd__mux2_1
Xhold2907 _7560_/Q VGND VGND VPWR VPWR hold2907/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3677__A1 _7539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2918 hold2918/A VGND VGND VPWR VPWR _4273_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2929 _7113_/Q VGND VGND VPWR VPWR hold2929/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4153_ _6942_/Q _7221_/Q _6839_/B VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4084_ _6895_/Q _6879_/Q _6839_/B VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__o21a_2
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6379__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4986_ _5339_/A _5339_/C VGND VGND VPWR VPWR _4986_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4680__C _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3577__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6725_ _6715_/X _6717_/X _6724_/X _6431_/Y _6959_/Q VGND VGND VPWR VPWR _6725_/X
+ sky130_fd_sc_hd__o32a_1
X_3937_ _7311_/Q _5983_/A _3669_/C _3936_/X VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3601__A1 _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6656_ _7177_/Q _6058_/X _6457_/X _7061_/Q _6651_/X VGND VGND VPWR VPWR _6656_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout415_A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3868_ _7312_/Q _3521_/X _4231_/S input72/X _3867_/X VGND VGND VPWR VPWR _3868_/X
+ sky130_fd_sc_hd__a221o_1
X_5607_ _5607_/A0 _5647_/A0 _5611_/S VGND VGND VPWR VPWR _5607_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4157__A2 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6587_ _7300_/Q _6420_/A _6576_/X _6578_/X _6586_/X VGND VGND VPWR VPWR _6587_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6551__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3799_ _7441_/Q _4509_/A _5983_/A _4545_/A _7194_/Q VGND VGND VPWR VPWR _3799_/X
+ sky130_fd_sc_hd__a32o_1
X_5538_ _5538_/A _5538_/B _5538_/C VGND VGND VPWR VPWR _5568_/B sky130_fd_sc_hd__and3_1
XANTENNA__3904__A2 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5469_ _5070_/X _5468_/X _5260_/C VGND VGND VPWR VPWR _5469_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7208_ _7630_/CLK _7208_/D _6780_/B VGND VGND VPWR VPWR _7208_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__7267__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7139_ _7156_/CLK _7139_/D fanout598/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfstp_4
Xfanout354 hold55/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__buf_12
Xfanout376 _3514_/X VGND VGND VPWR VPWR _5603_/B sky130_fd_sc_hd__buf_12
XANTENNA__6606__A1 _7309_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout387 _5911_/A VGND VGND VPWR VPWR _5983_/A sky130_fd_sc_hd__buf_12
Xfanout398 _4932_/B VGND VGND VPWR VPWR _5339_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__4574__D _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A wb_adr_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3840__A1 _7184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3840__B2 _7154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6144__A _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5593__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6790__A0 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5983__A _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6137__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input80_A spi_sck VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_2
XFILLER_0_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6542__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4608__B1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4084__A1 _6895_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5596__C _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4840_ _4888_/B _5282_/A _5058_/D _4856_/A VGND VGND VPWR VPWR _5404_/D sky130_fd_sc_hd__and4b_4
XFILLER_0_169_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4771_ _4700_/Y _4717_/Y _4770_/Y _4766_/Y VGND VGND VPWR VPWR _4776_/B sky130_fd_sc_hd__o211ai_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6510_ _7537_/Q _6427_/A _6574_/B _6747_/C _6509_/X VGND VGND VPWR VPWR _6510_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__3595__B1 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3722_ _6961_/Q _3657_/X _3717_/X _3719_/X _3721_/X VGND VGND VPWR VPWR _3732_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7490_ _7510_/CLK _7490_/D fanout603/X VGND VGND VPWR VPWR _7490_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6441_ _6435_/B _7598_/Q _7597_/Q _6462_/D VGND VGND VPWR VPWR _6441_/X sky130_fd_sc_hd__and4bb_4
XFILLER_0_99_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3653_ hold36/X _4388_/B _4346_/C VGND VGND VPWR VPWR _4340_/A sky130_fd_sc_hd__and3_4
XANTENNA__6533__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6372_ _7180_/Q _6110_/A _6091_/X _6110_/X _7175_/Q VGND VGND VPWR VPWR _6372_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3584_ _7405_/Q _5794_/A _3565_/X _7469_/Q _3583_/X VGND VGND VPWR VPWR _3587_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5323_ _5183_/C _5260_/D _5339_/C _5342_/A _5339_/D VGND VGND VPWR VPWR _5324_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5832__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5254_ _4707_/Y _4709_/Y _4774_/Y _4946_/Y VGND VGND VPWR VPWR _5254_/X sky130_fd_sc_hd__o22a_1
Xhold2704 hold2704/A VGND VGND VPWR VPWR _4389_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2715 _7057_/Q VGND VGND VPWR VPWR hold2715/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4205_ _4205_/A0 _5805_/A1 _4211_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3860__B _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2726 _7015_/Q VGND VGND VPWR VPWR hold843/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4448__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2737 _7319_/Q VGND VGND VPWR VPWR hold2737/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4311__A2 _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5185_ _5185_/A _5185_/B _5185_/C VGND VGND VPWR VPWR _5185_/Y sky130_fd_sc_hd__nand3_1
Xhold2748 _7271_/Q VGND VGND VPWR VPWR hold2748/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_3_6_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_6_0_csclk/X sky130_fd_sc_hd__clkbuf_8
Xhold2759 hold852/X VGND VGND VPWR VPWR _4454_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4136_ _7075_/Q _7072_/Q VGND VGND VPWR VPWR _4136_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4862__A3 _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4067_ _6890_/Q _7071_/Q _4067_/C VGND VGND VPWR VPWR _4067_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4075__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5272__B1 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4691__B _4758_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4183__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4969_ _4873_/X _5528_/A3 _4672_/X _4679_/Y _7109_/Q VGND VGND VPWR VPWR _4969_/Y
+ sky130_fd_sc_hd__o41ai_4
XANTENNA__6772__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1382_A _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3586__B1 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6708_ _7038_/Q _6651_/B _6651_/C _6707_/X VGND VGND VPWR VPWR _6708_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_62_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5327__A1 _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6639_ _7350_/Q _6452_/X _6468_/X _7414_/Q _6638_/X VGND VGND VPWR VPWR _6647_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6524__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1647_A _7240_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4212__A _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3889__B2 _7328_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5027__B _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5742__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4866__B _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4585__C _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3510__B1 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4882__A _4932_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3813__B2 _7231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3498__A _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__B1 _5013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6358__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6763__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7424__SET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5318__A1 _4583_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6515__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output284_A _7242_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7487__SET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3664__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6818__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2030_A _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4057__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6990_ _7409_/CLK _6990_/D fanout577/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_189_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_8_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5941_ _5941_/A0 _5986_/A1 hold23/X VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3804__A1 _7521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4942__D _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5872_ _5872_/A0 _5998_/A1 _5874_/S VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5006__B1 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7611_ _7627_/CLK _7611_/D fanout566/X VGND VGND VPWR VPWR _7611_/Q sky130_fd_sc_hd__dfrtp_1
X_4823_ _5295_/A _4823_/B _4823_/C _5038_/A VGND VGND VPWR VPWR _4824_/C sky130_fd_sc_hd__nand4_1
XFILLER_0_29_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6754__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5827__S _5829_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4754_ _4803_/A _5297_/B VGND VGND VPWR VPWR _4760_/D sky130_fd_sc_hd__nand2_1
X_7542_ _7542_/CLK _7542_/D fanout581/X VGND VGND VPWR VPWR _7542_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_172_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3705_ _7045_/Q _4370_/A _3665_/X _7126_/Q VGND VGND VPWR VPWR _3705_/X sky130_fd_sc_hd__a22o_1
X_7473_ _7499_/CLK _7473_/D fanout577/X VGND VGND VPWR VPWR _7473_/Q sky130_fd_sc_hd__dfrtp_4
X_4685_ _4593_/A _4591_/Y _4593_/Y VGND VGND VPWR VPWR _4822_/D sky130_fd_sc_hd__o21ai_4
XFILLER_0_43_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3583__A3 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3636_ input8/X _3486_/X _3529_/X _7532_/Q _3635_/X VGND VGND VPWR VPWR _3642_/B
+ sky130_fd_sc_hd__a221o_1
X_6424_ _6427_/A _6455_/B _6424_/C VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__and3_4
XFILLER_0_113_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6355_ _6355_/A1 _4116_/X _6067_/X _6354_/X VGND VGND VPWR VPWR _6355_/X sky130_fd_sc_hd__o31a_1
X_3567_ _7334_/Q _5713_/A _3563_/X _3566_/X _3560_/X VGND VGND VPWR VPWR _3568_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6809__A1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3202 _7618_/Q VGND VGND VPWR VPWR _6572_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5306_ _5306_/A _5306_/B VGND VGND VPWR VPWR _5308_/B sky130_fd_sc_hd__nand2_1
Xhold3213 _7615_/Q VGND VGND VPWR VPWR _6473_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3224 hold51/A VGND VGND VPWR VPWR _4024_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6286_ _7011_/Q _6136_/B _6120_/B _6332_/B VGND VGND VPWR VPWR _6286_/X sky130_fd_sc_hd__a31o_1
Xhold3235 _6401_/X VGND VGND VPWR VPWR _7614_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_3498_ _4473_/A _5590_/A _5830_/C VGND VGND VPWR VPWR _3498_/X sky130_fd_sc_hd__and3_4
Xhold2501 _4263_/X VGND VGND VPWR VPWR hold972/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3246 _6066_/X VGND VGND VPWR VPWR _7601_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3590__B _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6285__A2 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2512 hold668/X VGND VGND VPWR VPWR _4324_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3257 _6903_/Q VGND VGND VPWR VPWR _4036_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5237_ _5208_/Y _5237_/B _5237_/C VGND VGND VPWR VPWR _5237_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA_fanout482_A _5735_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2523 _7022_/Q VGND VGND VPWR VPWR hold666/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3268 _6900_/Q VGND VGND VPWR VPWR _4044_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3279 _6879_/Q VGND VGND VPWR VPWR _4082_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2534 hold690/X VGND VGND VPWR VPWR _4505_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1800 hold344/X VGND VGND VPWR VPWR _5699_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2545 _7277_/Q VGND VGND VPWR VPWR hold755/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2556 hold777/X VGND VGND VPWR VPWR _5909_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1811 _7054_/Q VGND VGND VPWR VPWR hold372/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1822 _5986_/X VGND VGND VPWR VPWR hold305/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2567 hold793/X VGND VGND VPWR VPWR _5783_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5168_ _4849_/X _5061_/X _5167_/Y _5294_/A VGND VGND VPWR VPWR _5168_/X sky130_fd_sc_hd__o31a_1
Xhold2578 _5972_/X VGND VGND VPWR VPWR hold804/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1833 _6970_/Q VGND VGND VPWR VPWR hold326/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2589 hold712/X VGND VGND VPWR VPWR _5823_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1844 _5861_/X VGND VGND VPWR VPWR hold301/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1855 hold457/X VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4119_ _6751_/S _4107_/Y _4105_/Y _7256_/Q _6929_/Q VGND VGND VPWR VPWR _6931_/D
+ sky130_fd_sc_hd__a32o_1
Xhold1866 _7489_/Q VGND VGND VPWR VPWR hold426/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6109__D _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1877 _7425_/Q VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5099_ _4798_/Y _4960_/A _5098_/Y VGND VGND VPWR VPWR _5099_/Y sky130_fd_sc_hd__o21ai_1
Xhold1888 _6952_/Q VGND VGND VPWR VPWR hold404/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5245__B1 _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1899 hold432/X VGND VGND VPWR VPWR _5707_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6588__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6745__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__S _5739_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3559__B1 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1764_A _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6422__A _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6760__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3574__A3 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5038__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3484__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3731__B1 _3727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4596__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input43_A mgmt_gpio_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3931__D _3931_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6579__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5787__A1 _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5251__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4117__A _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6736__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5647__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6200__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4211__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3675__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4470_ _5914_/A1 _4470_/A1 _4472_/S VGND VGND VPWR VPWR _4470_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2078_A _7259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold407 hold407/A VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5199__A_N _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire393 _6411_/Y VGND VGND VPWR VPWR _6431_/B sky130_fd_sc_hd__clkbuf_2
Xhold418 hold418/A VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6503__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3421_ _7474_/Q VGND VGND VPWR VPWR _3421_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold429 hold429/A VGND VGND VPWR VPWR _7450_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6140_ _7416_/Q _6072_/X _6097_/X _7440_/Q _6139_/X VGND VGND VPWR VPWR _6140_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6267__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _7589_/Q _7588_/Q _6136_/C VGND VGND VPWR VPWR _6071_/X sky130_fd_sc_hd__and3b_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2412_A _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5138_/D _5180_/A _5216_/A VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__and3_1
Xhold1107 hold2993/X VGND VGND VPWR VPWR hold2994/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _4517_/X VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1129 hold2973/X VGND VGND VPWR VPWR hold2974/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_178_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6973_ _7630_/CLK _6973_/D VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3789__B1 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5924_ _5996_/A1 _5924_/A1 _5928_/S VGND VGND VPWR VPWR _5924_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3569__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4450__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5855_ hold61/X _5855_/A1 _5856_/S VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4806_ _5100_/A _5260_/B VGND VGND VPWR VPWR _4806_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__4202__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5786_ hold567/X hold464/X _5793_/S VGND VGND VPWR VPWR _5786_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6742__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7525_ _7572_/CLK _7525_/D fanout596/X VGND VGND VPWR VPWR _7525_/Q sky130_fd_sc_hd__dfrtp_4
X_4737_ _5100_/A _5079_/B VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__5950__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7456_ _7581_/CLK hold64/X fanout585/X VGND VGND VPWR VPWR _7456_/Q sky130_fd_sc_hd__dfstp_2
X_4668_ _4984_/B _4805_/B _4668_/C _4797_/B VGND VGND VPWR VPWR _4974_/C sky130_fd_sc_hd__nand4_4
XFILLER_0_160_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2__f_wb_clk_i clkbuf_3_1_0_wb_clk_i/X VGND VGND VPWR VPWR _6999_/CLK sky130_fd_sc_hd__clkbuf_16
X_3619_ _7614_/Q _7253_/Q _7255_/Q VGND VGND VPWR VPWR _3619_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_4_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6407_ _6427_/A _6574_/B _6747_/C VGND VGND VPWR VPWR _6408_/D sky130_fd_sc_hd__and3_4
XFILLER_0_101_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5702__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold930 _5953_/X VGND VGND VPWR VPWR _7540_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold941 hold941/A VGND VGND VPWR VPWR hold941/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4599_ _5282_/A _4888_/B VGND VGND VPWR VPWR _5073_/A sky130_fd_sc_hd__nand2b_4
X_7387_ _7575_/CLK _7387_/D fanout595/X VGND VGND VPWR VPWR _7387_/Q sky130_fd_sc_hd__dfrtp_4
Xhold952 _4350_/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold963 hold963/A VGND VGND VPWR VPWR hold963/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold974 _4307_/X VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6338_ _7013_/Q _6136_/B _6120_/B _6337_/X VGND VGND VPWR VPWR _6338_/X sky130_fd_sc_hd__a31o_1
Xhold3010 _7191_/Q VGND VGND VPWR VPWR hold773/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold985 hold985/A VGND VGND VPWR VPWR hold985/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold996 _5773_/X VGND VGND VPWR VPWR _7380_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3021 _7047_/Q VGND VGND VPWR VPWR hold3021/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3032 hold787/X VGND VGND VPWR VPWR _5608_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3043 _7010_/Q VGND VGND VPWR VPWR hold785/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3054 hold745/X VGND VGND VPWR VPWR _4308_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6269_ _7534_/Q _6094_/A _6091_/X _6121_/X _7310_/Q VGND VGND VPWR VPWR _6269_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4269__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3065 hold3065/A VGND VGND VPWR VPWR _4510_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2320 _4258_/X VGND VGND VPWR VPWR hold613/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2331 _7323_/Q VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3076 _7375_/Q VGND VGND VPWR VPWR hold3076/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3087 hold3087/A VGND VGND VPWR VPWR _4341_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2342 hold979/X VGND VGND VPWR VPWR _5818_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2353 _7505_/Q VGND VGND VPWR VPWR hold935/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3098 _7006_/Q VGND VGND VPWR VPWR hold3098/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2364 _7199_/Q VGND VGND VPWR VPWR hold947/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1630 _7189_/Q VGND VGND VPWR VPWR hold324/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2375 hold907/X VGND VGND VPWR VPWR _4361_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1641 hold340/X VGND VGND VPWR VPWR _4506_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2386 hold616/X VGND VGND VPWR VPWR _4372_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1652 _7008_/Q VGND VGND VPWR VPWR hold320/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2397 hold985/X VGND VGND VPWR VPWR _5791_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1663 hold1663/A VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6417__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1674 hold34/X VGND VGND VPWR VPWR _3505_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1685 _5863_/X VGND VGND VPWR VPWR hold339/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1696 _7369_/Q VGND VGND VPWR VPWR hold414/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5769__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_168_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6136__B _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4582__D _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4441__A1 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6718__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6194__A1 _7323_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6194__B2 _7339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5941__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4400__A _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6249__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5209__B1 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3970_ _7495_/Q _5902_/A _3969_/X _3931_/X _3968_/X VGND VGND VPWR VPWR _3970_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4432__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6709__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2195_A _7518_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5640_ _5722_/A _5640_/B _5640_/C _5640_/D VGND VGND VPWR VPWR _5642_/S sky130_fd_sc_hd__and4_1
XANTENNA__6185__A1 _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6185__B2 _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5571_ _5038_/B _5339_/B _5030_/C _5570_/X _5435_/D VGND VGND VPWR VPWR _5572_/C
+ sky130_fd_sc_hd__a311oi_2
XFILLER_0_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7310_ _7542_/CLK _7310_/D fanout581/X VGND VGND VPWR VPWR _7310_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4522_ _4522_/A0 _5840_/A1 _4526_/S VGND VGND VPWR VPWR _4522_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold204 hold204/A VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6488__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold215 hold215/A VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7241_ _7363_/CLK _7241_/D fanout575/X VGND VGND VPWR VPWR _7241_/Q sky130_fd_sc_hd__dfstp_2
Xhold226 hold226/A VGND VGND VPWR VPWR _7500_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4453_ _4453_/A0 _5852_/A0 _4454_/S VGND VGND VPWR VPWR _4453_/X sky130_fd_sc_hd__mux2_1
Xhold237 hold237/A VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_111_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold248 hold248/A VGND VGND VPWR VPWR _7506_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3404_ _5071_/A VGND VGND VPWR VPWR _5089_/B sky130_fd_sc_hd__inv_8
Xhold259 hold259/A VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4310__A _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7172_ _7176_/CLK _7172_/D fanout588/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_4
X_4384_ _5583_/A0 _4384_/A1 _4387_/S VGND VGND VPWR VPWR _4384_/X sky130_fd_sc_hd__mux2_1
X_6123_ _7279_/Q _6036_/Y _6775_/B1 _6931_/Q VGND VGND VPWR VPWR _6123_/X sky130_fd_sc_hd__o211a_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6050_/Y _6051_/C _7597_/Q _6019_/Y VGND VGND VPWR VPWR _6054_/X sky130_fd_sc_hd__a211o_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5005_/A _5005_/B _5005_/C VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__nand3_4
XANTENNA_hold2996_A _7363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6660__A2 _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4671__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6902__CLK _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__A3 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _6956_/CLK _6956_/D fanout604/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5907_ hold84/X _5907_/A1 _5910_/S VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__mux2_1
X_6887_ _4169_/B2 _6887_/D _6837_/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout612_A _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6176__A1 _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5838_ _5838_/A0 hold17/X _5838_/S VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6176__B2 _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6403__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5769_ _5769_/A0 _5985_/A1 _5775_/S VGND VGND VPWR VPWR _5769_/X sky130_fd_sc_hd__mux2_1
X_7508_ _7566_/CLK _7508_/D fanout603/X VGND VGND VPWR VPWR _7508_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6479__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7439_ _7505_/CLK _7439_/D fanout601/X VGND VGND VPWR VPWR _7439_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5687__A0 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold760 hold760/A VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5151__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold771 hold771/A VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold782 _5889_/X VGND VGND VPWR VPWR _7483_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold793 hold793/A VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5439__B1 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input145_A wb_dat_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2150 hold141/X VGND VGND VPWR VPWR _5853_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2161 _6939_/Q VGND VGND VPWR VPWR hold410/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_189_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2172 _5757_/X VGND VGND VPWR VPWR hold395/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2183 hold436/X VGND VGND VPWR VPWR _5658_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2194 hold614/X VGND VGND VPWR VPWR _5930_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1460 hold171/X VGND VGND VPWR VPWR _5926_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1471 _5671_/X VGND VGND VPWR VPWR hold198/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1482 _5872_/X VGND VGND VPWR VPWR hold180/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1493 _5887_/X VGND VGND VPWR VPWR hold214/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7644__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4414__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4965__A2 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5914__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput309 _7672_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
XFILLER_0_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3672__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5142__A2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6642__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5850__A0 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5387__A_N _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2208_A _7310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6810_ _6809_/X _6810_/A1 _6822_/S VGND VGND VPWR VPWR _7640_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4405__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6741_ _7160_/Q _6419_/A _6447_/X _7185_/Q _6740_/X VGND VGND VPWR VPWR _6749_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3953_ _7132_/Q _5785_/A _5619_/B _3506_/X _7351_/Q VGND VGND VPWR VPWR _3953_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4950__D _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6158__A1 _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6158__B2 _7393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6672_ _6962_/Q _6422_/X _6656_/X _6666_/X _6671_/X VGND VGND VPWR VPWR _6672_/X
+ sky130_fd_sc_hd__a2111o_1
X_3884_ _7528_/Q _3529_/X _3661_/X _7032_/Q _3883_/X VGND VGND VPWR VPWR _3884_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5623_ _5640_/C _5623_/B _5640_/D VGND VGND VPWR VPWR _5629_/S sky130_fd_sc_hd__and3_4
XFILLER_0_171_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5835__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3916__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5381__A2 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5554_ _5554_/A _5554_/B _5554_/C VGND VGND VPWR VPWR _5572_/B sky130_fd_sc_hd__and3_1
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_170_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3863__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4505_ _4505_/A0 _5805_/A1 _4508_/S VGND VGND VPWR VPWR _4505_/X sky130_fd_sc_hd__mux2_1
X_5485_ _5408_/Y _4713_/X _5143_/C _5303_/A VGND VGND VPWR VPWR _5569_/B sky130_fd_sc_hd__o211a_1
XANTENNA__5669__A0 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4436_ _4436_/A0 _5979_/A0 _4439_/S VGND VGND VPWR VPWR _4436_/X sky130_fd_sc_hd__mux2_1
X_7224_ _7231_/CLK _7224_/D _4128_/B VGND VGND VPWR VPWR _7224_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6330__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5133__A2 _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4341__A0 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout503 hold47/X VGND VGND VPWR VPWR _4551_/D sky130_fd_sc_hd__buf_12
Xfanout514 _7596_/Q VGND VGND VPWR VPWR _6462_/D sky130_fd_sc_hd__clkbuf_16
X_4367_ _4367_/A0 _5950_/A1 _4369_/S VGND VGND VPWR VPWR _4367_/X sky130_fd_sc_hd__mux2_1
X_7155_ _7156_/CLK _7155_/D _6833_/A VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout525 hold3283/X VGND VGND VPWR VPWR _4025_/A sky130_fd_sc_hd__clkbuf_16
X_6106_ _6119_/A _6106_/B _6136_/B VGND VGND VPWR VPWR _6106_/X sky130_fd_sc_hd__and3_4
XFILLER_0_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7086_ _7513_/CLK _7086_/D fanout600/X VGND VGND VPWR VPWR _7665_/A sky130_fd_sc_hd__dfrtp_1
Xfanout558 _4626_/B VGND VGND VPWR VPWR _5038_/A sky130_fd_sc_hd__buf_12
Xfanout569 fanout587/X VGND VGND VPWR VPWR fanout569/X sky130_fd_sc_hd__buf_12
X_4298_ _4302_/S _4298_/B VGND VGND VPWR VPWR _4298_/Y sky130_fd_sc_hd__nand2_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6633__A2 _6404_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6037_ _6036_/Y _6051_/C _6019_/Y VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__a21o_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6939_ _6956_/CLK _6939_/D fanout603/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6149__A1 _7529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6554__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5745__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3907__B1 _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_csclk _4169_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__4134__A_N _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5046__A _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3492__C _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6321__A1 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold590 hold590/A VGND VGND VPWR VPWR hold590/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4885__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3686__A2 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4635__A1 _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3989__A3 _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1290 hold3045/X VGND VGND VPWR VPWR hold3046/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4399__A0 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3667__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3610__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5899__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5270_ _4698_/Y _5563_/A1 _4946_/Y _4789_/Y _4709_/Y VGND VGND VPWR VPWR _5473_/B
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4323__A0 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4221_ _4253_/A0 _5986_/A1 _4231_/S VGND VGND VPWR VPWR _4221_/X sky130_fd_sc_hd__mux2_1
Xhold2908 hold2908/A VGND VGND VPWR VPWR _5976_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3677__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2919 _7568_/Q VGND VGND VPWR VPWR hold2919/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4874__B2 _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4152_ _6947_/Q input77/X _4173_/B VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__mux2_8
XANTENNA__6076__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6615__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4083_ _7600_/Q _7250_/Q _7255_/Q VGND VGND VPWR VPWR _4117_/B sky130_fd_sc_hd__mux2_8
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4985_ _5328_/A _5328_/B _5339_/C VGND VGND VPWR VPWR _5030_/C sky130_fd_sc_hd__and3_4
XFILLER_0_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3577__C _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6724_ _6431_/A _6431_/B _6431_/C _6723_/X VGND VGND VPWR VPWR _6724_/X sky130_fd_sc_hd__a31o_1
X_3936_ _7543_/Q _4491_/B _4212_/A _3654_/X _7117_/Q VGND VGND VPWR VPWR _3936_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_6655_ _7066_/Q _6463_/A _6441_/X _6425_/X _7016_/Q VGND VGND VPWR VPWR _6655_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3867_ _7336_/Q _3531_/X _3667_/X _7022_/Q _3863_/X VGND VGND VPWR VPWR _3867_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_33_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5606_ _5606_/A0 _5950_/A1 _5611_/S VGND VGND VPWR VPWR _5606_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4157__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6551__A1 _7331_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6586_ _7540_/Q _6408_/D _6582_/X _6585_/X VGND VGND VPWR VPWR _6586_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6551__B2 _7347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3798_ _7569_/Q _5983_/A _5965_/A _3654_/X _7119_/Q VGND VGND VPWR VPWR _3798_/X
+ sky130_fd_sc_hd__a32o_1
X_5537_ _4706_/Y _4735_/Y _4760_/D _5536_/Y VGND VGND VPWR VPWR _5538_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5468_ _5100_/A _5079_/B _4790_/B _5038_/A _5134_/A VGND VGND VPWR VPWR _5468_/X
+ sky130_fd_sc_hd__a32o_1
X_7207_ _7207_/CLK _7207_/D _6780_/B VGND VGND VPWR VPWR _7207_/Q sky130_fd_sc_hd__dfrtp_1
X_4419_ _4419_/A0 _4418_/X _4423_/S VGND VGND VPWR VPWR _4419_/X sky130_fd_sc_hd__mux2_1
X_5399_ _5399_/A _5399_/B _5399_/C _5399_/D VGND VGND VPWR VPWR _5481_/B sky130_fd_sc_hd__nand4_1
XFILLER_0_10_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7138_ _7447_/CLK _7138_/D fanout598/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout355 hold55/X VGND VGND VPWR VPWR _5947_/B sky130_fd_sc_hd__clkbuf_16
Xfanout366 _6873_/B VGND VGND VPWR VPWR _6869_/B sky130_fd_sc_hd__buf_6
Xfanout377 _4346_/C VGND VGND VPWR VPWR _5731_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__6606__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout388 _3933_/A VGND VGND VPWR VPWR _5785_/B sky130_fd_sc_hd__buf_12
X_7069_ _7190_/CLK _7069_/D _6871_/A VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4617__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1794_A _7554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4871__C _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7159__SET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_179_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input108_A wb_adr_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6144__B _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4250__C1 hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_18_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6542__A1 _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6542__B2 _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4599__B _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4553__A0 _5940_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input73_A pad_flash_io0_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4608__A1 _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4084__A2 _6879_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5596__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6230__B1 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4770_ _5387_/C _5113_/A _5404_/C _5410_/B VGND VGND VPWR VPWR _4770_/Y sky130_fd_sc_hd__nand4_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5893__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3595__B2 _7533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3721_ input16/X _3490_/X _5581_/A _7213_/Q _3720_/X VGND VGND VPWR VPWR _3721_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6440_ _7575_/Q _6427_/X _6432_/X _6439_/X _6430_/X VGND VGND VPWR VPWR _6440_/Y
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_0_125_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3652_ _4491_/A _4491_/B _4491_/C VGND VGND VPWR VPWR _3652_/X sky130_fd_sc_hd__and3_2
XANTENNA__6533__B2 _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6371_ _7044_/Q _6089_/X _6144_/C _7064_/Q _6100_/X VGND VGND VPWR VPWR _6371_/X
+ sky130_fd_sc_hd__a32o_1
X_3583_ _7525_/Q _5785_/B _5938_/C _4231_/S input41/X VGND VGND VPWR VPWR _3583_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_141_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3898__A2 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5322_ _5496_/B _5320_/X _5321_/X _5294_/Y VGND VGND VPWR VPWR _5322_/Y sky130_fd_sc_hd__a31oi_2
XANTENNA__6297__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5253_ _5107_/A _5282_/B wire529/X _5107_/X VGND VGND VPWR VPWR _5278_/D sky130_fd_sc_hd__a31oi_1
Xhold2705 _7435_/Q VGND VGND VPWR VPWR hold757/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4204_ _4204_/A0 _5948_/A1 _4211_/S VGND VGND VPWR VPWR _4204_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3860__C _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2716 hold2716/A VGND VGND VPWR VPWR _4390_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5184_ _4605_/Y _5528_/A3 _5046_/A _5183_/Y VGND VGND VPWR VPWR _5184_/X sky130_fd_sc_hd__o31a_1
Xhold2727 hold843/X VGND VGND VPWR VPWR _4339_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_139_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2738 hold2738/A VGND VGND VPWR VPWR _5705_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2749 hold2749/A VGND VGND VPWR VPWR _5651_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4135_ _6896_/Q _4135_/B VGND VGND VPWR VPWR _4135_/X sky130_fd_sc_hd__and2b_4
Xclkbuf_leaf_63_csclk _7496_/CLK VGND VGND VPWR VPWR _7457_/CLK sky130_fd_sc_hd__clkbuf_16
X_4066_ _6891_/Q _4098_/A1 _7071_/Q _4067_/C _4065_/Y VGND VGND VPWR VPWR _4066_/Y
+ sky130_fd_sc_hd__o41ai_1
XANTENNA__5272__A1 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4691__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3822__A2 hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6221__B1 _6090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4968_ _4873_/X _5528_/A3 _4672_/X _4679_/Y _7109_/Q VGND VGND VPWR VPWR _4968_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_136_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6707_ _7063_/Q _6574_/B _6441_/X _6058_/X _7179_/Q VGND VGND VPWR VPWR _6707_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3919_ _7304_/Q _5686_/A _3914_/X _3915_/X _3918_/X VGND VGND VPWR VPWR _3919_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_0_163_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4899_ _4667_/A _4608_/Y _4657_/C wire533/X _5213_/C VGND VGND VPWR VPWR _4899_/Y
+ sky130_fd_sc_hd__o2111ai_2
X_6638_ _7478_/Q _6424_/C _6441_/X _6443_/X _7454_/Q VGND VGND VPWR VPWR _6638_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5327__A2 _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6524__A1 _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6524__B2 _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4535__A0 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4212__B _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6569_ _6569_/A _6569_/B _6569_/C _6569_/D VGND VGND VPWR VPWR _6570_/C sky130_fd_sc_hd__nor4_2
XANTENNA__3889__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7505_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6288__B1 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4866__C _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7417__RESET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3510__B2 input33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6099__B_N _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4882__B _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5263__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3813__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3498__B _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5015__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5318__A2 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6515__B2 _7449_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6279__B1 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3453__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__A3 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7158__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5254__B2 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5940_ _5940_/A0 _5940_/A1 hold23/X VGND VGND VPWR VPWR _5940_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3804__A2 _5929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5871_ _5871_/A0 _5997_/A1 _5874_/S VGND VGND VPWR VPWR _5871_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5006__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6203__B1 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7610_ _7610_/CLK _7610_/D fanout568/X VGND VGND VPWR VPWR _7610_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4822_ _5138_/A _5138_/C _5138_/D _4822_/D VGND VGND VPWR VPWR _5531_/D sky130_fd_sc_hd__nand4_4
XFILLER_0_90_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7541_ _7542_/CLK _7541_/D fanout581/X VGND VGND VPWR VPWR _7541_/Q sky130_fd_sc_hd__dfrtp_2
X_4753_ _4778_/A _4767_/B _4753_/C VGND VGND VPWR VPWR _5297_/B sky130_fd_sc_hd__and3_2
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4313__A _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3704_ _6878_/Q _5875_/A _5632_/B _3703_/X VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_172_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7472_ _7499_/CLK _7472_/D fanout578/X VGND VGND VPWR VPWR _7472_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4684_ _4825_/A _4593_/A _4592_/X VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_160_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6423_ _6463_/A _6455_/B _6651_/B VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__and3_4
Xclkbuf_4_1__f_wb_clk_i clkbuf_3_0_0_wb_clk_i/X VGND VGND VPWR VPWR _7593_/CLK sky130_fd_sc_hd__clkbuf_16
X_3635_ _7492_/Q _5947_/B hold12/A _3565_/X _7468_/Q VGND VGND VPWR VPWR _3635_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6354_ _6751_/S _7611_/Q _6777_/S _6353_/X VGND VGND VPWR VPWR _6354_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_113_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3566_ _7366_/Q _5803_/A hold12/A _3565_/X _7470_/Q VGND VGND VPWR VPWR _3566_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3203 _6548_/X VGND VGND VPWR VPWR _7618_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3740__A1 _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5305_ _4716_/Y _4723_/Y _4978_/Y _4713_/X _5304_/X VGND VGND VPWR VPWR _5306_/B
+ sky130_fd_sc_hd__o221a_1
Xhold3214 _6473_/X VGND VGND VPWR VPWR _7615_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3740__B2 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3497_ _5722_/A _4449_/B _5947_/B VGND VGND VPWR VPWR _5902_/A sky130_fd_sc_hd__and3_4
X_6285_ _7001_/Q _6116_/C _6120_/B _6332_/C _7031_/Q VGND VGND VPWR VPWR _6285_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3225 _7072_/Q VGND VGND VPWR VPWR _4113_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3236 _7075_/Q VGND VGND VPWR VPWR _3403_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3247 _6898_/Q VGND VGND VPWR VPWR _4048_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2502 _6914_/Q VGND VGND VPWR VPWR hold959/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3590__C _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2513 _7408_/Q VGND VGND VPWR VPWR hold672/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3258 _6904_/Q VGND VGND VPWR VPWR _4033_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5236_ _4799_/C _4885_/X _4927_/B VGND VGND VPWR VPWR _5237_/C sky130_fd_sc_hd__a21oi_1
Xhold2524 hold666/X VGND VGND VPWR VPWR _4348_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3269 _7108_/Q VGND VGND VPWR VPWR _6827_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_166_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2535 _7493_/Q VGND VGND VPWR VPWR hold801/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1801 _5699_/X VGND VGND VPWR VPWR hold345/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2546 hold755/X VGND VGND VPWR VPWR _5657_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6690__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2557 _7461_/Q VGND VGND VPWR VPWR hold789/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4983__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1812 hold372/X VGND VGND VPWR VPWR _4386_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2568 _7541_/Q VGND VGND VPWR VPWR hold831/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1823 _7538_/Q VGND VGND VPWR VPWR hold380/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5167_ _5167_/A _5529_/A _5496_/B _5496_/A VGND VGND VPWR VPWR _5167_/Y sky130_fd_sc_hd__nand4_1
Xhold2579 _7437_/Q VGND VGND VPWR VPWR hold805/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout475_A hold2072/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1834 hold326/X VGND VGND VPWR VPWR _4275_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1845 _7465_/Q VGND VGND VPWR VPWR hold322/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_75_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1856 _7410_/Q VGND VGND VPWR VPWR hold342/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4118_ _4107_/A _6751_/S _6051_/C _4116_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__a211o_1
X_5098_ _4887_/B _5091_/A _4797_/X _5097_/Y VGND VGND VPWR VPWR _5098_/Y sky130_fd_sc_hd__a31oi_2
Xhold1867 hold426/X VGND VGND VPWR VPWR _5896_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1878 hold498/X VGND VGND VPWR VPWR _5824_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5245__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1889 hold404/X VGND VGND VPWR VPWR _4254_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6442__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4049_ _6908_/Q _7071_/Q _6910_/Q _6909_/Q VGND VGND VPWR VPWR _4050_/S sky130_fd_sc_hd__and4b_1
XFILLER_0_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6745__B2 _7155_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3559__A1 _7542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6422__B _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5181__B1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4877__B _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3731__A1 _4177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3040_A _6961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6276__A3 _6093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input36_A mgmt_gpio_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3495__B1 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__buf_12
XANTENNA__3798__A1 _7569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3798__B2 _7119_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4117__B _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6197__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6736__A1 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6200__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6332__B _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3675__C hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire350 _6102_/Y VGND VGND VPWR VPWR _6122_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold408 hold408/A VGND VGND VPWR VPWR hold408/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold419 _5584_/X VGND VGND VPWR VPWR _7211_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3420_ _7482_/Q VGND VGND VPWR VPWR _3420_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_111_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4787__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3722__A1 _6961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6332_/B _6119_/B _6116_/C _6112_/D VGND VGND VPWR VPWR _6070_/X sky130_fd_sc_hd__and4bb_4
XANTENNA__6267__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5475__A1 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A _5021_/B _5021_/C _5021_/D VGND VGND VPWR VPWR _5023_/B sky130_fd_sc_hd__nand4_1
Xhold1108 hold2995/X VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1119 hold2960/X VGND VGND VPWR VPWR hold2961/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6972_ _7206_/CLK _6972_/D VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3789__A1 _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5923_ _5986_/A1 _5923_/A1 _5928_/S VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5838__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5854_ _5998_/A1 _5854_/A1 _5856_/S VGND VGND VPWR VPWR _5854_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4805_ _4984_/B _4805_/B _5260_/B VGND VGND VPWR VPWR _5453_/B sky130_fd_sc_hd__and3_4
XFILLER_0_44_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5785_ _5785_/A _5785_/B _5992_/D VGND VGND VPWR VPWR _5793_/S sky130_fd_sc_hd__and3_4
X_7524_ _7572_/CLK _7524_/D fanout596/X VGND VGND VPWR VPWR _7524_/Q sky130_fd_sc_hd__dfrtp_4
X_4736_ _4795_/C _4740_/D _4909_/D VGND VGND VPWR VPWR _5074_/B sky130_fd_sc_hd__and3b_4
XFILLER_0_145_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7455_ _7487_/CLK _7455_/D fanout593/X VGND VGND VPWR VPWR _7455_/Q sky130_fd_sc_hd__dfstp_2
X_4667_ _4667_/A _4667_/B _4667_/C VGND VGND VPWR VPWR _4667_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_160_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6406_ _7594_/Q _7597_/Q _7598_/Q _6455_/B VGND VGND VPWR VPWR _6408_/C sky130_fd_sc_hd__and4bb_4
X_3618_ _7332_/Q _3933_/A _5731_/B _3521_/X _7316_/Q VGND VGND VPWR VPWR _3618_/X
+ sky130_fd_sc_hd__a32o_1
Xhold920 _4543_/X VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4697__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold931 hold931/A VGND VGND VPWR VPWR hold931/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7386_ _7575_/CLK _7386_/D fanout596/X VGND VGND VPWR VPWR _7386_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4598_ _5282_/A _4888_/B VGND VGND VPWR VPWR _5399_/A sky130_fd_sc_hd__and2b_4
Xhold942 _4458_/X VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3713__A1 _7291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold953 hold953/A VGND VGND VPWR VPWR hold953/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3713__B2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6337_ _6964_/Q _6144_/A _6136_/C _6379_/B1 _7124_/Q VGND VGND VPWR VPWR _6337_/X
+ sky130_fd_sc_hd__a32o_1
Xhold964 hold964/A VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout592_A fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3000 _5633_/X VGND VGND VPWR VPWR _7257_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold975 hold975/A VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3549_ _4551_/A _5992_/C _4388_/B VGND VGND VPWR VPWR _4422_/S sky130_fd_sc_hd__and3_4
XFILLER_0_177_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3011 hold773/X VGND VGND VPWR VPWR _4544_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold986 _5791_/X VGND VGND VPWR VPWR _7396_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3022 hold3022/A VGND VGND VPWR VPWR _4378_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3033 _7327_/Q VGND VGND VPWR VPWR hold3033/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold997 hold997/A VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_177_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3044 hold785/X VGND VGND VPWR VPWR _4333_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6268_ _7478_/Q _6032_/Y _6267_/X _6116_/B VGND VGND VPWR VPWR _6268_/X sky130_fd_sc_hd__a211o_1
Xhold2310 hold547/X VGND VGND VPWR VPWR _4439_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3055 _7146_/Q VGND VGND VPWR VPWR hold771/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5466__A1 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2321 _7320_/Q VGND VGND VPWR VPWR hold576/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3066 _4510_/X VGND VGND VPWR VPWR hold3066/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2332 hold98/X VGND VGND VPWR VPWR _5709_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6663__B1 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3077 hold3077/A VGND VGND VPWR VPWR _5768_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5219_ _4741_/Y _4886_/Y _4896_/Y _4903_/Y _5218_/Y VGND VGND VPWR VPWR _5219_/Y
+ sky130_fd_sc_hd__o2111ai_2
Xhold2343 _5818_/X VGND VGND VPWR VPWR hold980/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3088 _7575_/Q VGND VGND VPWR VPWR hold3088/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2354 hold935/X VGND VGND VPWR VPWR _5914_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3099 hold3099/A VGND VGND VPWR VPWR _4329_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6199_ _7483_/Q _6112_/X _6197_/X _6198_/X _6196_/X VGND VGND VPWR VPWR _6212_/B
+ sky130_fd_sc_hd__a2111o_2
Xhold1620 hold231/X VGND VGND VPWR VPWR _5888_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2365 hold947/X VGND VGND VPWR VPWR _4554_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1631 hold324/X VGND VGND VPWR VPWR _4542_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2376 _7129_/Q VGND VGND VPWR VPWR hold953/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1642 _4506_/X VGND VGND VPWR VPWR hold341/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2387 _7190_/Q VGND VGND VPWR VPWR hold919/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2398 _7100_/Q VGND VGND VPWR VPWR hold633/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1653 hold320/X VGND VGND VPWR VPWR _4331_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1664 _5918_/X VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6417__B _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1675 _4518_/X VGND VGND VPWR VPWR hold319/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1686 _7234_/Q VGND VGND VPWR VPWR hold269/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1697 hold414/X VGND VGND VPWR VPWR _5761_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6136__C _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5748__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6718__A1 _7184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6194__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3952__A1 _7391_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3792__A _3792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_31_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3704__A1 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4879__B_N _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6654__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4128__A _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4968__B1 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_168_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6709__A1 _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3640__B1 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2090_A _6926_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4196__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5570_ _4996_/A _5038_/B _5425_/X _5189_/X VGND VGND VPWR VPWR _5570_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_26_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3943__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4521_ _5866_/B _4521_/B _4551_/D VGND VGND VPWR VPWR _4526_/S sky130_fd_sc_hd__and3_2
XANTENNA__4798__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold205 hold205/A VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7240_ _7363_/CLK _7240_/D fanout575/X VGND VGND VPWR VPWR _7240_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6488__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4452_ _4452_/A0 _5914_/A1 _4454_/S VGND VGND VPWR VPWR _4452_/X sky130_fd_sc_hd__mux2_1
Xhold216 hold216/A VGND VGND VPWR VPWR _7524_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold227 hold227/A VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold238 hold238/A VGND VGND VPWR VPWR _7466_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5696__A1 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold249 hold249/A VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3403_ _3403_/A VGND VGND VPWR VPWR _3403_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4948__D _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7171_ _7213_/CLK _7171_/D fanout590/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4383_ _5714_/A0 _4383_/A1 _4387_/S VGND VGND VPWR VPWR _4383_/X sky130_fd_sc_hd__mux2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6122_/A _6122_/B VGND VGND VPWR VPWR _6122_/Y sky130_fd_sc_hd__nand2_4
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6052_/X _6051_/C _6050_/Y _6019_/Y _6462_/D VGND VGND VPWR VPWR _7596_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _4825_/A _5089_/B _4675_/A _4675_/B _4675_/C VGND VGND VPWR VPWR _5005_/C
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_178_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6956_/CLK _6955_/D fanout604/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5620__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5906_ _5987_/A1 _5906_/A1 _5910_/S VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__mux2_1
X_6886_ _4169_/B2 _6886_/D _6836_/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3631__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5837_ _5837_/A0 _5999_/A1 _5838_/S VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6176__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5768_ _5768_/A0 _5993_/A1 _5775_/S VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout605_A fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7507_ _7521_/CLK _7507_/D fanout600/X VGND VGND VPWR VPWR _7507_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3934__A1 _4175_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4719_ _4795_/C _4909_/D _4786_/C _4740_/D VGND VGND VPWR VPWR _5387_/D sky130_fd_sc_hd__and4bb_4
X_5699_ _5699_/A0 _5951_/A1 _5703_/S VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7438_ _7582_/CLK _7438_/D fanout585/X VGND VGND VPWR VPWR _7438_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold750 _4351_/X VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7369_ _7476_/CLK _7369_/D fanout586/X VGND VGND VPWR VPWR _7369_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold761 hold761/A VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold772 _4490_/X VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold783 hold783/A VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold794 _5783_/X VGND VGND VPWR VPWR _7389_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5439__A1 _5107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6636__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2140 hold145/X VGND VGND VPWR VPWR _5979_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2151 _5853_/X VGND VGND VPWR VPWR hold142/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4111__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2162 hold410/X VGND VGND VPWR VPWR _4230_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2173 hold395/X VGND VGND VPWR VPWR _7366_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input138_A wb_dat_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2184 _5658_/X VGND VGND VPWR VPWR hold437/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2195 _7518_/Q VGND VGND VPWR VPWR hold444/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1450 hold188/X VGND VGND VPWR VPWR _7492_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1461 _5926_/X VGND VGND VPWR VPWR hold172/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1472 hold198/X VGND VGND VPWR VPWR _7289_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1483 hold180/X VGND VGND VPWR VPWR _7468_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1494 hold214/X VGND VGND VPWR VPWR _7481_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3870__B1 hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3003_A _7440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5611__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4965__A3 _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_171_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5678__A1 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4350__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6627__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3461__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6642__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6057__B _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5602__A1 _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6073__A _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6740_ _7059_/Q _6447_/C _6651_/C _6435_/X _7049_/Q VGND VGND VPWR VPWR _6740_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3952_ _7391_/Q _5785_/A _5785_/B _3951_/X VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3613__B1 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6671_ _7157_/Q _6419_/A _6670_/X _6430_/X VGND VGND VPWR VPWR _6671_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_133_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6158__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3883_ _7123_/Q _4473_/A _4551_/A _4551_/C _3882_/X VGND VGND VPWR VPWR _3883_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5622_ _3933_/Y _5948_/A1 _5622_/B1 _5640_/D VGND VGND VPWR VPWR _5622_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5553_ _5553_/A1 _5339_/C _5328_/X _5552_/X _5015_/X VGND VGND VPWR VPWR _5554_/C
+ sky130_fd_sc_hd__a311oi_1
XFILLER_0_170_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2737_A _7319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4504_ _4504_/A0 _5714_/A0 _4508_/S VGND VGND VPWR VPWR _4504_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3863__C _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5484_ hold69/A _5580_/A2 _5482_/Y _5560_/B _5464_/Y VGND VGND VPWR VPWR _7205_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7223_ _7231_/CLK _7223_/D _4128_/B VGND VGND VPWR VPWR _7223_/Q sky130_fd_sc_hd__dfstp_2
X_4435_ _4435_/A0 _5996_/A1 _4439_/S VGND VGND VPWR VPWR _4435_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5851__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout504 hold48/X VGND VGND VPWR VPWR _5992_/D sky130_fd_sc_hd__buf_12
X_7154_ _7156_/CLK _7154_/D _6833_/A VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfstp_4
Xfanout515 _7595_/Q VGND VGND VPWR VPWR _6435_/B sky130_fd_sc_hd__clkbuf_16
X_4366_ _4366_/A0 _5805_/A1 _4369_/S VGND VGND VPWR VPWR _4366_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout526 _6931_/Q VGND VGND VPWR VPWR _6051_/C sky130_fd_sc_hd__buf_12
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6618__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6105_ _7303_/Q _6121_/A _6136_/C _6071_/X _7287_/Q VGND VGND VPWR VPWR _6105_/X
+ sky130_fd_sc_hd__a32o_1
X_7085_ _7513_/CLK _7085_/D fanout600/X VGND VGND VPWR VPWR _7664_/A sky130_fd_sc_hd__dfrtp_1
X_4297_ _4302_/S _3795_/B _4296_/Y VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout388_A _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6116_/C _6136_/C _6121_/C VGND VGND VPWR VPWR _6036_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__6633__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5841__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7575_/CLK _6938_/D fanout595/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6414__C _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6869_ _6873_/A _6869_/B VGND VGND VPWR VPWR _6869_/X sky130_fd_sc_hd__and2_1
XANTENNA__6149__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5357__B1 _5102_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7095__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3907__B2 _7143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5761__S _5766_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6321__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4332__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold580 hold580/A VGND VGND VPWR VPWR hold580/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold591 _5748_/X VGND VGND VPWR VPWR _7358_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6609__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5832__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3989__A4 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1280 hold3136/X VGND VGND VPWR VPWR hold3137/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1291 hold3047/X VGND VGND VPWR VPWR _7263_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_184_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3610__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6560__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6312__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2053_A _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4220_ _4220_/A0 _4219_/X _4232_/S VGND VGND VPWR VPWR _4220_/X sky130_fd_sc_hd__mux2_1
Xhold2909 _7399_/Q VGND VGND VPWR VPWR hold2909/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3677__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4151_ _6933_/Q _4168_/D _6899_/Q VGND VGND VPWR VPWR _4151_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4287__S _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6076__A1 _7511_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4082_ _6894_/Q _4082_/A2 _7073_/Q _4123_/B VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_37_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5823__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_csclk_A clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6379__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4984_ _4984_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _5339_/C sky130_fd_sc_hd__and3_4
XFILLER_0_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6723_ _7144_/Q _6468_/X _6719_/X _6720_/X _6722_/X VGND VGND VPWR VPWR _6723_/X
+ sky130_fd_sc_hd__a2111o_1
X_3935_ input52/X _5785_/B _4491_/B hold72/A _7559_/Q VGND VGND VPWR VPWR _3935_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2854_A _6947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6654_ _7051_/Q _6434_/X _6466_/X _7209_/Q _6653_/X VGND VGND VPWR VPWR _6654_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3866_ input53/X _5785_/B _5992_/C _4422_/S input44/X VGND VGND VPWR VPWR _3866_/X
+ sky130_fd_sc_hd__a32o_4
XANTENNA__6000__A1 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5605_ _5605_/A0 _5805_/A1 _5611_/S VGND VGND VPWR VPWR _5605_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_160_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6585_ _7316_/Q _6419_/D _6424_/X _7572_/Q _6584_/X VGND VGND VPWR VPWR _6585_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5354__A3 _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3797_ _3797_/A1 _3996_/A _3795_/Y _3796_/X VGND VGND VPWR VPWR _3797_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6551__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5536_ _5158_/A _5295_/C _5297_/B _5410_/A VGND VGND VPWR VPWR _5536_/Y sky130_fd_sc_hd__o211ai_1
X_5467_ _5467_/A _5467_/B _5467_/C VGND VGND VPWR VPWR _5521_/B sky130_fd_sc_hd__and3_1
XFILLER_0_78_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5106__A3 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4314__A1 _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7206_ _7206_/CLK _7206_/D _6780_/B VGND VGND VPWR VPWR _7206_/Q sky130_fd_sc_hd__dfrtp_1
X_4418_ _4446_/A0 _5998_/A1 _4422_/S VGND VGND VPWR VPWR _4418_/X sky130_fd_sc_hd__mux2_1
X_5398_ _4709_/Y _4748_/Y _5528_/A3 _4832_/Y _4826_/Y VGND VGND VPWR VPWR _5482_/A
+ sky130_fd_sc_hd__a311o_1
XANTENNA__4197__S _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7137_ _7447_/CLK _7137_/D fanout601/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_4
X_4349_ _4349_/A0 _5950_/A1 _4351_/S VGND VGND VPWR VPWR _4349_/X sky130_fd_sc_hd__mux2_1
Xfanout356 hold1491/X VGND VGND VPWR VPWR _5938_/C sky130_fd_sc_hd__buf_12
XANTENNA__6409__C _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout367 _6872_/B VGND VGND VPWR VPWR _6873_/B sky130_fd_sc_hd__buf_4
Xfanout378 _3669_/C VGND VGND VPWR VPWR _4346_/C sky130_fd_sc_hd__clkbuf_16
X_7068_ _7268_/CLK _7068_/D _6873_/A VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfstp_2
Xfanout389 _3472_/X VGND VGND VPWR VPWR _3933_/A sky130_fd_sc_hd__buf_12
XANTENNA__5814__A1 _5967_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6019_ _6051_/C _6929_/Q VGND VGND VPWR VPWR _6019_/Y sky130_fd_sc_hd__nor2_8
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4871__A_N _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__B _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4871__D _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6144__C _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7205__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4101__A_N _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4250__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5983__C hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6542__A2 _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input66_A mgmt_gpio_in[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4305__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4608__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5805__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6230__B2 _7452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _3470_/X _3485_/X _4491_/C _3669_/X _6971_/Q VGND VGND VPWR VPWR _3720_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3595__A2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3651_ _4449_/B _5938_/C _4388_/B VGND VGND VPWR VPWR _3651_/X sky130_fd_sc_hd__and3_2
XFILLER_0_130_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_0__f_wb_clk_i clkbuf_3_0_0_wb_clk_i/X VGND VGND VPWR VPWR _7601_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6533__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2170_A _7366_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4544__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2268_A _7539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6370_ _6367_/X _6368_/X _6369_/X _6144_/C VGND VGND VPWR VPWR _6370_/X sky130_fd_sc_hd__o31a_1
X_3582_ _7381_/Q _3498_/X _3564_/X _7365_/Q _3581_/X VGND VGND VPWR VPWR _3587_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3898__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5321_ _4595_/Y _4601_/Y _4622_/Y _4846_/Y _4956_/B VGND VGND VPWR VPWR _5321_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6297__B2 _7132_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5252_ _5252_/A _5252_/B _5252_/C VGND VGND VPWR VPWR _5252_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_139_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4203_ _5640_/B _5619_/A _5612_/C _5640_/D VGND VGND VPWR VPWR _4211_/S sky130_fd_sc_hd__and4_4
Xhold2706 hold757/X VGND VGND VPWR VPWR _5835_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2717 _7335_/Q VGND VGND VPWR VPWR hold2717/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3860__D _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5183_ _5183_/A _5203_/B _5183_/C _5339_/D VGND VGND VPWR VPWR _5183_/Y sky130_fd_sc_hd__nand4_1
Xhold2728 _7186_/Q VGND VGND VPWR VPWR hold837/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2739 _7070_/Q VGND VGND VPWR VPWR hold835/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4134_ _6897_/Q _4134_/B VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__and2b_4
XFILLER_0_155_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4065_ _4062_/B _4098_/A1 _6891_/Q _4062_/Y VGND VGND VPWR VPWR _4065_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3807__B1 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3822__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6221__A1 _7324_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4967_ _4966_/X _4965_/X _4964_/Y _4854_/X VGND VGND VPWR VPWR _4967_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_0_58_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6772__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3586__A2 _3506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6706_ _7013_/Q _6423_/X _6462_/X _7033_/Q _6705_/X VGND VGND VPWR VPWR _6706_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3918_ input96/X _3933_/A _5659_/B _3916_/X _3917_/X VGND VGND VPWR VPWR _3918_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout420_A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5980__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4898_ _5005_/A _4948_/B _4898_/C _5222_/B VGND VGND VPWR VPWR _4898_/Y sky130_fd_sc_hd__nand4_4
XANTENNA_fanout518_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6637_ _7302_/Q _6420_/A _6632_/X _6634_/X _6636_/X VGND VGND VPWR VPWR _6647_/A
+ sky130_fd_sc_hd__a2111o_1
X_3849_ input45/X _4422_/S _3846_/X _3847_/X _3848_/X VGND VGND VPWR VPWR _3849_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6524__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6568_ _7547_/Q _6419_/A _6435_/X _7515_/Q _6567_/X VGND VGND VPWR VPWR _6569_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4212__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3889__A3 _3519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5519_ _4717_/Y _4722_/Y _5083_/X _4718_/Y VGND VGND VPWR VPWR _5521_/D sky130_fd_sc_hd__o211a_1
X_6499_ _7489_/Q _6463_/A _6441_/X _6425_/X _7337_/Q VGND VGND VPWR VPWR _6499_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6288__A1 _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6288__B2 _6967_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1702_A _7529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3510__A2 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5799__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7457__RESET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input120_A wb_adr_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4471__A0 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3498__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6763__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold3285_A _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6515__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4526__A1 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6279__A1 _7350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5254__A2 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5870_ _5870_/A0 _5996_/A1 _5874_/S VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6203__A1 _7331_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5006__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_csclk_A _7267_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4821_ _5058_/D _4856_/A _5072_/B VGND VGND VPWR VPWR _4821_/Y sky130_fd_sc_hd__nand3_4
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6754__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7540_ _7542_/CLK _7540_/D fanout581/X VGND VGND VPWR VPWR _7540_/Q sky130_fd_sc_hd__dfrtp_2
X_4752_ _4706_/Y _4741_/Y _4751_/Y _4687_/Y _4746_/Y VGND VGND VPWR VPWR _4760_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_173_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3703_ _7387_/Q _5776_/A _3658_/X _7116_/Q VGND VGND VPWR VPWR _3703_/X sky130_fd_sc_hd__a22o_1
X_7471_ _7471_/CLK _7471_/D fanout597/X VGND VGND VPWR VPWR _7471_/Q sky130_fd_sc_hd__dfstp_2
X_4683_ _4562_/Y _4585_/Y _4687_/C VGND VGND VPWR VPWR _5138_/A sky130_fd_sc_hd__o21a_4
XANTENNA__6506__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5714__A0 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4517__A1 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6422_ _6467_/A _6747_/C _6459_/B VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__and3_4
X_3634_ _7500_/Q _5902_/A _3526_/X _7508_/Q _3633_/X VGND VGND VPWR VPWR _3642_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6353_ _6959_/Q _6036_/Y _6341_/X _6352_/X _6775_/B1 VGND VGND VPWR VPWR _6353_/X
+ sky130_fd_sc_hd__o221a_1
X_3565_ hold22/A _5875_/A _5640_/B VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__and3_4
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5304_ _4667_/A _4692_/Y _4712_/Y _4716_/Y _4755_/Y VGND VGND VPWR VPWR _5304_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3740__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6284_ _6283_/X _6284_/A1 _6777_/S VGND VGND VPWR VPWR _7609_/D sky130_fd_sc_hd__mux2_1
Xhold3204 _7626_/Q VGND VGND VPWR VPWR _6776_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3215 _7612_/Q VGND VGND VPWR VPWR _6355_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3496_ _3496_/A hold54/X VGND VGND VPWR VPWR _3496_/Y sky130_fd_sc_hd__nor2_8
Xhold3226 _7622_/Q VGND VGND VPWR VPWR _6675_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3237 _4120_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5235_ _5235_/A _5444_/D _5235_/C VGND VGND VPWR VPWR _5237_/B sky130_fd_sc_hd__and3_1
Xhold3248 _6882_/Q VGND VGND VPWR VPWR _3400_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2503 hold959/X VGND VGND VPWR VPWR _4195_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2514 hold672/X VGND VGND VPWR VPWR _5805_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3259 _7628_/Q VGND VGND VPWR VPWR _6779_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2525 _7421_/Q VGND VGND VPWR VPWR hold809/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2536 hold801/X VGND VGND VPWR VPWR _5900_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2547 _5657_/X VGND VGND VPWR VPWR hold756/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1802 _7338_/Q VGND VGND VPWR VPWR hold368/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1813 _4386_/X VGND VGND VPWR VPWR hold373/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6690__B2 _7143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5166_ _5205_/A1 _4849_/B _5295_/C _5060_/A VGND VGND VPWR VPWR _5496_/B sky130_fd_sc_hd__a31oi_4
Xhold2558 hold789/X VGND VGND VPWR VPWR _5864_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2569 hold831/X VGND VGND VPWR VPWR _5954_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1824 hold380/X VGND VGND VPWR VPWR _5951_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1835 _7274_/Q VGND VGND VPWR VPWR hold286/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4117_ _6751_/S _4117_/B VGND VGND VPWR VPWR _4117_/Y sky130_fd_sc_hd__nand2_2
Xhold1846 hold322/X VGND VGND VPWR VPWR _5869_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1857 hold342/X VGND VGND VPWR VPWR _5807_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5097_ _5097_/A _5097_/B _5444_/B VGND VGND VPWR VPWR _5097_/Y sky130_fd_sc_hd__nand3_1
Xhold1868 _7453_/Q VGND VGND VPWR VPWR hold120/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout468_A hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1879 _5824_/X VGND VGND VPWR VPWR hold499/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6442__B2 _7287_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4048_ _4062_/A _3998_/Y _3403_/Y _4113_/B1 _4048_/B1 VGND VGND VPWR VPWR _6898_/D
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5650__C1 hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5999_ _5999_/A0 _5999_/A1 hold37/X VGND VGND VPWR VPWR _5999_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6745__A2 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3559__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6422__C _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold213_A _7481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7669_ _7669_/A VGND VGND VPWR VPWR _7669_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5705__A0 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4508__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5038__C _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5181__A1 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3731__A2 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input168_A wb_sel_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6130__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput290 _6924_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XANTENNA__4893__B _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input29_A mask_rev_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3798__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6197__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6736__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6332__C _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6051__D _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3970__A2 _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_csclk _7496_/CLK VGND VGND VPWR VPWR _7476_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold409 hold409/A VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5172__B2 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7144_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7379__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5024_/A1 _4669_/X _4974_/B _5295_/C _5180_/A VGND VGND VPWR VPWR _5021_/D
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__5475__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 hold2947/X VGND VGND VPWR VPWR hold2948/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_45_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6971_ _7196_/CLK _6971_/D fanout588/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5922_ _5985_/A1 _5922_/A1 _5928_/S VGND VGND VPWR VPWR _5922_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3789__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7197_/CLK sky130_fd_sc_hd__clkbuf_16
X_5853_ _5979_/A0 _5853_/A1 _5856_/S VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6188__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5935__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4804_ _4700_/Y _4798_/Y _4803_/Y _4800_/Y VGND VGND VPWR VPWR _4809_/C sky130_fd_sc_hd__o211ai_1
XFILLER_0_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5784_ _5991_/A1 _5784_/A1 hold49/X VGND VGND VPWR VPWR _5784_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_152_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4735_ _5404_/B _5404_/C VGND VGND VPWR VPWR _4735_/Y sky130_fd_sc_hd__nand2_1
X_7523_ _7563_/CLK _7523_/D fanout599/X VGND VGND VPWR VPWR _7523_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5854__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7454_ _7572_/CLK _7454_/D fanout596/X VGND VGND VPWR VPWR _7454_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4666_ _4740_/D _4795_/C VGND VGND VPWR VPWR _4667_/C sky130_fd_sc_hd__nand2b_4
XANTENNA__4978__B _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6405_ _6462_/D _7595_/Q _6574_/B _6651_/B VGND VGND VPWR VPWR _6408_/B sky130_fd_sc_hd__and4_4
X_3617_ _4491_/A _3931_/D _5659_/B VGND VGND VPWR VPWR _3617_/X sky130_fd_sc_hd__and3_4
Xhold910 _5809_/X VGND VGND VPWR VPWR _7412_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7385_ _7577_/CLK _7385_/D fanout583/X VGND VGND VPWR VPWR _7385_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6360__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold921 hold921/A VGND VGND VPWR VPWR hold921/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4597_ _4743_/A _4856_/A VGND VGND VPWR VPWR _4843_/A sky130_fd_sc_hd__nand2b_4
XANTENNA__4697__C _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold932 _4332_/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold943 hold943/A VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3713__A2 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6336_ _6969_/Q _6136_/B _6136_/C _6332_/C _7033_/Q VGND VGND VPWR VPWR _6336_/X
+ sky130_fd_sc_hd__a32o_1
Xhold954 _4470_/X VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3548_ _4551_/A _3576_/B _3576_/C VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__and3_2
Xhold3001 _7664_/A VGND VGND VPWR VPWR hold3001/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold965 hold965/A VGND VGND VPWR VPWR hold965/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold976 _4464_/X VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3012 _7161_/Q VGND VGND VPWR VPWR hold779/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold987 hold987/A VGND VGND VPWR VPWR hold987/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3023 _7025_/Q VGND VGND VPWR VPWR hold749/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold998 _5701_/X VGND VGND VPWR VPWR _7316_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3034 hold3034/A VGND VGND VPWR VPWR _5714_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4994__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6267_ _7454_/Q _6144_/A _6116_/A _6379_/B1 _7526_/Q VGND VGND VPWR VPWR _6267_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2300 _5710_/X VGND VGND VPWR VPWR hold902/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3045 _7263_/Q VGND VGND VPWR VPWR hold3045/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout585_A fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3479_ _7398_/Q _5785_/A _3933_/A _5848_/A _7454_/Q VGND VGND VPWR VPWR _3479_/X
+ sky130_fd_sc_hd__a32o_4
Xhold2311 _7084_/Q VGND VGND VPWR VPWR hold2311/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3056 hold771/X VGND VGND VPWR VPWR _4490_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5466__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2322 hold576/X VGND VGND VPWR VPWR _5706_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3067 _6934_/Q VGND VGND VPWR VPWR hold3067/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5218_ _5079_/X _5216_/X _5213_/B VGND VGND VPWR VPWR _5218_/Y sky130_fd_sc_hd__o21ai_1
Xhold2333 _7307_/Q VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3078 _7383_/Q VGND VGND VPWR VPWR hold3078/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2344 _7300_/Q VGND VGND VPWR VPWR hold899/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6198_ _6144_/C _6089_/X _7379_/Q _6119_/X _7403_/Q VGND VGND VPWR VPWR _6198_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3089 hold3089/A VGND VGND VPWR VPWR _5993_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2355 _7364_/Q VGND VGND VPWR VPWR hold897/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1610 hold39/X VGND VGND VPWR VPWR _5775_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2366 _4554_/X VGND VGND VPWR VPWR hold948/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1621 _7330_/Q VGND VGND VPWR VPWR hold243/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1632 _4542_/X VGND VGND VPWR VPWR hold325/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2377 hold953/X VGND VGND VPWR VPWR _4470_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5149_ _4687_/Y _4777_/X _4821_/Y _4698_/Y _4723_/Y VGND VGND VPWR VPWR _5150_/C
+ sky130_fd_sc_hd__o32a_1
Xhold1643 _7362_/Q VGND VGND VPWR VPWR hold257/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2388 hold919/X VGND VGND VPWR VPWR _4543_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2399 hold633/X VGND VGND VPWR VPWR _4448_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1654 _4331_/X VGND VGND VPWR VPWR hold321/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1665 hold77/X VGND VGND VPWR VPWR _7509_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6417__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1676 hold319/X VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1687 hold269/X VGND VGND VPWR VPWR _5602_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1698 _5761_/X VGND VGND VPWR VPWR hold415/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6179__B1 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6718__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5926__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5049__B _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5764__S _5766_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3952__A2 _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4888__B _4888_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3150_A _7187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4901__A1 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3704__A2 _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4400__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6103__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7401__RESET_B fanout586/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output302_A _3619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6709__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6185__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_183_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5393__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6590__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4520_ _4520_/A0 _5586_/A0 _4520_/S VGND VGND VPWR VPWR _4520_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3943__A2 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4451_ _4451_/A0 _5583_/A0 _4454_/S VGND VGND VPWR VPWR _4451_/X sky130_fd_sc_hd__mux2_1
Xhold206 hold206/A VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold217 hold217/A VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6342__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold228 _5890_/X VGND VGND VPWR VPWR _7484_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_151_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3402_ _7071_/Q VGND VGND VPWR VPWR _4062_/A sky130_fd_sc_hd__inv_4
Xhold239 hold239/A VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7170_ _7170_/CLK _7170_/D fanout574/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_2
X_4382_ _4551_/A _5866_/B _4388_/B _4551_/D VGND VGND VPWR VPWR _4387_/S sky130_fd_sc_hd__nand4_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _6121_/A _6136_/C _6121_/C VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__and3_4
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold37_A hold37/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _7594_/Q _7593_/Q _6435_/B _6462_/D VGND VGND VPWR VPWR _6052_/X sky130_fd_sc_hd__a31o_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _4675_/A _4675_/B _4675_/C _4591_/B VGND VGND VPWR VPWR _5005_/B sky130_fd_sc_hd__a31o_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5849__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2884_A _7464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4959__B2 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6954_ _7575_/CLK hold3/X fanout595/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5905_ _5950_/A1 _5905_/A1 _5910_/S VGND VGND VPWR VPWR _5905_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3631__A1 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6885_ _4169_/B2 _6885_/D _6835_/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3631__B2 input40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5908__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5836_ _5836_/A0 _5998_/A1 _5838_/S VGND VGND VPWR VPWR _5836_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6176__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4989__A _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5767_ _5785_/A _5911_/A _5992_/D VGND VGND VPWR VPWR _5775_/S sky130_fd_sc_hd__and3_4
XANTENNA__6581__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7506_ _7513_/CLK _7506_/D fanout602/X VGND VGND VPWR VPWR _7506_/Q sky130_fd_sc_hd__dfrtp_4
X_4718_ _4803_/A _4765_/B VGND VGND VPWR VPWR _4718_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3934__A2 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5698_ _5698_/A0 _5896_/A0 _5703_/S VGND VGND VPWR VPWR _5698_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4649_ _4591_/Y _4616_/Y _4675_/A _4675_/B VGND VGND VPWR VPWR _4726_/C sky130_fd_sc_hd__nand4bb_4
XANTENNA__6333__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7437_ _7577_/CLK _7437_/D fanout584/X VGND VGND VPWR VPWR _7437_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_141_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold740 hold740/A VGND VGND VPWR VPWR hold740/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold751 hold751/A VGND VGND VPWR VPWR hold751/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7368_ _7432_/CLK hold75/X fanout586/X VGND VGND VPWR VPWR _7368_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold762 hold762/A VGND VGND VPWR VPWR _7427_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold773 hold773/A VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold784 _5738_/X VGND VGND VPWR VPWR _7349_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6319_ _7183_/Q _6097_/X _6317_/X _6318_/X _6316_/X VGND VGND VPWR VPWR _6327_/A
+ sky130_fd_sc_hd__a2111o_1
X_7299_ _7299_/CLK _7299_/D fanout576/X VGND VGND VPWR VPWR _7299_/Q sky130_fd_sc_hd__dfrtp_4
Xhold795 hold795/A VGND VGND VPWR VPWR hold795/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5439__A2 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6636__B2 _7510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2130 _7661_/A VGND VGND VPWR VPWR hold825/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2141 _5979_/X VGND VGND VPWR VPWR hold146/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2152 _7650_/A VGND VGND VPWR VPWR hold817/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2163 _4230_/X VGND VGND VPWR VPWR hold411/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2174 _7318_/Q VGND VGND VPWR VPWR hold484/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1440 _5680_/X VGND VGND VPWR VPWR hold192/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2185 _7294_/Q VGND VGND VPWR VPWR hold392/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1451 _7305_/Q VGND VGND VPWR VPWR hold189/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2196 hold444/X VGND VGND VPWR VPWR _5928_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1462 hold172/X VGND VGND VPWR VPWR _7516_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1473 _6889_/Q VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1484 _7669_/A VGND VGND VPWR VPWR hold185/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3870__A1 _7138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3870__B2 _7560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5759__S _5766_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1495 _7534_/Q VGND VGND VPWR VPWR hold1495/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4890__C _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3622__A1 _7234_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input96_A usr1_vdd_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5375__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6572__B1 _6570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6324__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6057__C _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6260__C1 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3951_ _7152_/Q _4473_/A _5632_/B _3661_/X _7031_/Q VGND VGND VPWR VPWR _3951_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6073__B _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3613__A1 _7556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3613__B2 _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2298_A _7324_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6670_ _7142_/Q _6468_/X _6667_/X _6669_/X VGND VGND VPWR VPWR _6670_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_133_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3882_ _7352_/Q _4473_/A _4212_/A _4370_/A _7042_/Q VGND VGND VPWR VPWR _3882_/X
+ sky130_fd_sc_hd__a32o_1
X_5621_ hold36/X _5590_/A _5619_/A _5621_/B1 VGND VGND VPWR VPWR _5621_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5366__A1 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6563__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3916__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5552_ _5180_/B _5342_/B _5013_/C _5183_/A VGND VGND VPWR VPWR _5552_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4503_ hold56/X _5632_/B _4551_/D VGND VGND VPWR VPWR _4508_/S sky130_fd_sc_hd__and3_2
XANTENNA__3863__D _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6315__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5483_ _5073_/A _4605_/Y _4826_/Y _5374_/X _7107_/Q VGND VGND VPWR VPWR _5560_/B
+ sky130_fd_sc_hd__o311a_1
X_4434_ _4434_/A0 _5986_/A1 _4439_/S VGND VGND VPWR VPWR _4434_/X sky130_fd_sc_hd__mux2_1
X_7222_ _7231_/CLK _7222_/D _4128_/B VGND VGND VPWR VPWR _7222_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7153_ _7156_/CLK _7153_/D _6833_/A VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfrtp_4
X_4365_ _4365_/A0 _5714_/A0 _4369_/S VGND VGND VPWR VPWR _4365_/X sky130_fd_sc_hd__mux2_1
Xfanout505 hold47/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__buf_6
Xfanout516 _7592_/Q VGND VGND VPWR VPWR _6332_/B sky130_fd_sc_hd__clkbuf_16
Xfanout527 _6930_/Q VGND VGND VPWR VPWR _6751_/S sky130_fd_sc_hd__buf_12
X_6104_ _7327_/Q _6079_/X _6091_/X _7399_/Q _6103_/X VGND VGND VPWR VPWR _6104_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7084_ _7644_/CLK _7084_/D _4309_/B VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_4
X_4296_ _4302_/S _4296_/B VGND VGND VPWR VPWR _4296_/Y sky130_fd_sc_hd__nand2_1
X_6035_ _6119_/A _6106_/B VGND VGND VPWR VPWR _6035_/Y sky130_fd_sc_hd__nor2_8
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4719__B_N _4909_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6937_ _7551_/CLK _6937_/D fanout595/X VGND VGND VPWR VPWR _7655_/A sky130_fd_sc_hd__dfrtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_74_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6414__D _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6868_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6868_/X sky130_fd_sc_hd__and2_1
XFILLER_0_181_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5819_ _5819_/A0 _5999_/A1 _5820_/S VGND VGND VPWR VPWR _5819_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6799_ _7111_/Q _6799_/A2 _6799_/B1 _7110_/Q VGND VGND VPWR VPWR _6799_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_161_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3907__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold570 hold570/A VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold581 hold581/A VGND VGND VPWR VPWR _7430_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold592 hold592/A VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input150_A wb_dat_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5293__B1 _4428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1270 hold3152/X VGND VGND VPWR VPWR hold3153/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3843__A1 _7481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input11_A mask_rev_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3843__B2 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1281 hold3138/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1292 hold3146/X VGND VGND VPWR VPWR hold3147/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6388__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5348__A1 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4795__C _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4150_ _6934_/Q _4150_/A1 _6898_/Q VGND VGND VPWR VPWR _4150_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6783__S _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4081_ _4076_/B _4050_/S _4080_/X _4121_/A VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_128_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3501__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6379__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4983_ _5038_/A _5339_/A _5399_/C VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__and3_1
XFILLER_0_144_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6722_ _7124_/Q _6420_/C _6467_/X _7154_/Q _6721_/X VGND VGND VPWR VPWR _6722_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3934_ _4175_/A _4248_/S _3652_/X _7147_/Q VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3865_ _7223_/Q hold36/A _5722_/A _5587_/C VGND VGND VPWR VPWR _3865_/X sky130_fd_sc_hd__and4_2
X_6653_ _7046_/Q _6435_/X _6443_/X _7192_/Q _6652_/X VGND VGND VPWR VPWR _6653_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6536__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5604_ _5604_/A0 _5948_/A1 _5611_/S VGND VGND VPWR VPWR _5604_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_116_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3796_ _7216_/Q _3856_/A _7073_/Q _6893_/Q VGND VGND VPWR VPWR _3796_/X sky130_fd_sc_hd__o211a_1
X_6584_ _7593_/Q _7580_/Q _6408_/C _6583_/X VGND VGND VPWR VPWR _6584_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5535_ _5535_/A _5535_/B _5535_/C VGND VGND VPWR VPWR _5539_/B sky130_fd_sc_hd__and3_1
XFILLER_0_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5862__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5466_ _4709_/Y _4722_/Y _4720_/Y _5563_/A1 VGND VGND VPWR VPWR _5467_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_14_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4417_ _4417_/A0 _4416_/X _4423_/S VGND VGND VPWR VPWR _4417_/X sky130_fd_sc_hd__mux2_1
X_7205_ _7206_/CLK _7205_/D _6780_/B VGND VGND VPWR VPWR _7205_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4314__A2 _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5397_ _4668_/C _4827_/X _5110_/X _5396_/X VGND VGND VPWR VPWR _5397_/X sky130_fd_sc_hd__a211o_1
XANTENNA_fanout498_A _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3522__B1 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4348_ _4348_/A0 _5805_/A1 _4351_/S VGND VGND VPWR VPWR _4348_/X sky130_fd_sc_hd__mux2_1
X_7136_ _7176_/CLK _7136_/D fanout588/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_input3_A debug_out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout357 _5875_/A VGND VGND VPWR VPWR _4509_/A sky130_fd_sc_hd__buf_12
XANTENNA__6409__D _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout368 _6839_/B VGND VGND VPWR VPWR _6872_/B sky130_fd_sc_hd__clkbuf_4
X_7067_ _7178_/CLK _7067_/D fanout606/X VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout379 hold1829/X VGND VGND VPWR VPWR _3669_/C sky130_fd_sc_hd__buf_12
X_4279_ _4289_/S _3996_/B _4278_/Y VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__o21ai_1
X_6018_ _6018_/A _6018_/B _6018_/C VGND VGND VPWR VPWR _7587_/D sky130_fd_sc_hd__and3_1
XFILLER_0_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3411__A _7554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__C _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6775__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3589__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6527__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6542__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5750__A1 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5772__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3761__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4896__B _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input59_A mgmt_gpio_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5502__A1 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3513__B1 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3570__A_N _3491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3816__B2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6766__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6230__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6518__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3650_ _5866_/B _4449_/B _4551_/C VGND VGND VPWR VPWR _4533_/A sky130_fd_sc_hd__and3_4
XANTENNA__6070__C _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6533__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3581_ _7493_/Q _5947_/B hold12/A _4422_/S input50/X VGND VGND VPWR VPWR _3581_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5741__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5320_ _4956_/A _4834_/Y _5529_/A _5422_/D _5319_/X VGND VGND VPWR VPWR _5320_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6297__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5251_ _4966_/A _5342_/A _5342_/B _4847_/X VGND VGND VPWR VPWR _5252_/A sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_22_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4202_ _4202_/A0 _5955_/A1 _4202_/S VGND VGND VPWR VPWR _4202_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2428_A _7184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5182_ _5034_/C _5018_/B _5180_/X _5181_/X _5179_/Y VGND VGND VPWR VPWR _5185_/A
+ sky130_fd_sc_hd__a2111oi_1
Xhold2707 _5835_/X VGND VGND VPWR VPWR hold758/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2718 hold2718/A VGND VGND VPWR VPWR _5723_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2729 hold837/X VGND VGND VPWR VPWR _4538_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4133_ input85/X _4076_/B _6897_/Q VGND VGND VPWR VPWR _4133_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4064_ _4064_/A1 _4063_/Y _4062_/B _4064_/B1 _4062_/Y VGND VGND VPWR VPWR _6892_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4480__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6221__A2 _6116_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2964_A _7367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4966_ _4966_/A _5248_/A _5248_/C VGND VGND VPWR VPWR _4966_/X sky130_fd_sc_hd__and3_1
XFILLER_0_176_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_163_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6705_ _7028_/Q _6651_/B _6459_/C _6408_/B _7043_/Q VGND VGND VPWR VPWR _6705_/X
+ sky130_fd_sc_hd__a32o_1
X_3917_ input12/X _3490_/X _3542_/X _6920_/Q _3865_/X VGND VGND VPWR VPWR _3917_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__6509__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4897_ _4622_/Y _4956_/A _4726_/Y _4895_/Y VGND VGND VPWR VPWR _4897_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5158__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6636_ _7526_/Q _6446_/X _6466_/X _7510_/Q _6635_/X VGND VGND VPWR VPWR _6636_/X
+ sky130_fd_sc_hd__a221o_1
X_3848_ _7226_/Q hold12/A _5659_/B _5713_/A _7329_/Q VGND VGND VPWR VPWR _3848_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5732__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4997__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3779_ _7009_/Q _3659_/X _4485_/A _7145_/Q VGND VGND VPWR VPWR _3779_/X sky130_fd_sc_hd__a22o_1
X_6567_ _7499_/Q _6447_/C _6429_/X _6455_/X _7459_/Q VGND VGND VPWR VPWR _6567_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3743__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5518_ _5518_/A _5518_/B _5518_/C VGND VGND VPWR VPWR _5562_/C sky130_fd_sc_hd__and3_1
X_6498_ _6497_/X _6522_/A1 _6777_/S VGND VGND VPWR VPWR _6498_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_131_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6288__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5449_ _4667_/A _4667_/C _5065_/Y _4913_/B _5228_/D VGND VGND VPWR VPWR _5450_/C
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4299__A1 _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7119_ _7447_/CLK _7119_/D fanout601/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input113_A wb_adr_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _4169_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4223__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__B _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5971__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire533 _4856_/Y VGND VGND VPWR VPWR wire533/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5723__A1 _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6279__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_189_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4462__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6203__A2 _6022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5006__A3 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7218__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4820_ _5058_/D _4856_/A _5072_/B VGND VGND VPWR VPWR _5138_/D sky130_fd_sc_hd__and3_4
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4214__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6754__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4751_ _4604_/Y _5158_/A _4790_/B _5077_/B _4898_/C VGND VGND VPWR VPWR _4751_/Y
+ sky130_fd_sc_hd__a221oi_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5962__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3702_ _7371_/Q _5758_/A _3698_/X _3699_/X _3701_/X VGND VGND VPWR VPWR _3732_/A
+ sky130_fd_sc_hd__a2111o_2
X_4682_ _4593_/A _5071_/A _5005_/A VGND VGND VPWR VPWR _4687_/C sky130_fd_sc_hd__a21boi_4
XFILLER_0_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7470_ _7510_/CLK _7470_/D fanout603/X VGND VGND VPWR VPWR _7470_/Q sky130_fd_sc_hd__dfrtp_4
X_6421_ _6455_/B _6467_/A _6651_/B VGND VGND VPWR VPWR _6421_/X sky130_fd_sc_hd__and3_4
X_3633_ _7484_/Q hold56/A _4212_/A _3520_/X _7444_/Q VGND VGND VPWR VPWR _3633_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4610__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3564_ _3564_/A _5590_/A _3931_/D VGND VGND VPWR VPWR _3564_/X sky130_fd_sc_hd__and3_4
X_6352_ _7028_/Q _6099_/X _6343_/X _6347_/X _6351_/X VGND VGND VPWR VPWR _6352_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5303_ _5303_/A _5538_/A _5405_/D _5303_/D VGND VGND VPWR VPWR _5306_/A sky130_fd_sc_hd__and4_1
XFILLER_0_12_767 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6283_ _6649_/S _7608_/Q _6281_/X _6282_/X VGND VGND VPWR VPWR _6283_/X sky130_fd_sc_hd__a22o_1
Xhold3205 _7617_/Q VGND VGND VPWR VPWR _6523_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_3495_ _7414_/Q _4473_/A _3590_/C _3494_/X _7478_/Q VGND VGND VPWR VPWR _3495_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3216 _6355_/X VGND VGND VPWR VPWR _7612_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3227 _7623_/Q VGND VGND VPWR VPWR _6676_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3238 _7613_/Q VGND VGND VPWR VPWR _6378_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5234_ _4929_/A _5180_/A _5342_/B _5102_/B _4790_/C VGND VGND VPWR VPWR _5235_/C
+ sky130_fd_sc_hd__a32oi_1
Xhold2504 _7400_/Q VGND VGND VPWR VPWR hold724/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3249 _7221_/Q VGND VGND VPWR VPWR _3573_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2515 _7349_/Q VGND VGND VPWR VPWR hold783/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2526 hold809/X VGND VGND VPWR VPWR _5819_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6690__A2 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5493__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5165_ _4595_/Y _4748_/Y _4832_/Y _4834_/Y _4709_/Y VGND VGND VPWR VPWR _5529_/A
+ sky130_fd_sc_hd__o32a_2
Xhold2537 _7134_/Q VGND VGND VPWR VPWR hold991/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2548 _7275_/Q VGND VGND VPWR VPWR hold151/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_75_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1803 hold368/X VGND VGND VPWR VPWR _5726_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2559 _7356_/Q VGND VGND VPWR VPWR hold2559/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1814 _7433_/Q VGND VGND VPWR VPWR hold420/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1825 _6905_/Q VGND VGND VPWR VPWR _4028_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4983__C _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1836 hold286/X VGND VGND VPWR VPWR _5654_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4116_ _6751_/S _4117_/B VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__and2_4
X_5096_ _5096_/A _5248_/C VGND VGND VPWR VPWR _5097_/B sky130_fd_sc_hd__nand2_1
Xhold1847 _5869_/X VGND VGND VPWR VPWR hold323/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1858 _5807_/X VGND VGND VPWR VPWR hold343/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6905__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1869 hold120/X VGND VGND VPWR VPWR _5855_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4047_ _6899_/Q _4121_/A _4047_/S VGND VGND VPWR VPWR _4047_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6442__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4453__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5650__B1 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4205__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A0 _5998_/A1 hold37/X VGND VGND VPWR VPWR _5998_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_137_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3559__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5953__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4949_ _4949_/A _4949_/B _4949_/C VGND VGND VPWR VPWR _4949_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3964__B1 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7668_ _7668_/A VGND VGND VPWR VPWR _7668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6619_ _7397_/Q _6420_/C _6467_/X _7421_/Q _6600_/X VGND VGND VPWR VPWR _6619_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_172_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7599_ _7627_/CLK _7599_/D fanout566/X VGND VGND VPWR VPWR _7599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3716__B1 _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5181__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput280 _6920_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
XANTENNA__6130__B2 _7488_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput291 _6925_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XANTENNA__4141__B1 _4140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6681__A2 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3495__A2 _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4444__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3798__A3 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5944__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3955__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_170_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output282_A _7240_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3707__B1 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5172__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire396 _5138_/C VGND VGND VPWR VPWR _4850_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6672__A2 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6791__S _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6970_ _7196_/CLK _6970_/D fanout589/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4435__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5921_ _5993_/A1 _5921_/A1 _5928_/S VGND VGND VPWR VPWR _5921_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3789__A3 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5852_ _5852_/A0 _5852_/A1 _5856_/S VGND VGND VPWR VPWR _5852_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6188__A1 _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6188__B2 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4803_ _4803_/A _4823_/B VGND VGND VPWR VPWR _4803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5783_ _5999_/A1 _5783_/A1 hold49/X VGND VGND VPWR VPWR _5783_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7522_ _7522_/CLK _7522_/D fanout605/X VGND VGND VPWR VPWR _7522_/Q sky130_fd_sc_hd__dfrtp_4
X_4734_ _4772_/A _4801_/B VGND VGND VPWR VPWR _4734_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7453_ _7572_/CLK _7453_/D fanout596/X VGND VGND VPWR VPWR _7453_/Q sky130_fd_sc_hd__dfrtp_4
X_4665_ _4740_/D _4795_/C VGND VGND VPWR VPWR _4797_/B sky130_fd_sc_hd__and2b_4
XFILLER_0_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6404_ _7597_/Q _7598_/Q VGND VGND VPWR VPWR _6404_/Y sky130_fd_sc_hd__nor2_8
X_3616_ _7348_/Q _5947_/A _5731_/B VGND VGND VPWR VPWR _3616_/X sky130_fd_sc_hd__and3_1
Xhold900 _5683_/X VGND VGND VPWR VPWR _7300_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7384_ _7577_/CLK hold50/X fanout584/X VGND VGND VPWR VPWR _7384_/Q sky130_fd_sc_hd__dfstp_2
Xhold911 hold911/A VGND VGND VPWR VPWR hold911/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4596_ _4887_/D _4747_/B VGND VGND VPWR VPWR _4748_/C sky130_fd_sc_hd__and2b_2
Xhold922 _5692_/X VGND VGND VPWR VPWR _7308_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6360__B2 _7185_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4371__A0 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold933 hold933/A VGND VGND VPWR VPWR hold933/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold944 hold944/A VGND VGND VPWR VPWR _7441_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6335_ _7003_/Q _6116_/C _6120_/B _6317_/C _7114_/Q VGND VGND VPWR VPWR _6335_/X
+ sky130_fd_sc_hd__a32o_1
X_3547_ _6926_/Q _3542_/X _3543_/X _7294_/Q _3546_/X VGND VGND VPWR VPWR _3568_/B
+ sky130_fd_sc_hd__a221o_4
XANTENNA__3713__A3 _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold955 hold955/A VGND VGND VPWR VPWR hold955/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold966 _5782_/X VGND VGND VPWR VPWR _7388_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3002 hold3002/A VGND VGND VPWR VPWR _4432_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold977 hold977/A VGND VGND VPWR VPWR hold977/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3013 hold779/X VGND VGND VPWR VPWR _4508_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3024 hold749/X VGND VGND VPWR VPWR _4351_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold988 _4500_/X VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold999 hold999/A VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6266_ _7398_/Q _6379_/B1 _6094_/A _6265_/X _6263_/X VGND VGND VPWR VPWR _6266_/X
+ sky130_fd_sc_hd__a2111o_1
X_3478_ _4551_/A hold22/A _5866_/B VGND VGND VPWR VPWR _5848_/A sky130_fd_sc_hd__and3_4
Xhold3035 _7118_/Q VGND VGND VPWR VPWR hold3035/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_86_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3046 hold3046/A VGND VGND VPWR VPWR _5641_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2301 _7510_/Q VGND VGND VPWR VPWR hold563/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3057 _7067_/Q VGND VGND VPWR VPWR hold3057/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2312 _4429_/B VGND VGND VPWR VPWR _3468_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6663__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2323 _6969_/Q VGND VGND VPWR VPWR hold895/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3068 hold3068/A VGND VGND VPWR VPWR _4220_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5217_ _5213_/C _5342_/B _4940_/D _5079_/X VGND VGND VPWR VPWR _5217_/X sky130_fd_sc_hd__a31o_1
Xhold2334 hold88/X VGND VGND VPWR VPWR _5691_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout480_A _5735_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3079 hold3079/A VGND VGND VPWR VPWR _5777_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1600 hold263/X VGND VGND VPWR VPWR _5779_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6197_ _7411_/Q _6144_/C _6116_/C _6144_/B VGND VGND VPWR VPWR _6197_/X sky130_fd_sc_hd__o211a_1
XANTENNA_fanout578_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2345 hold899/X VGND VGND VPWR VPWR _5683_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2356 hold897/X VGND VGND VPWR VPWR _5755_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1611 _5775_/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1622 hold243/X VGND VGND VPWR VPWR _5717_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2367 _7028_/Q VGND VGND VPWR VPWR hold961/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2378 _7478_/Q VGND VGND VPWR VPWR hold606/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1633 _7548_/Q VGND VGND VPWR VPWR hold261/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5148_ _5148_/A _5308_/A _5148_/C VGND VGND VPWR VPWR _5150_/B sky130_fd_sc_hd__nor3_1
Xhold1644 hold257/X VGND VGND VPWR VPWR _5753_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2389 _7004_/Q VGND VGND VPWR VPWR hold945/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1655 hold321/X VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1666 _7442_/Q VGND VGND VPWR VPWR hold245/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_98_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1677 _7572_/Q VGND VGND VPWR VPWR hold233/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5079_ _5100_/A _5079_/B _5248_/C VGND VGND VPWR VPWR _5079_/X sky130_fd_sc_hd__and3_1
Xhold1688 _5602_/X VGND VGND VPWR VPWR hold270/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1699 _7517_/Q VGND VGND VPWR VPWR hold1699/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_79_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4515__A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6179__A1 _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6179__B2 _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6718__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5049__C _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__1111_ clkbuf_0__1111_/X VGND VGND VPWR VPWR _3734_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3952__A3 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4888__C _5282_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5065__B _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3704__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5780__S hold49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4400__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input41_A mgmt_gpio_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6654__A2 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5081__A _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5862__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2890 hold2890/A VGND VGND VPWR VPWR _5637_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4968__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3640__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5378__C1 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5917__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_183_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4450_ _4450_/A0 _5840_/A1 _4454_/S VGND VGND VPWR VPWR _4450_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold207 hold207/A VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold218 hold218/A VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold229 hold229/A VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3401_ _6890_/Q VGND VGND VPWR VPWR _3401_/Y sky130_fd_sc_hd__inv_2
X_4381_ _4381_/A0 _5586_/A0 _4381_/S VGND VGND VPWR VPWR _4381_/X sky130_fd_sc_hd__mux2_1
X_6120_ _6121_/A _6120_/B _6121_/C VGND VGND VPWR VPWR _6120_/X sky130_fd_sc_hd__and3_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6462_/D _6435_/B _6051_/C _6434_/B VGND VGND VPWR VPWR _6051_/Y sky130_fd_sc_hd__nand4_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5853__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5002_ _5024_/A1 _4669_/X _4974_/B _5038_/C _5158_/A VGND VGND VPWR VPWR _5025_/D
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_147_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4408__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4959__A2 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6953_ _7575_/CLK _6953_/D fanout595/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5904_ _5967_/A1 _5904_/A1 _5910_/S VGND VGND VPWR VPWR _5904_/X sky130_fd_sc_hd__mux2_1
X_6884_ _4169_/B2 _6884_/D _6834_/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3631__A2 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _5835_/A0 _5997_/A1 _5838_/S VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5865__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_173_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5766_ _5955_/A1 _5766_/A1 _5766_/S VGND VGND VPWR VPWR _5766_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6581__B2 _7492_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7505_ _7505_/CLK _7505_/D fanout601/X VGND VGND VPWR VPWR _7505_/Q sky130_fd_sc_hd__dfrtp_4
X_4717_ _5260_/C _4717_/B VGND VGND VPWR VPWR _4717_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5697_ _5697_/A0 _5967_/A1 _5703_/S VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7436_ _7556_/CLK _7436_/D fanout594/X VGND VGND VPWR VPWR _7436_/Q sky130_fd_sc_hd__dfrtp_4
X_4648_ _4648_/A _4825_/A VGND VGND VPWR VPWR _4726_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4344__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold730 hold730/A VGND VGND VPWR VPWR hold730/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold741 hold741/A VGND VGND VPWR VPWR _7467_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7367_ _7575_/CLK _7367_/D fanout595/X VGND VGND VPWR VPWR _7367_/Q sky130_fd_sc_hd__dfstp_4
X_4579_ _4795_/C _4740_/D _4772_/A _4805_/B VGND VGND VPWR VPWR _4643_/C sky130_fd_sc_hd__and4_4
XFILLER_0_141_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap460 _4730_/C VGND VGND VPWR VPWR _4801_/B sky130_fd_sc_hd__buf_6
Xhold752 hold752/A VGND VGND VPWR VPWR _7233_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold763 hold763/A VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold774 _4544_/X VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6318_ _7067_/Q _6110_/A _6332_/C _6092_/X _7178_/Q VGND VGND VPWR VPWR _6318_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_70_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold785 hold785/A VGND VGND VPWR VPWR hold785/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7298_ _7501_/CLK _7298_/D fanout580/X VGND VGND VPWR VPWR _7298_/Q sky130_fd_sc_hd__dfrtp_4
Xhold796 _5801_/X VGND VGND VPWR VPWR _7405_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6636__A2 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5439__A3 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6249_ _7421_/Q _6072_/X _6099_/X _7357_/Q _6248_/X VGND VGND VPWR VPWR _6257_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2120 _4441_/X VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3414__A _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2131 hold825/X VGND VGND VPWR VPWR _4419_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2142 _7395_/Q VGND VGND VPWR VPWR hold164/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2153 hold817/X VGND VGND VPWR VPWR _4241_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2164 _7654_/A VGND VGND VPWR VPWR hold868/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1430 _7273_/Q VGND VGND VPWR VPWR hold181/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2175 hold484/X VGND VGND VPWR VPWR _5703_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1441 hold192/X VGND VGND VPWR VPWR _7297_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2186 hold392/X VGND VGND VPWR VPWR _5676_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2197 _5928_/X VGND VGND VPWR VPWR hold445/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1452 hold189/X VGND VGND VPWR VPWR _5689_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_99_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1463 _7205_/Q VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1474 hold15/X VGND VGND VPWR VPWR _4201_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 hold185/X VGND VGND VPWR VPWR _4437_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7499_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3870__A2 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1496 hold1496/A VGND VGND VPWR VPWR _5946_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3622__A2 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_csclk clkbuf_3_1_0_csclk/X VGND VGND VPWR VPWR _7266_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5775__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3093_A _7487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_192_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input89_A spimemio_flash_io2_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3689__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7201_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6088__B1 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6627__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4638__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_29_csclk _7267_/CLK VGND VGND VPWR VPWR _7513_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_187_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6079__B_N _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3950_ _7359_/Q _5803_/A hold12/A _3946_/X _3949_/X VGND VGND VPWR VPWR _3961_/C
+ sky130_fd_sc_hd__a311o_1
XANTENNA__6073__C _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3613__A2 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3881_ _6875_/Q _5866_/B _5632_/B _3880_/X VGND VGND VPWR VPWR _3881_/X sky130_fd_sc_hd__a31o_1
XANTENNA_hold2193_A _7519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5620_ _5620_/A0 _5948_/A1 _5620_/S VGND VGND VPWR VPWR _5620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6563__B2 _7339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5551_ _4975_/X _5424_/X _5340_/A _5169_/X _5438_/D VGND VGND VPWR VPWR _5551_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__4602__B _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4502_ _5979_/A0 _4502_/A1 _4502_/S VGND VGND VPWR VPWR _4502_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5482_ _5482_/A _5482_/B _5560_/A VGND VGND VPWR VPWR _5482_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__4326__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7221_ _7075_/CLK _7221_/D _6873_/X VGND VGND VPWR VPWR _7221_/Q sky130_fd_sc_hd__dfrtn_1
X_4433_ _4433_/A0 _5985_/A1 _4439_/S VGND VGND VPWR VPWR _4433_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7152_ _7156_/CLK _7152_/D _6833_/A VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfrtp_4
X_4364_ _5803_/A _5623_/B _5902_/B VGND VGND VPWR VPWR _4369_/S sky130_fd_sc_hd__and3_2
XFILLER_0_6_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout506 hold1418/X VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__buf_6
Xfanout517 _7592_/Q VGND VGND VPWR VPWR _6112_/C sky130_fd_sc_hd__buf_4
X_6103_ _7335_/Q _6121_/A _6120_/B _6332_/C _7359_/Q VGND VGND VPWR VPWR _6103_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6618__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout528 _6930_/Q VGND VGND VPWR VPWR _6649_/S sky130_fd_sc_hd__buf_8
X_7083_ _7513_/CLK _7083_/D fanout600/X VGND VGND VPWR VPWR _7663_/A sky130_fd_sc_hd__dfrtp_1
X_4295_ _4302_/S _3856_/B _4294_/Y VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__4629__A1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6034_ _6119_/A _6019_/Y _6033_/X VGND VGND VPWR VPWR _7591_/D sky130_fd_sc_hd__a21o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4644__A4 _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3852__A2 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5054__A1 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6251__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5054__B2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _7551_/CLK _6936_/D fanout595/X VGND VGND VPWR VPWR _7654_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout443_A _6035_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3604__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6867_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6867_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5818_ _5818_/A0 _5953_/A1 _5820_/S VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6798_ _6797_/X _6798_/B _6798_/C VGND VGND VPWR VPWR _6822_/S sky130_fd_sc_hd__nand3b_4
XFILLER_0_134_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3907__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5749_ _5803_/A hold12/X _5902_/B VGND VGND VPWR VPWR _5757_/S sky130_fd_sc_hd__and3_4
XFILLER_0_134_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6306__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7419_ _7471_/CLK _7419_/D fanout593/X VGND VGND VPWR VPWR _7419_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4868__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold560 _5734_/X VGND VGND VPWR VPWR _7345_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold571 hold571/A VGND VGND VPWR VPWR _7326_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold582 hold582/A VGND VGND VPWR VPWR hold582/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold593 hold593/A VGND VGND VPWR VPWR _7280_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6609__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input143_A wb_dat_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6490__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6455__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1260 hold3069/X VGND VGND VPWR VPWR hold3070/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1271 hold3154/X VGND VGND VPWR VPWR _7471_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1282 hold3104/X VGND VGND VPWR VPWR hold3105/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1293 _4335_/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6242__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4703__A _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5348__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4556__A0 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4795__D _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4080_ _6908_/Q _6882_/Q _4062_/A _4001_/Y VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6076__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5284__A1 _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6481__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3834__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6084__B _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5036__A1 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6233__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3501__B _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4982_ _4996_/A _5339_/D _5339_/A _5295_/C VGND VGND VPWR VPWR _5044_/C sky130_fd_sc_hd__nand4_2
X_6721_ _7058_/Q _6600_/B _6651_/C _6452_/X _7023_/Q VGND VGND VPWR VPWR _6721_/X
+ sky130_fd_sc_hd__a32o_1
X_3933_ _3933_/A _5619_/A VGND VGND VPWR VPWR _3933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6652_ _7137_/Q _6419_/C _6446_/X _7187_/Q VGND VGND VPWR VPWR _6652_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3864_ hold36/A _5722_/A _5587_/C VGND VGND VPWR VPWR _3864_/X sky130_fd_sc_hd__and3_1
XANTENNA__6536__A1 _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6536__B2 _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4547__A0 _5583_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5603_ _5612_/B _5603_/B _5640_/D VGND VGND VPWR VPWR _5611_/S sky130_fd_sc_hd__and3_4
XFILLER_0_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6583_ _7436_/Q _6747_/B _6645_/C _6408_/A _7556_/Q VGND VGND VPWR VPWR _6583_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3795_ _3923_/S _3795_/B VGND VGND VPWR VPWR _3795_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5534_ _4811_/A _5410_/C _5410_/A _5160_/D _5317_/C VGND VGND VPWR VPWR _5535_/C
+ sky130_fd_sc_hd__a311oi_1
XFILLER_0_42_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5465_ _4601_/Y _4700_/Y _4844_/Y _5077_/Y VGND VGND VPWR VPWR _5467_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_169_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7204_ _7206_/CLK _7204_/D _6780_/B VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfrtp_1
X_4416_ _4445_/A0 _5586_/A0 _4422_/S VGND VGND VPWR VPWR _4416_/X sky130_fd_sc_hd__mux2_1
X_5396_ _4817_/X _5453_/C _5394_/Y _5395_/X VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__a211o_1
X_7135_ _7186_/CLK _7135_/D fanout588/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfrtp_4
X_4347_ _4347_/A0 _5948_/A1 _4351_/S VGND VGND VPWR VPWR _4347_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_185_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout358 _5875_/A VGND VGND VPWR VPWR _5866_/B sky130_fd_sc_hd__buf_12
XFILLER_0_185_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7066_ _7191_/CLK _7066_/D _6871_/A VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout369 _4078_/Y VGND VGND VPWR VPWR _6839_/B sky130_fd_sc_hd__buf_12
X_4278_ _4289_/S _4278_/B VGND VGND VPWR VPWR _4278_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6472__B1 _7279_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6017_ _7585_/Q _7586_/Q _7587_/Q _6017_/D VGND VGND VPWR VPWR _6018_/C sky130_fd_sc_hd__nand4_1
XANTENNA__3825__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3443__2/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__6775__A1 _6961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5578__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919_ _7255_/CLK _6919_/D fanout565/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4250__A2 hold284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6527__A1 _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6527__B2 _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4538__A0 _5586_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_190_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1842_A _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold390 hold390/A VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3513__B2 _7310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3816__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 hold2921/X VGND VGND VPWR VPWR hold2922/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_185_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6518__A1 _7393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5248__B _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3580_ _7501_/Q _5902_/A _3542_/X _6925_/Q _3579_/X VGND VGND VPWR VPWR _3587_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3752__A1 _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3752__B2 _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6297__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5250_ _4743_/A _5399_/A _4953_/X _5249_/Y VGND VGND VPWR VPWR _5252_/C sky130_fd_sc_hd__a31o_1
XANTENNA__6151__C1 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4201_ _4201_/A0 _7644_/Q _7084_/Q VGND VGND VPWR VPWR _4201_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_139_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2708 _7213_/Q VGND VGND VPWR VPWR hold819/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5181_ _5295_/C _5183_/C _5180_/A _5216_/A VGND VGND VPWR VPWR _5181_/X sky130_fd_sc_hd__o211a_1
Xhold2719 _5723_/X VGND VGND VPWR VPWR hold2719/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2323_A _6969_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4132_ _4132_/A VGND VGND VPWR VPWR _4132_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold12_A hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4063_ _3401_/Y _6892_/Q _7071_/Q VGND VGND VPWR VPWR _4063_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3512__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3807__A2 _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6206__B1 _6073_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_171_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6221__A3 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4965_ _4966_/A _5342_/A _5138_/D _4847_/X VGND VGND VPWR VPWR _4965_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_80_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2957_A _7511_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6704_ _7114_/Q _6651_/B _6426_/X _6703_/X VGND VGND VPWR VPWR _6704_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_74_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3916_ _7368_/Q _5758_/A _5776_/A _7384_/Q _3860_/X VGND VGND VPWR VPWR _3916_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6509__B2 _7569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4896_ _4966_/A _5158_/A _5222_/B _5222_/C VGND VGND VPWR VPWR _4896_/Y sky130_fd_sc_hd__nand4_4
X_6635_ _7342_/Q _6425_/X _6460_/X _7390_/Q VGND VGND VPWR VPWR _6635_/X sky130_fd_sc_hd__a22o_1
X_3847_ _7246_/Q _5947_/A _3519_/B _3598_/X VGND VGND VPWR VPWR _3847_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3991__B2 _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6566_ _7555_/Q _6408_/A _6408_/D _7539_/Q _6565_/X VGND VGND VPWR VPWR _6569_/C
+ sky130_fd_sc_hd__a221o_1
X_3778_ _7059_/Q hold56/A _4521_/B _3739_/X VGND VGND VPWR VPWR _3782_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3743__A1 _7562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5517_ _5563_/A1 _4796_/Y _5471_/X _5516_/X VGND VGND VPWR VPWR _5518_/B sky130_fd_sc_hd__o31a_1
XANTENNA__3743__B2 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6497_ _6649_/S _7615_/Q _6495_/Y _6496_/X VGND VGND VPWR VPWR _6497_/X sky130_fd_sc_hd__a22o_1
X_5448_ _5445_/X _5448_/B _5508_/A _5448_/D VGND VGND VPWR VPWR _5452_/B sky130_fd_sc_hd__and4b_1
XANTENNA__6693__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5379_ _4703_/Y _4844_/Y _4737_/Y _5563_/A1 VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5902__A _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7118_ _7197_/CLK _7118_/D fanout601/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6445__B1 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7049_ _7176_/CLK _7049_/D fanout588/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3422__A _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_179_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6748__A1 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A wb_adr_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6452__B _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_182_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3982__A1 _7244_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3982__B2 _7487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5783__S hold49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input71_A mgmt_gpio_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4700__B _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6684__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5812__A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5239__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6436__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4998__B1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6739__A1 _7145_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6203__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4750_ _5260_/A _5260_/B _5094_/A VGND VGND VPWR VPWR _4898_/C sky130_fd_sc_hd__and3_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6081__C _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3701_ _7475_/Q _3494_/X _3529_/X _7531_/Q _3700_/X VGND VGND VPWR VPWR _3701_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4681_ _5158_/A _4952_/B VGND VGND VPWR VPWR _4681_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6420_ _6420_/A _6420_/B _6420_/C _6419_/Y VGND VGND VPWR VPWR _6431_/C sky130_fd_sc_hd__nor4b_4
XFILLER_0_71_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3632_ _3632_/A _3632_/B _3632_/C _3632_/D VGND VGND VPWR VPWR _3643_/B sky130_fd_sc_hd__nor4_2
XFILLER_0_114_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3725__A1 _7259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6351_ _7164_/Q _6075_/X _6350_/X _6332_/X _6349_/X VGND VGND VPWR VPWR _6351_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4610__B _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3563_ _7302_/Q hold12/A _3669_/C VGND VGND VPWR VPWR _3563_/X sky130_fd_sc_hd__and3_1
XFILLER_0_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5302_ _4741_/Y _4755_/Y _4687_/Y _5135_/Y _5297_/Y VGND VGND VPWR VPWR _5303_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6282_ _7286_/Q _6036_/Y _6775_/B1 VGND VGND VPWR VPWR _6282_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_12_779 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3494_ _5590_/A _5875_/A _5938_/B VGND VGND VPWR VPWR _3494_/X sky130_fd_sc_hd__and3_4
Xhold3206 _7644_/Q VGND VGND VPWR VPWR _6822_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3217 _7611_/Q VGND VGND VPWR VPWR _6331_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5233_ _4954_/C _4929_/A _4943_/B _5102_/B _4790_/C VGND VGND VPWR VPWR _5233_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3228 _7604_/Q VGND VGND VPWR VPWR _6170_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3239 _7620_/Q VGND VGND VPWR VPWR _6599_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2505 hold724/X VGND VGND VPWR VPWR _5796_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5722__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2516 hold783/X VGND VGND VPWR VPWR _5738_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4150__A1 _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2527 _5819_/X VGND VGND VPWR VPWR hold810/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5164_ _5164_/A _5164_/B VGND VGND VPWR VPWR _5167_/A sky130_fd_sc_hd__nor2_1
Xhold2538 hold991/X VGND VGND VPWR VPWR _4476_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1804 _5726_/X VGND VGND VPWR VPWR hold369/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2549 hold151/X VGND VGND VPWR VPWR _5655_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1815 hold420/X VGND VGND VPWR VPWR _5833_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4115_ _6827_/A _4115_/B VGND VGND VPWR VPWR _4115_/Y sky130_fd_sc_hd__nand2b_1
Xhold1826 _3448_/X VGND VGND VPWR VPWR _3449_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1837 _5654_/X VGND VGND VPWR VPWR hold287/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5095_ _4887_/B _5091_/A _5096_/A _5093_/Y VGND VGND VPWR VPWR _5097_/A sky130_fd_sc_hd__a31oi_1
Xhold1848 _7038_/Q VGND VGND VPWR VPWR hold506/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1859 hold343/X VGND VGND VPWR VPWR _7410_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4046_ _6910_/Q _6909_/Q _6908_/Q _7071_/Q VGND VGND VPWR VPWR _4047_/S sky130_fd_sc_hd__and4_1
XANTENNA__6442__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5650__A1 _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _5997_/A0 _5997_/A1 hold37/X VGND VGND VPWR VPWR _5997_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4948_ _4966_/A _4948_/B _4948_/C _5248_/C VGND VGND VPWR VPWR _4949_/B sky130_fd_sc_hd__and4_1
XFILLER_0_148_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7667_ _7667_/A VGND VGND VPWR VPWR _7667_/X sky130_fd_sc_hd__clkbuf_2
X_4879_ _4747_/B _4887_/B _4879_/C _4887_/D VGND VGND VPWR VPWR _5342_/B sky130_fd_sc_hd__and4bb_4
XFILLER_0_163_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6618_ _7549_/Q _6419_/A _6455_/X _7461_/Q _6602_/X VGND VGND VPWR VPWR _6618_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_160_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7598_ _7610_/CLK _7598_/D fanout568/X VGND VGND VPWR VPWR _7598_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_132_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3716__B2 _7499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6549_ _7571_/Q _6424_/X _6427_/X _7579_/Q VGND VGND VPWR VPWR _6549_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3417__A _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput270 _6913_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
XANTENNA__6130__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput281 _7239_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
Xoutput292 _6926_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XANTENNA__4141__A1 _7578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6447__B _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3495__A3 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5641__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5778__S hold49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_186_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6463__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6197__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5079__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3955__A1 _7527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire364 _4594_/Y VGND VGND VPWR VPWR _4836_/A sky130_fd_sc_hd__buf_2
XANTENNA_output275_A _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4380__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6657__B1 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5880__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5920_ _5920_/A _5992_/D VGND VGND VPWR VPWR _5928_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5851_ _5986_/A1 _5851_/A1 _5856_/S VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6092__B _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6188__A2 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4802_ _4802_/A _5404_/C VGND VGND VPWR VPWR _4802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5782_ _5953_/A1 _5782_/A1 hold49/X VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7521_ _7521_/CLK _7521_/D fanout600/X VGND VGND VPWR VPWR _7521_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4733_ _4733_/A _4733_/B _4984_/B VGND VGND VPWR VPWR _5404_/C sky130_fd_sc_hd__and3_4
XFILLER_0_29_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7452_ _7572_/CLK _7452_/D fanout596/X VGND VGND VPWR VPWR _7452_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4664_ _4568_/Y _4984_/C _4861_/B VGND VGND VPWR VPWR _4974_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5699__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6403_ _6463_/A _6427_/A _6747_/C VGND VGND VPWR VPWR _6408_/A sky130_fd_sc_hd__and3_4
XFILLER_0_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3615_ _7292_/Q _3543_/X _4422_/S input49/X _3614_/X VGND VGND VPWR VPWR _3623_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4340__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7383_ _7575_/CLK _7383_/D fanout595/X VGND VGND VPWR VPWR _7383_/Q sky130_fd_sc_hd__dfstp_4
Xhold901 hold901/A VGND VGND VPWR VPWR hold901/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6360__A2 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4595_ _5295_/A _5295_/D VGND VGND VPWR VPWR _4595_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_40_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold912 hold912/A VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold923 hold923/A VGND VGND VPWR VPWR hold923/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6334_ _7144_/Q _6121_/C _6116_/C _6136_/C VGND VGND VPWR VPWR _6334_/X sky130_fd_sc_hd__o211a_1
Xhold934 _5788_/X VGND VGND VPWR VPWR _7393_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3546_ _7422_/Q _4509_/A _4212_/A _3545_/X _7350_/Q VGND VGND VPWR VPWR _3546_/X
+ sky130_fd_sc_hd__a32o_1
Xhold945 hold945/A VGND VGND VPWR VPWR hold945/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold956 hold956/A VGND VGND VPWR VPWR _7227_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold967 hold967/A VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3003 _7440_/Q VGND VGND VPWR VPWR hold3003/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold978 _5764_/X VGND VGND VPWR VPWR _7372_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3014 _7657_/A VGND VGND VPWR VPWR hold3014/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6265_ _7390_/Q _6073_/X _6079_/X _7334_/Q _6264_/X VGND VGND VPWR VPWR _6265_/X
+ sky130_fd_sc_hd__a221o_1
Xhold989 hold989/A VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3025 _7233_/Q VGND VGND VPWR VPWR hold751/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3477_ _3557_/C hold54/X VGND VGND VPWR VPWR _3477_/Y sky130_fd_sc_hd__nor2_1
Xhold3036 hold3036/A VGND VGND VPWR VPWR _4457_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4994__C _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3047 _5641_/X VGND VGND VPWR VPWR hold3047/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2302 hold563/X VGND VGND VPWR VPWR _5919_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_86_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5216_ _5216_/A _5342_/B _5339_/C VGND VGND VPWR VPWR _5216_/X sky130_fd_sc_hd__and3_2
Xhold3058 hold3058/A VGND VGND VPWR VPWR _4402_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2313 _3468_/X VGND VGND VPWR VPWR _3474_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3069 _7066_/Q VGND VGND VPWR VPWR hold3069/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6196_ _7443_/Q _6097_/X _6121_/X _7307_/Q _6195_/X VGND VGND VPWR VPWR _6196_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6663__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2324 hold895/X VGND VGND VPWR VPWR _4274_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2335 _7064_/Q VGND VGND VPWR VPWR hold913/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5871__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1601 _5779_/X VGND VGND VPWR VPWR hold264/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2346 _7180_/Q VGND VGND VPWR VPWR hold925/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2357 _7037_/Q VGND VGND VPWR VPWR hold629/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1612 hold40/X VGND VGND VPWR VPWR _7382_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1623 _5717_/X VGND VGND VPWR VPWR hold244/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5147_ _4778_/A _4758_/X _5410_/B _5086_/B _4706_/A VGND VGND VPWR VPWR _5148_/C
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout473_A _4256_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2368 hold961/X VGND VGND VPWR VPWR _4355_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2379 hold606/X VGND VGND VPWR VPWR _5883_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1634 hold261/X VGND VGND VPWR VPWR _5962_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1645 _5753_/X VGND VGND VPWR VPWR hold258/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1656 _7386_/Q VGND VGND VPWR VPWR hold290/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1667 hold245/X VGND VGND VPWR VPWR _5843_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5078_ _4571_/Y _4843_/A _4727_/Y _4946_/Y _5077_/Y VGND VGND VPWR VPWR _5467_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_169_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1678 hold233/X VGND VGND VPWR VPWR _5989_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1689 _7091_/Q VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4029_ _6902_/Q _6901_/Q _6900_/Q _4025_/A VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_79_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4515__B _4551_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6179__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1490_A _3496_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3937__A1 _7311_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1755_A _7469_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6351__A2 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5154__A3 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4362__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6639__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6103__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3456__A_N _4429_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input34_A mask_rev_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2880 _7495_/Q VGND VGND VPWR VPWR hold2880/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2891 _5637_/X VGND VGND VPWR VPWR hold2891/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3625__B1 _5929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3640__A3 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_183_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6590__A2 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6342__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5971__S hold13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold208 hold208/A VGND VGND VPWR VPWR _7580_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold219 hold219/A VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3400_ _3400_/A VGND VGND VPWR VPWR _3400_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4353__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4380_ _4380_/A0 _5852_/A0 _4381_/S VGND VGND VPWR VPWR _4380_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2236_A _7406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _7594_/Q _7593_/Q _6462_/D _6435_/B VGND VGND VPWR VPWR _6050_/Y sky130_fd_sc_hd__nand4_4
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6087__B _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5024_/A1 _4669_/X _4974_/B _5295_/C _5038_/C VGND VGND VPWR VPWR _5025_/C
+ sky130_fd_sc_hd__o2111ai_4
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2403_A _6965_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5605__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7569__RESET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6307__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6952_ _7551_/CLK _6952_/D fanout595/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3520__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4959__A3 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5903_ _5903_/A0 _5903_/A1 _5910_/S VGND VGND VPWR VPWR _5903_/X sky130_fd_sc_hd__mux2_1
X_6883_ _4169_/B2 _6883_/D _6833_/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2772_A _7132_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ _5834_/A0 _5987_/A1 _5838_/S VGND VGND VPWR VPWR _5834_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6030__A1 _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7151__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5765_ _5954_/A1 _5765_/A1 _5766_/S VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6581__A2 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4989__C _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7504_ _7521_/CLK _7504_/D fanout600/X VGND VGND VPWR VPWR _7504_/Q sky130_fd_sc_hd__dfstp_4
X_4716_ _5260_/A _5079_/B VGND VGND VPWR VPWR _4716_/Y sky130_fd_sc_hd__nand2_4
X_5696_ _5696_/A0 _5903_/A0 _5703_/S VGND VGND VPWR VPWR _7311_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7435_ _7569_/CLK _7435_/D fanout593/X VGND VGND VPWR VPWR _7435_/Q sky130_fd_sc_hd__dfrtp_4
X_4647_ _4646_/A _4646_/B _4643_/Y _5071_/A VGND VGND VPWR VPWR _4647_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6333__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5881__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7366_ _7366_/CLK _7366_/D fanout579/X VGND VGND VPWR VPWR _7366_/Q sky130_fd_sc_hd__dfrtp_4
Xhold720 hold720/A VGND VGND VPWR VPWR hold720/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4578_ _4984_/C _4578_/B VGND VGND VPWR VPWR _4675_/C sky130_fd_sc_hd__nor2_8
Xhold731 _4196_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold742 hold742/A VGND VGND VPWR VPWR hold742/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap450 _5118_/B VGND VGND VPWR VPWR _5399_/D sky130_fd_sc_hd__clkbuf_2
Xmax_cap461 wire462/X VGND VGND VPWR VPWR _5580_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold753 hold753/A VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6317_ _7047_/Q _7592_/Q _6317_/C VGND VGND VPWR VPWR _6317_/X sky130_fd_sc_hd__and3_1
Xhold764 hold764/A VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout590_A fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3529_ hold22/A _5938_/B _5938_/C VGND VGND VPWR VPWR _3529_/X sky130_fd_sc_hd__and3_4
Xhold775 hold775/A VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7297_ _7539_/CLK _7297_/D fanout577/X VGND VGND VPWR VPWR _7297_/Q sky130_fd_sc_hd__dfrtp_4
Xhold786 _4333_/X VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold797 hold797/A VGND VGND VPWR VPWR hold797/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6248_ _7429_/Q _6112_/C _6074_/X _6120_/X _7341_/Q VGND VGND VPWR VPWR _6248_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2110 hold139/X VGND VGND VPWR VPWR _5745_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2121 _7262_/Q VGND VGND VPWR VPWR hold468/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2132 _4419_/X VGND VGND VPWR VPWR hold826/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5844__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6428__D _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2143 hold164/X VGND VGND VPWR VPWR _5790_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2154 _4241_/X VGND VGND VPWR VPWR hold818/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6179_ _7450_/Q _6144_/A _6116_/A _6317_/C _7514_/Q VGND VGND VPWR VPWR _6179_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1420 _5617_/X VGND VGND VPWR VPWR hold176/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2165 hold868/X VGND VGND VPWR VPWR _4224_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1431 hold181/X VGND VGND VPWR VPWR _5653_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2176 _7334_/Q VGND VGND VPWR VPWR hold388/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1442 _7202_/Q VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2187 _7662_/A VGND VGND VPWR VPWR hold480/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2198 _7350_/Q VGND VGND VPWR VPWR hold460/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1453 _5689_/X VGND VGND VPWR VPWR hold190/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1464 hold69/X VGND VGND VPWR VPWR _3461_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1475 _4201_/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1486 _4437_/X VGND VGND VPWR VPWR hold186/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3870__A3 _4521_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _5946_/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3430__A _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4280__A0 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4104__A_N _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5375__A3 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5780__A0 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_1__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6324__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5791__S _5793_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4335__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6088__B2 _7463_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6627__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5835__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_187_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5966__S hold13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3880_ _7376_/Q _3498_/X _3658_/X _7113_/Q VGND VGND VPWR VPWR _3880_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6563__A2 _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5550_ _5550_/A _5550_/B _5550_/C _5550_/D VGND VGND VPWR VPWR _5550_/Y sky130_fd_sc_hd__nand4_2
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6377__A1_N _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4501_ _5852_/A0 _4501_/A1 _4502_/S VGND VGND VPWR VPWR _4501_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5481_ _5481_/A _5481_/B _5481_/C VGND VGND VPWR VPWR _5560_/A sky130_fd_sc_hd__and3_1
XANTENNA__4747__A_N _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2353_A _7505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7220_ _4150_/A1 _7220_/D _6872_/X VGND VGND VPWR VPWR _7220_/Q sky130_fd_sc_hd__dfrtn_1
X_4432_ _4432_/A0 _5993_/A1 _4439_/S VGND VGND VPWR VPWR _4432_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7151_ _7151_/CLK _7151_/D fanout593/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfrtp_2
X_4363_ _4363_/A0 _5586_/A0 _4363_/S VGND VGND VPWR VPWR _4363_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3515__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6102_ _6102_/A _6102_/B _6102_/C _6102_/D VGND VGND VPWR VPWR _6102_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_111_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout518 _7592_/Q VGND VGND VPWR VPWR _6110_/A sky130_fd_sc_hd__clkbuf_16
X_7082_ _7505_/CLK _7082_/D fanout601/X VGND VGND VPWR VPWR _7662_/A sky130_fd_sc_hd__dfrtp_1
X_4294_ _4302_/S _4294_/B VGND VGND VPWR VPWR _4294_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5826__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6033_ _6119_/A _6028_/Y _6106_/B _6032_/B _6051_/C VGND VGND VPWR VPWR _6033_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4991__D _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_174_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4346__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2987_A _7123_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6251__B2 _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_3__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _7556_/CLK _6935_/D fanout594/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5876__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3604__A3 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6866_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6866_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout436_A _6093_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5817_ _5817_/A0 _5997_/A1 _5820_/S VGND VGND VPWR VPWR _5817_/X sky130_fd_sc_hd__mux2_1
X_6797_ _7111_/Q _6794_/Y _6795_/Y _7109_/Q _4430_/C VGND VGND VPWR VPWR _6797_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6554__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5762__A0 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5748_ _5748_/A0 _5991_/A1 _5748_/S VGND VGND VPWR VPWR _5748_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout603_A fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5679_ _5679_/A0 _5967_/A1 _5685_/S VGND VGND VPWR VPWR _5679_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7418_ _7555_/CLK _7418_/D fanout594/X VGND VGND VPWR VPWR _7418_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7349_ _7501_/CLK _7349_/D fanout581/X VGND VGND VPWR VPWR _7349_/Q sky130_fd_sc_hd__dfrtp_4
Xhold550 hold550/A VGND VGND VPWR VPWR _7417_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold561 hold561/A VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold572 hold572/A VGND VGND VPWR VPWR hold572/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3425__A _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold583 hold583/A VGND VGND VPWR VPWR _7390_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1718_A _7578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold594 hold594/A VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3540__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5817__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5640__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6490__B2 _7560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input136_A wb_dat_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1250 hold3095/X VGND VGND VPWR VPWR hold3096/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1261 _4401_/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1272 hold3111/X VGND VGND VPWR VPWR hold3112/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 _5582_/X VGND VGND VPWR VPWR _7209_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1294 hold3086/X VGND VGND VPWR VPWR hold3087/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5786__S _5793_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4703__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4308__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5808__A1 hold84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5284__A2 _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6481__B2 _7336_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput170 wb_we_i VGND VGND VPWR VPWR _6824_/C sky130_fd_sc_hd__buf_2
XANTENNA__3834__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4981_ _5339_/D _5138_/D _5034_/C VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__and3_2
XFILLER_0_187_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6720_ _7199_/Q _6463_/A _6771_/A3 _6463_/X _7164_/Q VGND VGND VPWR VPWR _6720_/X
+ sky130_fd_sc_hd__a32o_1
X_3932_ _7157_/Q hold56/A _5603_/B _3617_/X _7229_/Q VGND VGND VPWR VPWR _3932_/X
+ sky130_fd_sc_hd__a32o_1
X_6651_ _7036_/Q _6651_/B _6651_/C VGND VGND VPWR VPWR _6651_/X sky130_fd_sc_hd__and3_1
X_3863_ _3863_/A _5722_/A _4449_/B _5612_/B VGND VGND VPWR VPWR _3863_/X sky130_fd_sc_hd__and4_2
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6536__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5602_ _5602_/A0 _5863_/A0 _5602_/S VGND VGND VPWR VPWR _5602_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_143_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6582_ _7404_/Q _6409_/X _6420_/B _7308_/Q _6581_/X VGND VGND VPWR VPWR _6582_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3794_ _3744_/X _3750_/X _3794_/C _3794_/D VGND VGND VPWR VPWR _3795_/B sky130_fd_sc_hd__and4bb_4
XFILLER_0_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5533_ _5533_/A _5533_/B VGND VGND VPWR VPWR _5533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7539_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3770__A2 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5464_ _5294_/Y _5422_/X _5463_/X VGND VGND VPWR VPWR _5464_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7203_ _7206_/CLK _7203_/D _6780_/B VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfrtp_1
X_4415_ _4415_/A0 _4414_/X _4423_/S VGND VGND VPWR VPWR _4415_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5395_ _5395_/A1 _5113_/A wire529/X _5277_/X VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_10_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5511__A3 _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2902_A _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7134_ _7134_/CLK _7134_/D fanout588/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfstp_4
X_4346_ _5640_/B _5612_/C _4346_/C _5640_/D VGND VGND VPWR VPWR _4351_/S sky130_fd_sc_hd__and4_4
XANTENNA__3522__A2 _5875_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_75_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7231_/CLK sky130_fd_sc_hd__clkbuf_16
X_7065_ _7190_/CLK _7065_/D fanout573/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout359 hold400/X VGND VGND VPWR VPWR _5875_/A sky130_fd_sc_hd__buf_12
X_4277_ _4425_/C _6780_/B VGND VGND VPWR VPWR _4289_/S sky130_fd_sc_hd__nand2_8
XANTENNA__7513__RESET_B fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6016_ _7585_/Q _7586_/Q _6017_/D _7587_/Q VGND VGND VPWR VPWR _6018_/B sky130_fd_sc_hd__a31o_1
XANTENNA__6472__B2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3825__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6224__A1 _7468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6775__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__A2 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6918_ _7239_/CLK _6918_/D fanout566/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_92_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4250__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5619__B _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3994__C1 _3992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7134_/CLK sky130_fd_sc_hd__clkbuf_16
X_6849_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6849_/X sky130_fd_sc_hd__and2_1
XANTENNA__6527__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1570_A _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7521_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_115_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3761__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6160__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5502__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold380 hold380/A VGND VGND VPWR VPWR hold380/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3513__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold391 hold391/A VGND VGND VPWR VPWR _7247_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_189_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3816__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1080 hold2902/X VGND VGND VPWR VPWR hold2903/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 hold2923/X VGND VGND VPWR VPWR _7432_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6766__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6620__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6518__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4529__A1 _5805_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5248__C _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3752__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6151__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4200_ _4200_/A0 _5954_/A1 _4202_/S VGND VGND VPWR VPWR _4200_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6079__C _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2149_A _7451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5180_ _5180_/A _5180_/B _5216_/A VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__and3_1
Xhold2709 hold819/X VGND VGND VPWR VPWR _5586_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4131_ _6896_/Q _4131_/B VGND VGND VPWR VPWR _4132_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2316_A _7499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4062_ _4062_/A _4062_/B VGND VGND VPWR VPWR _4062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3512__B _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3807__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6206__A1 _7299_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6757__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4964_ _4963_/X _4960_/B _4855_/Y _4962_/Y VGND VGND VPWR VPWR _4964_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_0_59_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6703_ _6876_/Q _6600_/B _6459_/C _6421_/X _7008_/Q VGND VGND VPWR VPWR _6703_/X
+ sky130_fd_sc_hd__a32o_1
X_3915_ input35/X _5983_/A _5587_/C _5704_/A _7320_/Q VGND VGND VPWR VPWR _3915_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_80_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4895_ _4942_/A _5005_/A _5222_/B _4898_/C VGND VGND VPWR VPWR _4895_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__6509__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5717__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6634_ _7334_/Q _6423_/X _6454_/X _7494_/Q _6633_/X VGND VGND VPWR VPWR _6634_/X
+ sky130_fd_sc_hd__a221o_1
X_3846_ _4076_/B _4248_/S _3652_/X _7149_/Q _3845_/X VGND VGND VPWR VPWR _3846_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__3991__A2 _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3777_ _7282_/Q _3558_/X _3682_/X _7227_/Q _3776_/X VGND VGND VPWR VPWR _3782_/B
+ sky130_fd_sc_hd__a221o_4
X_6565_ _7307_/Q _6420_/B _6422_/X _7291_/Q VGND VGND VPWR VPWR _6565_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3743__A2 hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5516_ _5563_/A1 _4787_/Y _4946_/Y _4798_/Y _4709_/Y VGND VGND VPWR VPWR _5516_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_42_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6496_ _7280_/Q _6431_/Y _6775_/B1 VGND VGND VPWR VPWR _6496_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_112_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5447_ _4889_/A _4726_/Y _4889_/B _4888_/Y _5355_/D VGND VGND VPWR VPWR _5508_/A
+ sky130_fd_sc_hd__o41a_1
XANTENNA__6142__B1 _6090_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5378_ _4703_/Y _4844_/Y _4741_/Y _5451_/A1 VGND VGND VPWR VPWR _5378_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5902__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7117_ _7447_/CLK _7117_/D fanout598/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfrtp_4
X_4329_ _4329_/A0 _5714_/A0 _4333_/S VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_129_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7048_ _7176_/CLK _7048_/D fanout588/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6748__A2 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6452__C _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5420__A2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5708__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5068__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3982__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5184__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire546 wire546/A VGND VGND VPWR VPWR _4706_/A sky130_fd_sc_hd__buf_2
XANTENNA__6381__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input64_A mgmt_gpio_in[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6684__A1 _7027_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7435__RESET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4709__A _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6436__A1 _7319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6436__B2 _7511_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6739__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _7523_/Q _5785_/B _5938_/C _3673_/X _7201_/Q VGND VGND VPWR VPWR _3700_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_hold2099_A _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3973__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4680_ _5158_/A _5248_/A _5248_/B VGND VGND VPWR VPWR _4830_/A sky130_fd_sc_hd__and3_1
XFILLER_0_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3631_ _4173_/A _4248_/S _4231_/S input40/X _3630_/X VGND VGND VPWR VPWR _3632_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6372__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6350_ _7199_/Q _6332_/B _6079_/X _6072_/X _7154_/Q VGND VGND VPWR VPWR _6350_/X
+ sky130_fd_sc_hd__a32o_1
X_3562_ _5590_/A _3931_/D _5731_/B VGND VGND VPWR VPWR _3562_/X sky130_fd_sc_hd__and3_2
XANTENNA__3725__A2 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5301_ _5301_/A1 _4730_/Y _4731_/Y _5138_/Y _5300_/X VGND VGND VPWR VPWR _5405_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__6124__B1 _6122_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6281_ _6266_/X _6268_/X _6280_/Y VGND VGND VPWR VPWR _6281_/X sky130_fd_sc_hd__a21bo_4
X_3493_ _5803_/A _5590_/A _5640_/B VGND VGND VPWR VPWR _3493_/X sky130_fd_sc_hd__and3_2
Xhold3207 _7605_/Q VGND VGND VPWR VPWR _6192_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5232_ _4790_/C _4885_/X _4922_/B VGND VGND VPWR VPWR _5444_/D sky130_fd_sc_hd__a21oi_1
Xhold3218 _7602_/Q VGND VGND VPWR VPWR _6124_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3229 _7600_/Q VGND VGND VPWR VPWR _6064_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2506 _7153_/Q VGND VGND VPWR VPWR hold641/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_166_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5722__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2517 _7299_/Q VGND VGND VPWR VPWR hold128/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5163_ _5163_/A _5163_/B _5163_/C VGND VGND VPWR VPWR _5164_/B sky130_fd_sc_hd__nand3_1
Xhold2528 _7181_/Q VGND VGND VPWR VPWR hold126/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2539 _7178_/Q VGND VGND VPWR VPWR hold704/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1805 hold369/X VGND VGND VPWR VPWR _7338_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1816 _5833_/X VGND VGND VPWR VPWR hold421/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4114_ _4096_/X _4114_/B VGND VGND VPWR VPWR _4115_/B sky130_fd_sc_hd__nand2b_1
Xhold1827 _3449_/X VGND VGND VPWR VPWR _3500_/C sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_38_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5094_ _5094_/A _5096_/A VGND VGND VPWR VPWR _5473_/D sky130_fd_sc_hd__nand2_1
Xhold1838 _7017_/Q VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1849 hold506/X VGND VGND VPWR VPWR _4367_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4045_ _6910_/Q _6908_/Q _7071_/Q VGND VGND VPWR VPWR _4076_/C sky130_fd_sc_hd__and3_1
XANTENNA__5650__A2 hold284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _5996_/A0 _5996_/A1 hold37/X VGND VGND VPWR VPWR _5996_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_176_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_191_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4947_ _4948_/B _4948_/C _4947_/C _4954_/A VGND VGND VPWR VPWR _4947_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3964__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7666_ _7666_/A VGND VGND VPWR VPWR _7666_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout516_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4878_ _5213_/B _4954_/C _5183_/C _5213_/C VGND VGND VPWR VPWR _4906_/D sky130_fd_sc_hd__nand4_1
XFILLER_0_62_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6617_ _7565_/Q _6419_/C _6466_/X hold76/A _6601_/X VGND VGND VPWR VPWR _6617_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3829_ _7433_/Q _3525_/X _4485_/A _7144_/Q VGND VGND VPWR VPWR _3829_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6363__B1 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7597_ _7610_/CLK _7597_/D fanout568/X VGND VGND VPWR VPWR _7597_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_171_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6548_ _6547_/X _6572_/A2 _6573_/S VGND VGND VPWR VPWR _6548_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6115__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6479_ _7568_/Q _6424_/X _6474_/X _6478_/X _6430_/X VGND VGND VPWR VPWR _6479_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput260 _7224_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
Xoutput271 _6914_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_0_100_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput282 _7240_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
XANTENNA__5632__B _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4141__A2 _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput293 _6911_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_0_100_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6447__C _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3433__A _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6463__B _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_186_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_179_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3955__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5157__A1 _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6354__B1 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire365 _4145_/Y VGND VGND VPWR VPWR wire365/X sky130_fd_sc_hd__buf_6
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3707__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output268_A _7231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6657__A1 _7132_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6657__B2 _6988_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5969__S hold13/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4174__A _4174_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5850_ _5985_/A1 _5850_/A1 _5856_/S VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _4802_/A _4801_/B _4801_/C VGND VGND VPWR VPWR _4823_/B sky130_fd_sc_hd__and3_2
XFILLER_0_152_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6593__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5781_ _5997_/A1 _5781_/A1 hold49/X VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7520_ _7560_/CLK _7520_/D fanout599/X VGND VGND VPWR VPWR _7520_/Q sky130_fd_sc_hd__dfstp_4
X_4732_ _5038_/A _4822_/D _4755_/A _5005_/A VGND VGND VPWR VPWR _4732_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3946__A2 hold12/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold72_A hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7451_ _7505_/CLK _7451_/D fanout601/X VGND VGND VPWR VPWR _7451_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6345__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4663_ _4667_/A _4667_/B _4795_/C VGND VGND VPWR VPWR _4861_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3518__A _5785_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6402_ _6462_/D _6435_/B VGND VGND VPWR VPWR _6645_/C sky130_fd_sc_hd__nor2_8
X_3614_ _7548_/Q _5965_/A _4212_/A hold72/A _7564_/Q VGND VGND VPWR VPWR _3614_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_0_153_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4594_ _4825_/A _5071_/B _5071_/C _4755_/A VGND VGND VPWR VPWR _4594_/Y sky130_fd_sc_hd__nor4_2
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7382_ _7581_/CLK _7382_/D fanout584/X VGND VGND VPWR VPWR _7382_/Q sky130_fd_sc_hd__dfrtp_4
Xhold902 hold902/A VGND VGND VPWR VPWR _7324_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6360__A3 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold913 hold913/A VGND VGND VPWR VPWR hold913/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3545_ _5590_/A _5640_/B _5731_/B VGND VGND VPWR VPWR _3545_/X sky130_fd_sc_hd__and3_4
XFILLER_0_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold924 hold924/A VGND VGND VPWR VPWR _7284_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6333_ _7194_/Q _6144_/A _6120_/B _6379_/B1 _7189_/Q VGND VGND VPWR VPWR _6333_/X
+ sky130_fd_sc_hd__a32o_1
Xhold935 hold935/A VGND VGND VPWR VPWR hold935/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold946 _4326_/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold957 hold957/A VGND VGND VPWR VPWR hold957/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold968 _4207_/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3004 hold3004/A VGND VGND VPWR VPWR _5841_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6648__B2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6264_ _7294_/Q _6144_/A _6144_/B _6074_/X _7302_/Q VGND VGND VPWR VPWR _6264_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3015 hold3015/A VGND VGND VPWR VPWR _4411_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold979 hold979/A VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3476_ hold280/X hold53/X VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__nand2b_1
Xhold3026 hold751/X VGND VGND VPWR VPWR _5601_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5215_ _4622_/Y _4709_/Y _4726_/Y _5214_/X VGND VGND VPWR VPWR _5223_/A sky130_fd_sc_hd__o31a_1
Xhold3037 _7250_/Q VGND VGND VPWR VPWR hold736/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2303 _7284_/Q VGND VGND VPWR VPWR hold923/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3048 _7040_/Q VGND VGND VPWR VPWR hold720/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5320__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2314 _5724_/X VGND VGND VPWR VPWR hold587/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3059 _6941_/Q VGND VGND VPWR VPWR hold3059/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6195_ _7499_/Q _6094_/A _6084_/X _6116_/X _7315_/Q VGND VGND VPWR VPWR _6195_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2325 _7009_/Q VGND VGND VPWR VPWR hold931/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2336 hold913/X VGND VGND VPWR VPWR _4398_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1602 _7530_/Q VGND VGND VPWR VPWR hold235/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5146_ _5404_/C _5410_/B _4977_/X _4776_/A VGND VGND VPWR VPWR _5308_/A sky130_fd_sc_hd__a31o_1
Xhold2347 hold925/X VGND VGND VPWR VPWR _4531_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2358 hold629/X VGND VGND VPWR VPWR _4366_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1613 _7556_/Q VGND VGND VPWR VPWR hold255/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2369 _7540_/Q VGND VGND VPWR VPWR hold929/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1624 _6951_/Q VGND VGND VPWR VPWR hold249/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3882__A1 _7352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5879__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1635 _5962_/X VGND VGND VPWR VPWR hold262/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1646 hold258/X VGND VGND VPWR VPWR _7362_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5077_ _5387_/C _5077_/B VGND VGND VPWR VPWR _5077_/Y sky130_fd_sc_hd__nand2_4
Xhold1657 hold290/X VGND VGND VPWR VPWR _5780_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout466_A hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1668 _5843_/X VGND VGND VPWR VPWR hold246/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1679 _5989_/X VGND VGND VPWR VPWR hold234/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6820__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4028_ _4028_/A0 _4027_/Y _4040_/A VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6820__B2 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3634__B2 _7508_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4515__C hold56/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6179__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5979_ _5979_/A0 _5979_/A1 _5982_/S VGND VGND VPWR VPWR _5979_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3937__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7649_ _7649_/A VGND VGND VPWR VPWR _7649_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6336__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3428__A _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6639__A1 _7350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input166_A wb_sel_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6103__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4259__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2870 _6984_/Q VGND VGND VPWR VPWR _4298_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5789__S _5793_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input27_A mask_rev_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2881 hold2881/A VGND VGND VPWR VPWR _5903_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2892 _7197_/Q VGND VGND VPWR VPWR hold2892/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6811__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6811__B2 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3625__B2 _7524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4968__A4 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_168_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5378__A1 _4703_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6575__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4722__A _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5393__A4 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_user_clock user_clock VGND VGND VPWR VPWR clkbuf_0_user_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6342__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold209 hold209/A VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6084__A_N _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5138_/D _5038_/C _5216_/A VGND VGND VPWR VPWR _5026_/B sky130_fd_sc_hd__and3_1
XANTENNA__6087__C _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6802__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6802__B2 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6951_ _7551_/CLK _6951_/D fanout595/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4616__B _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3520__B _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5902_ _5902_/A _5902_/B VGND VGND VPWR VPWR _5910_/S sky130_fd_sc_hd__nand2_8
XANTENNA_hold2598_A _7512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6882_ _7075_/CLK _6882_/D _6832_/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5369__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5833_ _5833_/A0 _5896_/A0 _5838_/S VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_159_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6566__B1 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3919__A2 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5764_ _5953_/A1 _5764_/A1 _5766_/S VGND VGND VPWR VPWR _5764_/X sky130_fd_sc_hd__mux2_1
X_7503_ _7521_/CLK _7503_/D fanout601/X VGND VGND VPWR VPWR _7503_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4715_ _4795_/C _4909_/D _4805_/B _4740_/D VGND VGND VPWR VPWR _4715_/Y sky130_fd_sc_hd__nor4b_2
XANTENNA__6318__B1 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5695_ _5983_/A _5731_/B _5902_/B VGND VGND VPWR VPWR _5703_/S sky130_fd_sc_hd__and3_4
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7434_ _7556_/CLK _7434_/D fanout594/X VGND VGND VPWR VPWR _7434_/Q sky130_fd_sc_hd__dfrtp_4
X_4646_ _4646_/A _4646_/B VGND VGND VPWR VPWR _4646_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6333__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold710 hold710/A VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4577_ _4795_/C _4740_/D _4772_/A VGND VGND VPWR VPWR _4578_/B sky130_fd_sc_hd__nand3_4
X_7365_ _7366_/CLK _7365_/D fanout579/X VGND VGND VPWR VPWR _7365_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold721 _4369_/X VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold732 hold732/A VGND VGND VPWR VPWR hold732/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_102_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap451 _5113_/B VGND VGND VPWR VPWR _5118_/B sky130_fd_sc_hd__clkbuf_2
Xhold743 hold743/A VGND VGND VPWR VPWR _7475_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6316_ _6875_/Q _6112_/X _6121_/X _6989_/Q _6315_/X VGND VGND VPWR VPWR _6316_/X
+ sky130_fd_sc_hd__a221o_1
Xhold754 _4276_/X VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3528_ _7510_/Q _5983_/A _5947_/B _3527_/X _6918_/Q VGND VGND VPWR VPWR _3528_/X
+ sky130_fd_sc_hd__a32o_4
Xhold765 hold765/A VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold776 hold776/A VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7296_ _7539_/CLK _7296_/D fanout577/X VGND VGND VPWR VPWR _7296_/Q sky130_fd_sc_hd__dfstp_2
Xhold787 hold787/A VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold798 _4478_/X VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2100 hold655/X VGND VGND VPWR VPWR _4202_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6247_ _7317_/Q _6116_/X _6121_/X _7309_/Q _6246_/X VGND VGND VPWR VPWR _6257_/A
+ sky130_fd_sc_hd__a221o_1
X_3459_ _3511_/C _3557_/B _3557_/C VGND VGND VPWR VPWR _3564_/A sky130_fd_sc_hd__and3_4
Xhold2111 _5745_/X VGND VGND VPWR VPWR hold140/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2122 hold468/X VGND VGND VPWR VPWR _5639_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2133 _6949_/Q VGND VGND VPWR VPWR hold538/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2144 _5790_/X VGND VGND VPWR VPWR hold165/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1410 _5995_/X VGND VGND VPWR VPWR hold1410/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6178_ _6116_/B _6172_/X _6175_/X _6177_/X VGND VGND VPWR VPWR _6178_/X sky130_fd_sc_hd__a211o_4
Xhold2155 _7045_/Q VGND VGND VPWR VPWR hold160/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1421 hold176/X VGND VGND VPWR VPWR _7246_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2166 _4224_/X VGND VGND VPWR VPWR hold869/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1432 _5653_/X VGND VGND VPWR VPWR hold182/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2177 hold388/X VGND VGND VPWR VPWR _5721_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2188 hold480/X VGND VGND VPWR VPWR _4421_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1443 hold10/X VGND VGND VPWR VPWR _3468_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5129_ _5410_/A _4815_/B _5399_/C _5047_/A VGND VGND VPWR VPWR _5317_/A sky130_fd_sc_hd__a31o_1
Xhold2199 hold460/X VGND VGND VPWR VPWR _5739_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1454 hold190/X VGND VGND VPWR VPWR _7305_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1465 _3461_/X VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1476 hold16/X VGND VGND VPWR VPWR hold1476/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 _7206_/Q VGND VGND VPWR VPWR hold130/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 hold24/X VGND VGND VPWR VPWR _7534_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6557__B1 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6460__C _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7208__RESET_B _6780_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7645__CLK _4164_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6088__A2 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3846__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__buf_2
XFILLER_0_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_188_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5599__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6651__B _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5220__B1 _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6563__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5771__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4500_ _5914_/A1 _4500_/A1 _4502_/S VGND VGND VPWR VPWR _4500_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5480_ _4703_/Y _4826_/Y _4832_/Y _4846_/Y _4709_/Y VGND VGND VPWR VPWR _5481_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_41_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6315__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1 _3526_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4431_ _5785_/B _5992_/C _5992_/D VGND VGND VPWR VPWR _4439_/S sky130_fd_sc_hd__and3_4
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6720__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4362_ _4362_/A0 _5852_/A0 _4363_/S VGND VGND VPWR VPWR _4362_/X sky130_fd_sc_hd__mux2_1
X_7150_ _7395_/CLK _7150_/D fanout598/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3515__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6101_ _7351_/Q _6099_/X _6100_/X _7471_/Q _6098_/X VGND VGND VPWR VPWR _6102_/D
+ sky130_fd_sc_hd__a221o_1
X_7081_ _7505_/CLK _7081_/D fanout601/X VGND VGND VPWR VPWR _7661_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout519 _7592_/Q VGND VGND VPWR VPWR _6094_/A sky130_fd_sc_hd__clkbuf_16
X_4293_ _3922_/Y _4293_/A1 _4302_/S VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_0__1111_ _3733_/X VGND VGND VPWR VPWR clkbuf_0__1111_/X sky130_fd_sc_hd__clkbuf_16
X_6032_ _6106_/B _6032_/B VGND VGND VPWR VPWR _6032_/Y sky130_fd_sc_hd__nor2_8
XFILLER_0_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3531__A _5722_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4346__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6251__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5054__A3 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6934_ _7551_/CLK _6934_/D fanout595/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4262__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6865_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6865_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6539__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6003__A2 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5816_ _5816_/A0 _5987_/A1 _5820_/S VGND VGND VPWR VPWR _5816_/X sky130_fd_sc_hd__mux2_1
X_6796_ _6824_/C _6825_/A3 _7110_/Q VGND VGND VPWR VPWR _6798_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5747_ _5747_/A0 _5999_/A1 _5748_/S VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_146_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7673__A _7673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5678_ _5678_/A0 _5903_/A0 _5685_/S VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7417_ _7417_/CLK _7417_/D fanout586/X VGND VGND VPWR VPWR _7417_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_130_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4629_ _4814_/C _4568_/Y _5301_/A1 _4627_/Y VGND VGND VPWR VPWR _4768_/B sky130_fd_sc_hd__o31a_4
XANTENNA__6711__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1446_A _3537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold540 hold540/A VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4301__S _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7348_ _7478_/CLK _7348_/D fanout580/X VGND VGND VPWR VPWR _7348_/Q sky130_fd_sc_hd__dfrtp_4
Xhold551 hold551/A VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold562 _5733_/X VGND VGND VPWR VPWR _7344_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold573 _4343_/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold584 hold584/A VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold595 hold595/A VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7279_ _7309_/CLK _7279_/D fanout576/X VGND VGND VPWR VPWR _7279_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_hold1613_A _7556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5640__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6490__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3441__A _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1240 hold3082/X VGND VGND VPWR VPWR hold3083/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6455__C _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1251 hold3097/X VGND VGND VPWR VPWR _7543_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1262 hold3076/X VGND VGND VPWR VPWR hold3077/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1273 _4516_/X VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input129_A wb_adr_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1284 hold3150/X VGND VGND VPWR VPWR hold3151/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 _4341_/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6242__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input94_A uart_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5753__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5505__A1 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6481__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6818_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4492__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6218__C1 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6769__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6233__A2 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4244__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4980_ _4984_/B _4984_/A _4660_/Y _4690_/Y VGND VGND VPWR VPWR _4980_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_175_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3931_ _7162_/Q _4509_/A _5612_/C _3931_/D VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__and4_1
XFILLER_0_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4714__A_N _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6650_ _6649_/X _6675_/A2 _6777_/S VGND VGND VPWR VPWR _7622_/D sky130_fd_sc_hd__mux2_1
X_3862_ _7236_/Q _5612_/B _5603_/B VGND VGND VPWR VPWR _3862_/X sky130_fd_sc_hd__and3_2
XFILLER_0_85_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6536__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5601_ _5601_/A0 _5754_/A1 _5602_/S VGND VGND VPWR VPWR _5601_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5744__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6581_ _7340_/Q _6425_/X _6454_/X _7492_/Q _6580_/X VGND VGND VPWR VPWR _6581_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3793_ _3764_/X _3773_/X _3793_/C _3793_/D VGND VGND VPWR VPWR _3794_/D sky130_fd_sc_hd__and4bb_4
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5532_ _5532_/A _5532_/B _5532_/C _5532_/D VGND VGND VPWR VPWR _5533_/B sky130_fd_sc_hd__and4_1
XFILLER_0_14_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7213_/CLK sky130_fd_sc_hd__clkbuf_16
X_5463_ _5462_/X _5460_/X _5442_/X _5441_/X VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__3770__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3526__A _3537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7202_ _7206_/CLK _7202_/D _6780_/B VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_1
X_4414_ _4444_/A0 _5996_/A1 _4422_/S VGND VGND VPWR VPWR _4414_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5394_ _5394_/A _5476_/B _5394_/C VGND VGND VPWR VPWR _5394_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7133_ _7186_/CLK _7133_/D _6833_/A VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfrtp_4
X_4345_ _5754_/A1 _4345_/A1 _4345_/S VGND VGND VPWR VPWR _4345_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3522__A3 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7064_ _7190_/CLK _7064_/D fanout573/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_4
X_4276_ _4276_/A0 _5586_/A0 _4276_/S VGND VGND VPWR VPWR _4276_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6908__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6015_ _6018_/A _6015_/B _6015_/C VGND VGND VPWR VPWR _7586_/D sky130_fd_sc_hd__and3_1
XFILLER_0_185_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4483__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4076__B _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6224__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ _7239_/CLK _6917_/D fanout566/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6848_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6848_/X sky130_fd_sc_hd__and2_1
XANTENNA__5619__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6527__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5735__A1 _5735_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6779_ _7108_/D _4115_/B _6778_/Y _6779_/B2 VGND VGND VPWR VPWR _6779_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold1563_A _7524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3761__A3 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold370 hold370/A VGND VGND VPWR VPWR hold370/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold381 _5951_/X VGND VGND VPWR VPWR _7538_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3513__A3 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold392 hold392/A VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5671__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4474__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 hold2832/X VGND VGND VPWR VPWR hold2833/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5797__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1081 _4462_/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1092 hold2933/X VGND VGND VPWR VPWR hold2934/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4714__B _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4887__A_N _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5726__A1 _5987_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output298_A _7247_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4130_ _4130_/A VGND VGND VPWR VPWR _4130_/Y sky130_fd_sc_hd__inv_2
X_4061_ _7071_/Q _3856_/A _4057_/S _4067_/C VGND VGND VPWR VPWR _4062_/B sky130_fd_sc_hd__a211o_2
XANTENNA__4465__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2211_A _7470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3512__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6206__A2 _6022_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4217__A1 hold464/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_176_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4624__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4963_ _4571_/Y _5073_/B _4843_/A VGND VGND VPWR VPWR _4963_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_175_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6702_ _7174_/Q _6747_/B _6747_/C VGND VGND VPWR VPWR _6702_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3914_ _7552_/Q _5965_/A hold12/A _3501_/X _7576_/Q VGND VGND VPWR VPWR _3914_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4894_ _4932_/B _5213_/C _5260_/D _4940_/D VGND VGND VPWR VPWR _4894_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6633_ _7374_/Q _6404_/Y _6651_/C _6422_/X _7294_/Q VGND VGND VPWR VPWR _6633_/X
+ sky130_fd_sc_hd__a32o_1
X_3845_ input54/X _5785_/B _4491_/B hold72/A _7561_/Q VGND VGND VPWR VPWR _3845_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3991__A3 _5911_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3728__B1 hold72/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6331__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6564_ _7299_/Q _6420_/A _6454_/X hold96/A _6563_/X VGND VGND VPWR VPWR _6569_/B
+ sky130_fd_sc_hd__a221o_1
X_3776_ _6965_/Q _5603_/B _5640_/C _3657_/X _6960_/Q VGND VGND VPWR VPWR _3776_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_144_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_756 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5515_ _5294_/C _5294_/A _5294_/B _5493_/Y _5514_/X VGND VGND VPWR VPWR _5515_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_125_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6495_ _6479_/X _6495_/B _6495_/C VGND VGND VPWR VPWR _6495_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_131_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5446_ _4737_/Y _5065_/Y _5355_/B _5223_/A _4897_/X VGND VGND VPWR VPWR _5448_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__6142__B2 _7376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6693__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5377_ _5255_/X _4844_/Y _4703_/Y _4717_/Y VGND VGND VPWR VPWR _5384_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_10_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A _5903_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3900__B1 _3675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7116_ _7134_/CLK _7116_/D fanout588/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_4
X_4328_ _4449_/B _4388_/B _4346_/C _5640_/D VGND VGND VPWR VPWR _4333_/S sky130_fd_sc_hd__and4_4
XANTENNA_input1_A debug_mode VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6445__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7047_ _7151_/CLK _7047_/D fanout588/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_4
X_4259_ _5640_/B _5612_/C _5640_/C _5640_/D VGND VGND VPWR VPWR _4264_/S sky130_fd_sc_hd__and4_2
XANTENNA__6880__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5653__A0 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4456__A1 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4208__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4815__A _5387_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1680_A _7436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3982__A3 _3519_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire536 _5118_/C VGND VGND VPWR VPWR wire536/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5184__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4392__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input57_A mgmt_gpio_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6684__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5812__C hold48/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4709__B _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6436__A2 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4447__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5644__A0 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_74_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7255_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3973__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3630_ _7380_/Q _5803_/A _5983_/A _3503_/X input31/X VGND VGND VPWR VPWR _3630_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4383__A0 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3561_ hold36/X _5590_/A _5731_/B VGND VGND VPWR VPWR _5713_/A sky130_fd_sc_hd__and3_4
XANTENNA__3725__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5300_ _4956_/A _4709_/Y _4687_/Y _4605_/Y VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6280_ _6280_/A _6280_/B _6280_/C _6280_/D VGND VGND VPWR VPWR _6280_/Y sky130_fd_sc_hd__nor4_1
XANTENNA__3507__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3492_ _3505_/C _3505_/D _5590_/A VGND VGND VPWR VPWR _3492_/X sky130_fd_sc_hd__and3_4
XFILLER_0_11_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5231_ _5231_/A _5231_/B _5231_/C VGND VGND VPWR VPWR _5235_/A sky130_fd_sc_hd__nor3_1
Xhold3208 _6192_/X VGND VGND VPWR VPWR _7605_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3219 _7603_/Q VGND VGND VPWR VPWR _6169_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2507 hold641/X VGND VGND VPWR VPWR _4499_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5722__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2518 hold128/X VGND VGND VPWR VPWR _5682_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5162_ _4748_/Y _5528_/A3 _4826_/Y _4814_/Y VGND VGND VPWR VPWR _5491_/C sky130_fd_sc_hd__a211o_1
Xhold2529 hold126/X VGND VGND VPWR VPWR _4532_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_12_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7112_/CLK sky130_fd_sc_hd__clkbuf_16
X_4113_ _4121_/A _4047_/S _3400_/Y _4113_/B1 VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__a31o_1
Xhold1806 _7457_/Q VGND VGND VPWR VPWR hold412/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5093_ _4707_/Y _4946_/Y _5092_/Y VGND VGND VPWR VPWR _5093_/Y sky130_fd_sc_hd__o21ai_1
Xhold1817 _7175_/Q VGND VGND VPWR VPWR hold376/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4438__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1828 hold280/X VGND VGND VPWR VPWR _3511_/C sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5635__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1839 hold65/X VGND VGND VPWR VPWR _4342_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4044_ _4044_/A1 _4040_/D _4014_/B _4043_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_79_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6834__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5650__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7563_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_189_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_188_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5995_ _5995_/A0 _5995_/A1 hold37/A VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__mux2_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4946_ _5091_/A _5072_/B VGND VGND VPWR VPWR _4946_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_86_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_191_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7665_ _7665_/A VGND VGND VPWR VPWR _7665_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4877_ _4877_/A _5180_/B VGND VGND VPWR VPWR _5185_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6616_ _7445_/Q _6574_/B _6771_/A3 _6443_/X _7453_/Q VGND VGND VPWR VPWR _6616_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3828_ _3828_/A _3828_/B _3828_/C _3828_/D VGND VGND VPWR VPWR _3854_/A sky130_fd_sc_hd__nor4_1
XANTENNA_fanout411_A _4491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7596_ _7610_/CLK _7596_/D fanout567/X VGND VGND VPWR VPWR _7596_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5020__D1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4374__A0 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6547_ _6649_/S _7617_/Q _6545_/Y _6546_/X VGND VGND VPWR VPWR _6547_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3759_ _3759_/A _3759_/B _3759_/C _3759_/D VGND VGND VPWR VPWR _3794_/C sky130_fd_sc_hd__nor4_2
XFILLER_0_30_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6115__A1 _7447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6115__B2 _7519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6478_ _7400_/Q _6409_/X _6476_/X _6477_/X VGND VGND VPWR VPWR _6478_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6666__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5323__C1 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5429_ _5113_/A _5094_/A _5260_/D _5107_/A VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__o31a_1
Xoutput250 _4130_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
XFILLER_0_11_770 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput261 _7225_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
Xoutput272 _6915_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput283 _7241_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
Xoutput294 _6912_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_0_100_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6463__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input111_A wb_adr_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5079__C _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6354__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire344 _3888_/Y VGND VGND VPWR VPWR _3922_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3707__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6657__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5865__A0 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6290__B1 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4455__A _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6092__D _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4800_/A _4800_/B _4800_/C VGND VGND VPWR VPWR _4800_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_158_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ _5987_/A1 _5780_/A1 hold49/X VGND VGND VPWR VPWR _5780_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5396__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _5138_/A _4822_/D VGND VGND VPWR VPWR _4731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3946__A3 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7450_ _7505_/CLK _7450_/D fanout601/X VGND VGND VPWR VPWR _7450_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6345__A1 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4662_ _4984_/A _4984_/B _4660_/Y VGND VGND VPWR VPWR _4996_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5002__D1 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6401_ _6400_/X _6401_/A1 _6777_/S VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3613_ _7556_/Q _3508_/X _5920_/A _7516_/Q _3612_/X VGND VGND VPWR VPWR _3623_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3518__B hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7381_ _7429_/CLK _7381_/D fanout583/X VGND VGND VPWR VPWR _7381_/Q sky130_fd_sc_hd__dfrtp_4
X_4593_ _4593_/A _4825_/A VGND VGND VPWR VPWR _4593_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_153_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold903 hold903/A VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6332_ _7068_/Q _6332_/B _6332_/C VGND VGND VPWR VPWR _6332_/X sky130_fd_sc_hd__and3_1
Xhold914 hold914/A VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3544_ _5722_/A _4509_/A _3931_/D VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__and3_4
Xhold925 hold925/A VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold936 _5914_/X VGND VGND VPWR VPWR _7505_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold947 hold947/A VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold958 _4494_/X VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold969 hold969/A VGND VGND VPWR VPWR hold969/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6263_ _7318_/Q _6116_/C _6116_/A _6262_/X VGND VGND VPWR VPWR _6263_/X sky130_fd_sc_hd__a31o_1
Xhold3005 _5841_/X VGND VGND VPWR VPWR hold3005/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3475_ _4429_/B hold52/X _3453_/X VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__o21a_1
Xhold3016 _7228_/Q VGND VGND VPWR VPWR hold738/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5856__A0 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3027 _5601_/X VGND VGND VPWR VPWR hold752/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5214_ _4622_/Y _4726_/Y _4946_/Y _4898_/Y VGND VGND VPWR VPWR _5214_/X sky130_fd_sc_hd__o31a_1
Xhold3038 hold736/X VGND VGND VPWR VPWR _5624_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_50_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2304 hold923/X VGND VGND VPWR VPWR _5665_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3049 hold720/X VGND VGND VPWR VPWR _4369_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6194_ _7323_/Q _6082_/X _6120_/X _7339_/Q _6193_/X VGND VGND VPWR VPWR _6212_/A
+ sky130_fd_sc_hd__a221o_1
Xhold2315 hold587/X VGND VGND VPWR VPWR _7336_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2326 hold931/X VGND VGND VPWR VPWR _4332_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2337 _4398_/X VGND VGND VPWR VPWR hold914/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1603 hold235/X VGND VGND VPWR VPWR _5942_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2348 _7160_/Q VGND VGND VPWR VPWR hold927/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5145_ _5145_/A _5145_/B _5145_/C VGND VGND VPWR VPWR _5148_/A sky130_fd_sc_hd__nand3_1
Xhold1614 hold255/X VGND VGND VPWR VPWR _5971_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2359 _7339_/Q VGND VGND VPWR VPWR hold106/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1625 hold249/X VGND VGND VPWR VPWR _4253_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3882__A2 _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1636 hold262/X VGND VGND VPWR VPWR _7548_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1647 _7240_/Q VGND VGND VPWR VPWR hold273/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5076_ _5260_/C _5070_/X _5075_/Y VGND VGND VPWR VPWR _5084_/A sky130_fd_sc_hd__a21oi_1
Xhold1658 _5780_/X VGND VGND VPWR VPWR hold291/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1669 _6924_/Q VGND VGND VPWR VPWR _4209_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4027_ _4025_/A _4017_/B _4026_/Y _3447_/Y VGND VGND VPWR VPWR _4027_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__3634__A2 _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6033__B1 _6106_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5895__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4515__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6584__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5978_ _5987_/A1 _5978_/A1 _5982_/S VGND VGND VPWR VPWR _5978_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_177_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4929_ _4929_/A _5038_/C _5342_/B VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3937__A3 _3669_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7648_ _7648_/A VGND VGND VPWR VPWR _7648_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6336__A1 _6969_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6336__B2 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7579_ _7580_/CLK _7579_/D fanout597/X VGND VGND VPWR VPWR _7579_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1643_A _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmgmt_gpio_9_buff_inst _4150_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_8
XANTENNA__6639__A2 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3444__A _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7067__RESET_B fanout606/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1908_A _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input159_A wb_dat_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4259__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2860 _7636_/Q VGND VGND VPWR VPWR _6792_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2871 hold2871/A VGND VGND VPWR VPWR hold2871/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2882 _6986_/Q VGND VGND VPWR VPWR _4301_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5075__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2893 hold2893/A VGND VGND VPWR VPWR _4552_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6272__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5378__A2 _4844_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4722__B _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_182_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6950_ _7575_/CLK _6950_/D fanout595/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3520__C _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5901_ _5991_/A1 _5901_/A1 _5901_/S VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__mux2_1
X_6881_ _6881_/CLK _6881_/D _4079_/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5832_ _5832_/A0 _5985_/A1 _5838_/S VGND VGND VPWR VPWR _5832_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5369__A2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6566__B2 _7539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5763_ _5997_/A1 _5763_/A1 _5766_/S VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7502_ _7580_/CLK _7502_/D fanout594/X VGND VGND VPWR VPWR _7502_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3529__A hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4714_ _4795_/C _4740_/D VGND VGND VPWR VPWR _5079_/B sky130_fd_sc_hd__and2b_4
XANTENNA_hold2758_A _7116_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5694_ _5955_/A1 _5694_/A1 _5694_/S VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6318__B2 _7178_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7433_ _7457_/CLK _7433_/D fanout586/X VGND VGND VPWR VPWR _7433_/Q sky130_fd_sc_hd__dfrtp_4
X_4645_ _4675_/B _5089_/B _4675_/A _4645_/D VGND VGND VPWR VPWR _4646_/B sky130_fd_sc_hd__nand4_4
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold700 hold700/A VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7364_ _7501_/CLK _7364_/D fanout581/X VGND VGND VPWR VPWR _7364_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_141_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4576_ _4615_/A _4668_/C VGND VGND VPWR VPWR _4861_/A sky130_fd_sc_hd__nand2_2
Xhold711 _5772_/X VGND VGND VPWR VPWR _7379_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold722 hold722/A VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold733 hold733/A VGND VGND VPWR VPWR _7365_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold744 hold744/A VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6315_ _7057_/Q _6110_/A _6084_/X _6075_/X _7163_/Q VGND VGND VPWR VPWR _6315_/X
+ sky130_fd_sc_hd__a32o_1
X_3527_ _5590_/A _5640_/B _5612_/B VGND VGND VPWR VPWR _3527_/X sky130_fd_sc_hd__and3_2
Xhold755 hold755/A VGND VGND VPWR VPWR hold755/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7295_ _7539_/CLK _7295_/D fanout577/X VGND VGND VPWR VPWR _7295_/Q sky130_fd_sc_hd__dfstp_2
Xhold766 _4357_/X VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold777 hold777/A VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold788 _5608_/X VGND VGND VPWR VPWR _7239_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7160__RESET_B _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6246_ _7517_/Q _6332_/B _6073_/X _6085_/X _7501_/Q VGND VGND VPWR VPWR _6246_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold799 hold799/A VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3458_ _4429_/B _3458_/A2 _3456_/X VGND VGND VPWR VPWR _3458_/Y sky130_fd_sc_hd__a21oi_4
Xhold2101 _4202_/X VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2112 hold140/X VGND VGND VPWR VPWR _7355_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4501__A0 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2123 _5639_/X VGND VGND VPWR VPWR hold469/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6177_ _7314_/Q _6116_/X _6119_/X _7402_/Q _6176_/X VGND VGND VPWR VPWR _6177_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2134 hold538/X VGND VGND VPWR VPWR _4251_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1400 _6885_/Q VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout576_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2145 hold165/X VGND VGND VPWR VPWR _7395_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2156 hold160/X VGND VGND VPWR VPWR _4375_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1411 hold1411/A VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2167 _6925_/Q VGND VGND VPWR VPWR hold847/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1422 _7329_/Q VGND VGND VPWR VPWR hold193/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1433 hold182/X VGND VGND VPWR VPWR _7273_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5128_ _4695_/Y _4732_/Y _5531_/D _5531_/C VGND VGND VPWR VPWR _5163_/A sky130_fd_sc_hd__o211a_1
Xhold2178 _7670_/A VGND VGND VPWR VPWR hold885/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2189 _4421_/X VGND VGND VPWR VPWR hold481/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1444 _3467_/Y VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1455 _7270_/Q VGND VGND VPWR VPWR hold177/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6254__B1 _7469_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1466 hold70/X VGND VGND VPWR VPWR _3505_/C sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4095__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1477 hold1477/A VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1488 hold130/X VGND VGND VPWR VPWR _3458_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5059_ _5107_/A _5059_/B _5399_/D VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__and3_2
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 _7444_/Q VGND VGND VPWR VPWR hold173/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4823__A _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6557__B2 _7467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6460__D _6651_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3439__A _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6309__A1 _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_180_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6190__C1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6493__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3846__A2 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__buf_2
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6245__B1 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2690 hold763/X VGND VGND VPWR VPWR _4550_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_98_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6651__C _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4430_ _7105_/D _4430_/B _4430_/C _4430_/D VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__nand4b_1
XANTENNA_2 _3614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6720__A1 _7199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5523__A2 _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4361_ _4361_/A0 _5914_/A1 _4363_/S VGND VGND VPWR VPWR _4361_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6100_ _6106_/B _6116_/C _6332_/B _6119_/A VGND VGND VPWR VPWR _6100_/X sky130_fd_sc_hd__and4b_4
X_7080_ _7197_/CLK _7080_/D fanout601/X VGND VGND VPWR VPWR _7660_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__3515__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4292_ _4302_/S _3996_/B _4291_/Y VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__6484__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6031_ _6119_/A _6116_/C VGND VGND VPWR VPWR _6032_/B sky130_fd_sc_hd__nand2_4
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3531__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6787__A1 _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4346__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6933_ _6956_/CLK _6933_/D fanout603/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6864_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6864_/X sky130_fd_sc_hd__and2_1
XANTENNA__6539__A1 _7546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6539__B2 _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5815_ _5815_/A0 _5815_/A1 _5820_/S VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6795_ _6824_/C _6795_/B VGND VGND VPWR VPWR _6795_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5746_ _5746_/A0 _5953_/A1 _5748_/S VGND VGND VPWR VPWR _5746_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3773__A1 _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5677_ hold12/X _5731_/B hold47/X VGND VGND VPWR VPWR _5685_/S sky130_fd_sc_hd__and3_4
X_7416_ _7417_/CLK _7416_/D fanout586/X VGND VGND VPWR VPWR _7416_/Q sky130_fd_sc_hd__dfstp_2
X_4628_ _4747_/B _4795_/C _4772_/A VGND VGND VPWR VPWR _4628_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold530 _3485_/B VGND VGND VPWR VPWR _3557_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_7347_ _7539_/CLK hold87/X fanout577/X VGND VGND VPWR VPWR _7347_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4559_ _4086_/Y _5115_/A _4558_/X VGND VGND VPWR VPWR _5005_/A sky130_fd_sc_hd__a21o_4
Xhold541 _5949_/X VGND VGND VPWR VPWR _7536_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold552 _5950_/X VGND VGND VPWR VPWR _7537_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold563 hold563/A VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold574 hold574/A VGND VGND VPWR VPWR hold574/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7278_ _7278_/CLK _7278_/D fanout582/X VGND VGND VPWR VPWR _7278_/Q sky130_fd_sc_hd__dfrtp_1
Xhold585 hold585/A VGND VGND VPWR VPWR _7550_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold596 hold596/A VGND VGND VPWR VPWR hold596/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6475__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6229_ _7524_/Q _6112_/D _6119_/B _6136_/B _6121_/C VGND VGND VPWR VPWR _6229_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5640__C _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6490__A3 _6429_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1230 hold3052/X VGND VGND VPWR VPWR _7229_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6227__B1 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1241 _5939_/X VGND VGND VPWR VPWR _7527_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1252 hold3108/X VGND VGND VPWR VPWR hold3109/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1263 _5768_/X VGND VGND VPWR VPWR _7375_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1274 hold3139/X VGND VGND VPWR VPWR hold3140/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1285 _4540_/X VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 hold3160/X VGND VGND VPWR VPWR hold3161/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input87_A spimemio_flash_io1_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7471__SET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5505__A2 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4666__A_N _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3616__B _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output243_A _4152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3819__A2 _5902_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6481__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6805_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6821_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6218__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3930_ _3930_/A _5722_/A _4449_/B _5612_/B VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__and4_1
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3861_ _7264_/Q _5722_/A _5640_/B _5640_/C VGND VGND VPWR VPWR _3861_/X sky130_fd_sc_hd__and4_1
XFILLER_0_156_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5993__S hold37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5600_ _5600_/A0 _5647_/A0 _5602_/S VGND VGND VPWR VPWR _5600_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_183_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6580_ _7292_/Q _6422_/X _6457_/X _7476_/Q _6579_/X VGND VGND VPWR VPWR _6580_/X
+ sky130_fd_sc_hd__a221o_1
X_3792_ _3792_/A _3792_/B _3792_/C _3792_/D VGND VGND VPWR VPWR _3793_/D sky130_fd_sc_hd__nor4_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3755__A1 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5531_ _5531_/A _5531_/B _5531_/C _5531_/D VGND VGND VPWR VPWR _5532_/D sky130_fd_sc_hd__and4_1
XFILLER_0_14_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4910__B _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5462_ _4622_/Y _4654_/Y _4880_/Y _5461_/X _4854_/X VGND VGND VPWR VPWR _5462_/X
+ sky130_fd_sc_hd__o311a_2
X_7201_ _7201_/CLK _7201_/D _6839_/A VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4413_ _4413_/A0 _4412_/X _4423_/S VGND VGND VPWR VPWR _4413_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_111_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3526__B _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5393_ _5222_/A _4702_/Y _4755_/C _5453_/C _5100_/X VGND VGND VPWR VPWR _5393_/X
+ sky130_fd_sc_hd__o41a_1
X_7132_ _7176_/CLK _7132_/D fanout588/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_4
X_4344_ _5647_/A0 _4344_/A1 _4345_/S VGND VGND VPWR VPWR _4344_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6837__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7063_ _7189_/CLK _7063_/D fanout572/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfstp_2
X_4275_ _4275_/A0 _5852_/A0 _4276_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3542__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6014_ _7585_/Q _6017_/D _7586_/Q VGND VGND VPWR VPWR _6015_/C sky130_fd_sc_hd__a21o_1
XANTENNA__5680__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6209__B1 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_179_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6853__A _6871_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3691__B1 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout441_A _6424_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6916_ _7239_/CLK _6916_/D fanout566/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_65_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6847_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6847_/X sky130_fd_sc_hd__and2_1
XFILLER_0_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7522__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1389_A _7392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6778_ _7101_/Q _7102_/Q _6827_/A _7108_/Q _4115_/B VGND VGND VPWR VPWR _6778_/Y
+ sky130_fd_sc_hd__o41ai_1
XFILLER_0_107_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3746__A1 _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5729_ _5729_/A0 _5954_/A1 _5730_/S VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3746__B2 _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4820__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4312__S _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6145__C1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6696__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6160__A2 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold360 hold360/A VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold371 _4380_/X VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold382 hold382/A VGND VGND VPWR VPWR hold382/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6747__B _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold393 _5676_/X VGND VGND VPWR VPWR _7294_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6466__C _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input141_A wb_dat_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 hold2792/X VGND VGND VPWR VPWR hold2793/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 _4371_/X VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1082 hold2829/X VGND VGND VPWR VPWR hold2830/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 _4354_/X VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4283__A _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A1 _7648_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7263__RESET_B fanout569/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6687__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4618__B1_N _4795_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6151__A2 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4162__A1 _4164_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4060_ _7071_/Q _4001_/Y _4008_/Y _4059_/X VGND VGND VPWR VPWR _4067_/C sky130_fd_sc_hd__a31oi_4
XANTENNA__4177__B _4177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5662__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6206__A3 _6035_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5414__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_wire507_A wire508/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6611__B1 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4962_ _4962_/A _4962_/B VGND VGND VPWR VPWR _4962_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4624__C _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6701_ _6700_/X _6726_/A1 _6777_/S VGND VGND VPWR VPWR _6701_/X sky130_fd_sc_hd__mux2_1
X_3913_ _3913_/A _3913_/B _3913_/C _3913_/D VGND VGND VPWR VPWR _3921_/C sky130_fd_sc_hd__nor4_1
X_4893_ _5183_/A _5260_/D VGND VGND VPWR VPWR _4893_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6632_ _7558_/Q _6408_/A _6419_/D _7318_/Q VGND VGND VPWR VPWR _6632_/X sky130_fd_sc_hd__a22o_1
X_3844_ _7513_/Q _5920_/A _3838_/X _3840_/X _3843_/X VGND VGND VPWR VPWR _3844_/Y
+ sky130_fd_sc_hd__a2111oi_2
XANTENNA__3728__A1 _7141_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6563_ _7475_/Q _6424_/C _6441_/X _6425_/X _7339_/Q VGND VGND VPWR VPWR _6563_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3775_ _7402_/Q _5794_/A _3564_/X _7362_/Q _3774_/X VGND VGND VPWR VPWR _3782_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6390__A2 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3537__A _3537_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5514_ _5462_/X _5513_/X _5505_/X _5550_/C VGND VGND VPWR VPWR _5514_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_15_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6494_ _6494_/A _6494_/B _6494_/C _6494_/D VGND VGND VPWR VPWR _6495_/C sky130_fd_sc_hd__nor4_2
XANTENNA__6678__B1 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5445_ _5222_/A _5453_/C _5213_/B _5387_/D VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4153__A1 _7221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5376_ _4703_/Y _4844_/Y _5255_/X _4774_/Y VGND VGND VPWR VPWR _5384_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_2_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6693__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7115_ _7134_/CLK _7115_/D fanout589/X VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4327_ _5754_/A1 _4327_/A1 _4327_/S VGND VGND VPWR VPWR _4327_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout391_A hold2225/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_A hold43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7046_ _7151_/CLK _7046_/D fanout588/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfrtp_4
X_4258_ _4258_/A0 _5991_/A1 _4258_/S VGND VGND VPWR VPWR _4258_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5898__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4189_ _4189_/A0 hold166/X _7084_/Q VGND VGND VPWR VPWR _4189_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6602__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3719__A1 _7146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5184__A3 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6381__A2 _6072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1840_A _7521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1938_A _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire559 _4823_/C VGND VGND VPWR VPWR _5295_/D sky130_fd_sc_hd__buf_4
XFILLER_0_116_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6669__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6684__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5892__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold190 hold190/A VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4278__A _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4217__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A1 _7519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_185_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3560_ _7390_/Q _5776_/A _5704_/A _7326_/Q _3559_/X VGND VGND VPWR VPWR _3560_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6124__A2 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3491_ input28/X _3488_/X _3490_/X input19/X _3487_/X VGND VGND VPWR VPWR _3491_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_51_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5230_ _5213_/A _4929_/A _4943_/B _5102_/B _5091_/C VGND VGND VPWR VPWR _5231_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3209 _7619_/Q VGND VGND VPWR VPWR _6598_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5883__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5161_ _4748_/Y _5528_/A3 _4826_/Y _4814_/Y VGND VGND VPWR VPWR _5163_/C sky130_fd_sc_hd__a211o_1
XANTENNA__5722__D _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2508 _7227_/Q VGND VGND VPWR VPWR hold955/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2519 _7143_/Q VGND VGND VPWR VPWR hold694/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4112_ _6929_/Q _3409_/Y _4112_/B1 _6932_/Q VGND VGND VPWR VPWR _4112_/X sky130_fd_sc_hd__a22o_1
Xhold1807 hold412/X VGND VGND VPWR VPWR _5860_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5092_ _5260_/C _5091_/X _5067_/X _5090_/Y VGND VGND VPWR VPWR _5092_/Y sky130_fd_sc_hd__a211oi_1
Xhold1818 hold376/X VGND VGND VPWR VPWR _4525_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1829 _3511_/X VGND VGND VPWR VPWR hold1829/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4043_ _3399_/Y _4025_/A _3465_/Y _4040_/A VGND VGND VPWR VPWR _4043_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_79_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4127__S _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5994_ _5994_/A0 hold43/X hold37/X VGND VGND VPWR VPWR _5994_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4945_ _4945_/A _4960_/A VGND VGND VPWR VPWR _5248_/C sky130_fd_sc_hd__nor2_8
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2955_A _7331_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7664_ _7664_/A VGND VGND VPWR VPWR _7664_/X sky130_fd_sc_hd__clkbuf_2
X_4876_ _4861_/A _4861_/B _4974_/C _4974_/D VGND VGND VPWR VPWR _5216_/A sky130_fd_sc_hd__a22oi_4
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6615_ _7333_/Q _6423_/X _6606_/X _6610_/X _6614_/X VGND VGND VPWR VPWR _6615_/X
+ sky130_fd_sc_hd__a2111o_1
X_3827_ _7038_/Q _5803_/A _5623_/B _3824_/X _3826_/X VGND VGND VPWR VPWR _3828_/D
+ sky130_fd_sc_hd__a311o_1
X_7595_ _7610_/CLK _7595_/D fanout567/X VGND VGND VPWR VPWR _7595_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4370__B _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6363__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5020__C1 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5166__A3 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6546_ _7282_/Q _6431_/Y _6067_/A VGND VGND VPWR VPWR _6546_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5185__C _5185_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3758_ _7306_/Q _5686_/A _4467_/A _7130_/Q _3757_/X VGND VGND VPWR VPWR _3759_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6115__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6477_ _7512_/Q _6435_/X _6466_/X _7504_/Q VGND VGND VPWR VPWR _6477_/X sky130_fd_sc_hd__a22o_1
X_3689_ _7435_/Q _3525_/X _3651_/X _7050_/Q _3688_/X VGND VGND VPWR VPWR _3689_/X
+ sky130_fd_sc_hd__a221o_1
X_5428_ _5203_/B _5553_/A1 _5328_/X _5427_/X VGND VGND VPWR VPWR _5435_/D sky130_fd_sc_hd__a31o_1
Xoutput240 _7650_/X VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
Xoutput251 _4130_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
Xoutput262 _7226_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
XANTENNA__5874__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput273 _6916_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
X_5359_ _4915_/C _5346_/X _5228_/A VGND VGND VPWR VPWR _5573_/B sky130_fd_sc_hd__a21boi_1
Xoutput284 _7242_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xoutput295 _7244_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
XANTENNA__7375__SET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5626__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7029_ _7196_/CLK _7029_/D fanout590/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4826__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4545__B _5902_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input104_A wb_adr_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire345 _3844_/Y VGND VGND VPWR VPWR _3854_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__4365__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5617__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5093__A2 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6290__A1 _7187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4455__B _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6593__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4730_ _4984_/B _4802_/A _4730_/C VGND VGND VPWR VPWR _4730_/Y sky130_fd_sc_hd__nand3b_4
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4661_ _5058_/D _4888_/B _5282_/A _4805_/B VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__a31o_4
XANTENNA__6345__A2 _6332_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5002__C1 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6400_ _6751_/S _7613_/Q _6398_/X _6399_/X VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__a22o_1
X_3612_ _7240_/Q _3485_/X _5603_/B _3525_/X _7436_/Q VGND VGND VPWR VPWR _3612_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4356__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7380_ _7577_/CLK _7380_/D fanout583/X VGND VGND VPWR VPWR _7380_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3518__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4592_ _5115_/B _4591_/B _4675_/A _4675_/B _4586_/C VGND VGND VPWR VPWR _4592_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_71_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold904 hold904/A VGND VGND VPWR VPWR _7404_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6331_ _6330_/X _6331_/A1 _6777_/S VGND VGND VPWR VPWR _7611_/D sky130_fd_sc_hd__mux2_1
X_3543_ _5722_/A _5596_/B _5731_/B VGND VGND VPWR VPWR _3543_/X sky130_fd_sc_hd__and3_4
Xhold915 hold915/A VGND VGND VPWR VPWR hold915/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold926 _4531_/X VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold937 hold937/A VGND VGND VPWR VPWR hold937/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold948 hold948/A VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4410__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4108__A1 _6751_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold959 hold959/A VGND VGND VPWR VPWR hold959/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6262_ _7382_/Q _6089_/X _6093_/X _7366_/Q VGND VGND VPWR VPWR _6262_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_110_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3474_ _3474_/A _3576_/C VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__nor2_1
Xhold3006 _7012_/Q VGND VGND VPWR VPWR hold3006/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5213_ _5213_/A _5213_/B _5213_/C _5342_/B VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__and4_1
Xhold3017 hold738/X VGND VGND VPWR VPWR _5595_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3028 _7224_/Q VGND VGND VPWR VPWR hold3028/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3039 _5624_/X VGND VGND VPWR VPWR hold737/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6193_ hold96/A _6094_/A _6093_/X _6110_/X _7435_/Q VGND VGND VPWR VPWR _6193_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2305 _5665_/X VGND VGND VPWR VPWR hold924/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2316 _7499_/Q VGND VGND VPWR VPWR hold102/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2327 _7304_/Q VGND VGND VPWR VPWR hold588/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5144_ _4687_/Y _4713_/X _4821_/Y _4723_/Y _4716_/Y VGND VGND VPWR VPWR _5145_/C
+ sky130_fd_sc_hd__o32a_1
Xhold2338 _7280_/Q VGND VGND VPWR VPWR hold592/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1604 _5942_/X VGND VGND VPWR VPWR hold236/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2349 hold927/X VGND VGND VPWR VPWR _4507_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5608__A1 _5754_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1615 _5971_/X VGND VGND VPWR VPWR hold256/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1626 _4253_/X VGND VGND VPWR VPWR hold250/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_193_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1637 _7667_/A VGND VGND VPWR VPWR hold253/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3882__A3 _4212_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5075_ _4605_/Y _5451_/A1 _4709_/Y _5072_/Y _5074_/Y VGND VGND VPWR VPWR _5075_/Y
+ sky130_fd_sc_hd__o311ai_1
Xhold1648 hold273/X VGND VGND VPWR VPWR _5609_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1659 _6888_/Q VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3550__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4026_ _6904_/Q _4025_/B _6905_/Q VGND VGND VPWR VPWR _4026_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6033__A1 _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_176_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ _5986_/A1 _5977_/A1 _5982_/S VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_47_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4928_ _4933_/B _4928_/B VGND VGND VPWR VPWR _4930_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout619_A _4743_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6336__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4859_ _5248_/B _5453_/A _4859_/C VGND VGND VPWR VPWR _4949_/A sky130_fd_sc_hd__and3_1
XFILLER_0_16_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4347__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1469_A _3543_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5544__B1 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7578_ _7578_/CLK _7578_/D fanout604/X VGND VGND VPWR VPWR _7578_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6529_ _7578_/Q _6427_/X _6524_/X _6528_/X _6430_/X VGND VGND VPWR VPWR _6529_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4320__S _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5847__A1 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4259__C _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2850 hold2850/A VGND VGND VPWR VPWR hold2850/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_73_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6926_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2861 hold2861/A VGND VGND VPWR VPWR hold2861/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2872 _7046_/Q VGND VGND VPWR VPWR hold2872/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2883 hold2883/A VGND VGND VPWR VPWR hold2883/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5075__A2 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2894 _4552_/X VGND VGND VPWR VPWR hold2894/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_167_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6893__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4291__A _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7178_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_170_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4338__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output273_A _6916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_csclk _7267_/CLK VGND VGND VPWR VPWR _7560_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5838__A1 hold17/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__B1 _3846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4510__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5996__S hold37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5900_ _5999_/A1 _5900_/A1 _5901_/S VGND VGND VPWR VPWR _5900_/X sky130_fd_sc_hd__mux2_1
X_6880_ _4127_/A1 _6880_/D _6831_/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_2
X_5831_ _5831_/A0 _5993_/A1 _5838_/S VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6566__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5762_ _5987_/A1 _5762_/A1 _5766_/S VGND VGND VPWR VPWR _5762_/X sky130_fd_sc_hd__mux2_1
X_7501_ _7501_/CLK _7501_/D fanout581/X VGND VGND VPWR VPWR _7501_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3529__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4713_ _4733_/A _4733_/B _4801_/C _4712_/Y VGND VGND VPWR VPWR _4713_/X sky130_fd_sc_hd__a211o_2
XFILLER_0_17_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5693_ _5954_/A1 _5693_/A1 _5694_/S VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4329__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4644_ _4675_/A _4675_/B _4643_/C _4645_/D _5089_/B VGND VGND VPWR VPWR _4644_/Y
+ sky130_fd_sc_hd__a41oi_4
X_7432_ _7432_/CLK _7432_/D fanout593/X VGND VGND VPWR VPWR _7432_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_126_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4575_ _4887_/D _4887_/B _4879_/C _4805_/B VGND VGND VPWR VPWR _4984_/C sky130_fd_sc_hd__nand4_4
X_7363_ _7363_/CLK _7363_/D fanout575/X VGND VGND VPWR VPWR _7363_/Q sky130_fd_sc_hd__dfrtp_4
Xhold701 hold701/A VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold712 hold712/A VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_188_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3545__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold723 _4327_/X VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold734 hold734/A VGND VGND VPWR VPWR hold734/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6314_ _7062_/Q _6032_/Y _6313_/X _6144_/C VGND VGND VPWR VPWR _6314_/X sky130_fd_sc_hd__a211o_1
X_3526_ _3537_/A _5830_/C _5938_/C VGND VGND VPWR VPWR _3526_/X sky130_fd_sc_hd__and3_4
Xhold745 hold745/A VGND VGND VPWR VPWR hold745/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7294_ _7366_/CLK _7294_/D fanout579/X VGND VGND VPWR VPWR _7294_/Q sky130_fd_sc_hd__dfrtp_4
Xmax_cap464 _4426_/Y VGND VGND VPWR VPWR wire463/A sky130_fd_sc_hd__clkbuf_4
Xhold756 hold756/A VGND VGND VPWR VPWR _7277_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5829__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold767 hold767/A VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold778 _5909_/X VGND VGND VPWR VPWR _7501_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6245_ _7477_/Q _6032_/Y _6081_/X _7453_/Q _6244_/X VGND VGND VPWR VPWR _6245_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__7547__RESET_B fanout597/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold789 hold789/A VGND VGND VPWR VPWR hold789/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3457_ _4429_/B _3458_/A2 hold398/X VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__a21o_1
Xhold2102 _7443_/Q VGND VGND VPWR VPWR hold147/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2113 _7479_/Q VGND VGND VPWR VPWR hold474/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2124 _7507_/Q VGND VGND VPWR VPWR hold162/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6176_ _7370_/Q _6144_/C _6084_/X _6070_/X _7346_/Q VGND VGND VPWR VPWR _6176_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2135 _4251_/X VGND VGND VPWR VPWR hold539/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1401 hold4/X VGND VGND VPWR VPWR _4187_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2146 _7131_/Q VGND VGND VPWR VPWR hold2146/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2157 _4375_/X VGND VGND VPWR VPWR hold161/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1412 _7553_/Q VGND VGND VPWR VPWR hold1412/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5127_ _5127_/A _5295_/B _5138_/D VGND VGND VPWR VPWR _5164_/A sky130_fd_sc_hd__and3_1
Xhold2168 hold847/X VGND VGND VPWR VPWR _4210_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1423 hold193/X VGND VGND VPWR VPWR _5716_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout471_A _5863_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4376__A _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2179 hold885/X VGND VGND VPWR VPWR _5646_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1434 _7337_/Q VGND VGND VPWR VPWR hold201/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout569_A fanout587/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1445 hold11/X VGND VGND VPWR VPWR _3507_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1456 hold177/X VGND VGND VPWR VPWR _5649_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6254__B2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1467 _3504_/Y VGND VGND VPWR VPWR hold1467/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5058_ _4747_/B _5282_/A _5058_/C _5058_/D VGND VGND VPWR VPWR _5060_/B sky130_fd_sc_hd__and4b_1
Xhold1478 _5847_/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1489 _3458_/Y VGND VGND VPWR VPWR _3496_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _6910_/Q _6909_/Q _6908_/Q VGND VGND VPWR VPWR _4123_/B sky130_fd_sc_hd__and3_2
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6557__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6411__D1 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5765__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1586_A _3502_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5000__A _5138_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6309__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3791__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6190__B1 _6178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1920_A _7226_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input32_A mask_rev_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__buf_12
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2680 _7419_/Q VGND VGND VPWR VPWR hold767/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2691 _4550_/X VGND VGND VPWR VPWR hold764/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7431__SET_B fanout593/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__clkbuf_4
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1990 _7417_/Q VGND VGND VPWR VPWR hold549/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_187_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4225__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _3686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6720__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3534__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4360_ _4360_/A0 _5583_/A0 _4363_/S VGND VGND VPWR VPWR _4360_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4291_ _4302_/S _4291_/B VGND VGND VPWR VPWR _4291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6030_ _6106_/B _6019_/Y _6029_/X VGND VGND VPWR VPWR _7590_/D sky130_fd_sc_hd__a21o_1
XANTENNA__5287__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6484__B2 _7488_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3531__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6787__A2 _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4346__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6932_ _7601_/CLK _6932_/D fanout567/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6863_ _6873_/A _6869_/B VGND VGND VPWR VPWR _6863_/X sky130_fd_sc_hd__and2_1
XFILLER_0_190_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6539__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2770_A _6967_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5814_ _5814_/A0 _5967_/A1 _5820_/S VGND VGND VPWR VPWR _5814_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6794_ _6824_/B _6824_/C VGND VGND VPWR VPWR _6794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5745_ _5745_/A0 _5979_/A0 _5748_/S VGND VGND VPWR VPWR _5745_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5676_ _5955_/A1 _5676_/A1 _5676_/S VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7415_ _7415_/CLK _7415_/D fanout593/X VGND VGND VPWR VPWR _7415_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6172__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4627_ _4667_/A _5301_/A1 _4795_/C VGND VGND VPWR VPWR _4627_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_0_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6711__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold520 hold520/A VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4558_ _4825_/A _5071_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _4558_/X sky130_fd_sc_hd__and4_2
X_7346_ _7412_/CLK hold6/X fanout580/X VGND VGND VPWR VPWR _7346_/Q sky130_fd_sc_hd__dfrtp_4
Xhold531 hold531/A VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold542 hold542/A VGND VGND VPWR VPWR hold542/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold553 hold553/A VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold564 _5919_/X VGND VGND VPWR VPWR _7510_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold575 hold575/A VGND VGND VPWR VPWR _7237_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3509_ _7358_/Q _3564_/A _4212_/A _3508_/X _7558_/Q VGND VGND VPWR VPWR _3509_/X
+ sky130_fd_sc_hd__a32o_1
Xhold586 _7336_/Q VGND VGND VPWR VPWR hold586/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7277_ _7278_/CLK _7277_/D fanout580/X VGND VGND VPWR VPWR _7277_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4489_ _5647_/A0 _4489_/A1 _4490_/S VGND VGND VPWR VPWR _4489_/X sky130_fd_sc_hd__mux2_1
Xhold597 _4325_/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6475__A1 _7448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6475__B2 _7376_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6228_ _7388_/Q _6317_/C _6332_/B _6227_/X _6226_/X VGND VGND VPWR VPWR _6228_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4486__A0 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _7385_/Q _6112_/D _6106_/B _6144_/A _6112_/C VGND VGND VPWR VPWR _6159_/X
+ sky130_fd_sc_hd__a41o_1
Xhold1220 _4411_/X VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5640__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 hold3078/X VGND VGND VPWR VPWR hold3079/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1242 hold2939/X VGND VGND VPWR VPWR hold2940/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1253 hold3110/X VGND VGND VPWR VPWR _7551_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1264 hold3141/X VGND VGND VPWR VPWR hold3142/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1275 _4528_/X VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 hold3090/X VGND VGND VPWR VPWR hold3091/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1297 _4323_/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3764__A2 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4961__A1 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6163__B1 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3616__C _5731_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5910__A0 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6802_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6808_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6799_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6769__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5977__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4744__A _4879_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3860_ _7183_/Q _5875_/A _4449_/B _4551_/C VGND VGND VPWR VPWR _3860_/X sky130_fd_sc_hd__and4_1
XFILLER_0_86_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3791_ _7054_/Q _4509_/A _5619_/B _3788_/X _3790_/X VGND VGND VPWR VPWR _3792_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_183_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3755__A2 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5530_ _4956_/A _4834_/Y _5294_/C _5163_/C _5294_/B VGND VGND VPWR VPWR _5532_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4910__C _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5461_ _4965_/X _5461_/B VGND VGND VPWR VPWR _5461_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6154__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4412_ _4443_/A0 _5986_/A1 _4422_/S VGND VGND VPWR VPWR _4412_/X sky130_fd_sc_hd__mux2_1
X_7200_ _7201_/CLK _7200_/D _6839_/A VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5901__A0 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3526__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5392_ _5255_/X _4844_/Y _4703_/Y _4806_/Y _5563_/A1 VGND VGND VPWR VPWR _5394_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_151_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4343_ _5950_/A1 _4343_/A1 _4345_/S VGND VGND VPWR VPWR _4343_/X sky130_fd_sc_hd__mux2_1
X_7131_ _7395_/CLK _7131_/D fanout598/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7062_ _7190_/CLK hold44/X fanout573/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfrtp_4
X_4274_ _4274_/A0 _5914_/A1 _4276_/S VGND VGND VPWR VPWR _4274_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4468__A0 _5840_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6013_ _7585_/Q _7586_/Q _6017_/D VGND VGND VPWR VPWR _6015_/B sky130_fd_sc_hd__nand3_1
XANTENNA__3542__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6209__A1 _7459_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3691__A1 _7299_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_178_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_178_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5432__A2 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6915_ _6926_/CLK _6915_/D fanout566/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6846_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6846_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout434_A _6404_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6393__B1 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6777_ _6776_/X _6777_/A1 _6777_/S VGND VGND VPWR VPWR _7627_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_107_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3989_ input93/X _5722_/A _5938_/B _5612_/B _3930_/X VGND VGND VPWR VPWR _3989_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout601_A fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3746__A2 _4473_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5728_ _5728_/A0 _5863_/A0 _5730_/S VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4820__C _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5659_ _5947_/A _5659_/B _5902_/B VGND VGND VPWR VPWR _5667_/S sky130_fd_sc_hd__and3_4
XFILLER_0_143_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6696__A1 _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold350 hold350/A VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7329_ _7359_/CLK _7329_/D fanout576/X VGND VGND VPWR VPWR _7329_/Q sky130_fd_sc_hd__dfrtp_4
Xhold361 hold361/A VGND VGND VPWR VPWR _7402_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4829__A _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold372 hold372/A VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__A1 _7439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold383 _4392_/X VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6747__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold394 hold394/A VGND VGND VPWR VPWR hold394/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__B2 _7519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6466__D _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input134_A wb_dat_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _5985_/X VGND VGND VPWR VPWR _7568_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1061 hold2794/X VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1072 hold2864/X VGND VGND VPWR VPWR hold2865/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 hold2831/X VGND VGND VPWR VPWR _7439_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 hold2872/X VGND VGND VPWR VPWR hold2873/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__B1 _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4715__D_N _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3985__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6384__B1 _6144_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6439__A1 _7399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5139__A_N _5013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5414__A2 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4961_ _5180_/B _4953_/X _5252_/B _4959_/X VGND VGND VPWR VPWR _4962_/B sky130_fd_sc_hd__a211oi_1
X_6700_ _6649_/S _7623_/Q _6698_/Y _6699_/X VGND VGND VPWR VPWR _6700_/X sky130_fd_sc_hd__a22o_1
X_3912_ _7344_/Q _3545_/X _3562_/X _7296_/Q _3911_/X VGND VGND VPWR VPWR _3913_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_175_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3976__A2 _5640_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4892_ _4909_/C _4909_/D _4909_/A VGND VGND VPWR VPWR _4940_/D sky130_fd_sc_hd__and3_4
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6631_ _7582_/Q _6427_/X _6626_/X _6630_/X _6430_/X VGND VGND VPWR VPWR _6631_/Y
+ sky130_fd_sc_hd__a2111oi_4
XANTENNA__5178__A1 _5295_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3843_ _7481_/Q _3535_/X _3661_/X _7033_/Q _3842_/X VGND VGND VPWR VPWR _3843_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4921__B _4932_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4413__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3728__A2 _4491_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3774_ _7251_/Q _5640_/C _5623_/B _3648_/X _7039_/Q VGND VGND VPWR VPWR _3774_/X
+ sky130_fd_sc_hd__a32o_2
X_6562_ _7315_/Q _6419_/D _6451_/X _7483_/Q _6561_/X VGND VGND VPWR VPWR _6569_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3537__B _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5513_ _5113_/A _4953_/X _5366_/X _5512_/Y VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6127__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6493_ _7424_/Q _6463_/X _6468_/X _7408_/Q _6492_/X VGND VGND VPWR VPWR _6494_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6678__A1 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6678__B2 _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5444_ _5444_/A _5444_/B _5444_/C _5444_/D VGND VGND VPWR VPWR _5510_/B sky130_fd_sc_hd__and4_1
XANTENNA__5350__A1 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5375_ _4703_/Y _5255_/X _4844_/Y _4707_/Y VGND VGND VPWR VPWR _5473_/C sky130_fd_sc_hd__a31o_1
XANTENNA__3553__A hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7114_ _7134_/CLK _7114_/D fanout589/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfstp_4
X_4326_ _5647_/A0 _4326_/A1 _4327_/S VGND VGND VPWR VPWR _4326_/X sky130_fd_sc_hd__mux2_1
X_4257_ _4257_/A0 hold61/X _4258_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
X_7045_ _7134_/CLK _7045_/D _6833_/A VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout384_A _3492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4188_ _4188_/A0 _5852_/A0 _4190_/S VGND VGND VPWR VPWR _4188_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6063__C1 _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4815__C _5399_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5199__B _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1499_A _7444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3967__A2 _4509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6829_ wire463/A _6827_/Y _6828_/X _6826_/X VGND VGND VPWR VPWR _7646_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6366__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1666_A _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3719__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire538 _5072_/C VGND VGND VPWR VPWR _5282_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__6381__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6669__A1 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6669__B2 _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5341__A1 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold180 hold180/A VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold191 hold191/A VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4852__B1 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4294__A _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4741__B _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6372__A3 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_181_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3591__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3490_ _4449_/B _5612_/B _5612_/C VGND VGND VPWR VPWR _3490_/X sky130_fd_sc_hd__and3_4
XFILLER_0_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5160_ _5317_/A _5160_/B _5160_/C _5160_/D VGND VGND VPWR VPWR _5163_/B sky130_fd_sc_hd__nor4_1
Xhold2509 hold955/X VGND VGND VPWR VPWR _5594_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5999__S hold37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4111_ _7111_/Q _4084_/X _4425_/C VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__a21o_1
X_5091_ _5091_/A _5399_/A _5091_/C VGND VGND VPWR VPWR _5091_/X sky130_fd_sc_hd__and3_1
XFILLER_0_166_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1808 _5860_/X VGND VGND VPWR VPWR hold413/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1819 _4525_/X VGND VGND VPWR VPWR hold377/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4042_ _4042_/A _4042_/B VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4408__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6596__B1 _6775_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5993_ _5993_/A0 _5993_/A1 hold37/X VGND VGND VPWR VPWR _5993_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3949__A2 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4944_ _4944_/A _4944_/B _4944_/C VGND VGND VPWR VPWR _4949_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_164_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7663_ _7663_/A VGND VGND VPWR VPWR _7663_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6348__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4875_ _5328_/A _5328_/B _5203_/B VGND VGND VPWR VPWR _5038_/C sky130_fd_sc_hd__and3_4
XANTENNA__3548__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6614_ _7541_/Q _6427_/A _6574_/B _6747_/C _6613_/X VGND VGND VPWR VPWR _6614_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3826_ _7345_/Q _3545_/X _3649_/X _7068_/Q _3825_/X VGND VGND VPWR VPWR _3826_/X
+ sky130_fd_sc_hd__a221o_1
X_7594_ _7610_/CLK _7594_/D fanout568/X VGND VGND VPWR VPWR _7594_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6363__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6545_ _6529_/X _6545_/B _6545_/C VGND VGND VPWR VPWR _6545_/Y sky130_fd_sc_hd__nand3b_4
X_3757_ input55/X _5785_/B _5992_/C _3501_/X _7578_/Q VGND VGND VPWR VPWR _3757_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3582__B1 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6476_ _7520_/Q _6446_/X _6447_/X _7440_/Q _6475_/X VGND VGND VPWR VPWR _6476_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6115__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3688_ _7419_/Q _5875_/A _4212_/A _3687_/X VGND VGND VPWR VPWR _3688_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput230 _7667_/X VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
X_5427_ _4861_/X _5339_/C _5425_/X _5186_/X VGND VGND VPWR VPWR _5427_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5323__A1 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6520__B1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput241 _7651_/X VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
Xoutput252 _7671_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
XANTENNA_fanout599_A fanout602/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput263 _7227_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
Xoutput274 _6917_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
Xoutput285 _6927_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
X_5358_ _5213_/C _5038_/C _5342_/B _5357_/X VGND VGND VPWR VPWR _5361_/B sky130_fd_sc_hd__a31oi_1
XANTENNA_clkbuf_leaf_43_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3885__A1 _7392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput296 _7245_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
XANTENNA__3885__B2 _7504_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4309_ _4425_/B _4309_/B VGND VGND VPWR VPWR _4321_/S sky130_fd_sc_hd__nand2_8
X_5289_ _4858_/Y _4946_/Y _4622_/Y _4654_/Y VGND VGND VPWR VPWR _5461_/B sky130_fd_sc_hd__a211o_1
X_7028_ _7112_/CLK _7028_/D fanout589/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_0_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4617__B1_N _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6339__B1 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire346 _6733_/Y VGND VGND VPWR VPWR wire346/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_hold3164_A _7343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input62_A mgmt_gpio_in[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3876__A1 _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5078__B1 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6814__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6814__B2 _7109_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4736__B _4740_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout490 hold43/X VGND VGND VPWR VPWR _5967_/A1 sky130_fd_sc_hd__buf_12
XANTENNA__6290__A2 _6119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4455__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5848__A _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3800__A1 _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4660_ _5058_/D _4888_/B _5282_/A _4805_/B _4984_/B VGND VGND VPWR VPWR _4660_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_0_71_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6345__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3611_ input25/X _3488_/X _3490_/X input17/X _3610_/X VGND VGND VPWR VPWR _3623_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_114_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4591_ _5115_/B _4591_/B VGND VGND VPWR VPWR _4591_/Y sky130_fd_sc_hd__nor2_8
X_6330_ _6751_/S _6330_/A2 _6328_/X _6329_/X VGND VGND VPWR VPWR _6330_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_52_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3542_ _5640_/B _5612_/B _5612_/C VGND VGND VPWR VPWR _3542_/X sky130_fd_sc_hd__and3_4
XFILLER_0_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold905 hold905/A VGND VGND VPWR VPWR hold905/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold916 _4344_/X VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold927 hold927/A VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_101_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4108__A2 _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold938 hold938/A VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6261_ _6261_/A1 _4116_/X _6067_/X _6260_/X VGND VGND VPWR VPWR _7608_/D sky130_fd_sc_hd__o31a_1
XFILLER_0_12_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold949 hold949/A VGND VGND VPWR VPWR hold949/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6502__B1 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3473_ _4473_/A _4551_/A _5590_/A VGND VGND VPWR VPWR _3473_/X sky130_fd_sc_hd__and3_1
XANTENNA_hold2431_A _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3007 hold3007/A VGND VGND VPWR VPWR _4336_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5212_ _5068_/B _5387_/D _5248_/C _4904_/A VGND VGND VPWR VPWR _5349_/A sky130_fd_sc_hd__a31o_1
Xhold3018 _5595_/X VGND VGND VPWR VPWR hold739/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3029 hold3029/A VGND VGND VPWR VPWR _5591_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3867__A1 _7336_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6192_ _6192_/A1 _4116_/X _6067_/X _6191_/X VGND VGND VPWR VPWR _6192_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3867__B2 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2306 _7550_/Q VGND VGND VPWR VPWR hold584/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2317 hold102/X VGND VGND VPWR VPWR _5907_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5143_ _5143_/A _5143_/B _5143_/C VGND VGND VPWR VPWR _5145_/B sky130_fd_sc_hd__and3_1
Xhold2328 hold588/X VGND VGND VPWR VPWR _5688_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2339 hold592/X VGND VGND VPWR VPWR _5661_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1605 hold236/X VGND VGND VPWR VPWR _7530_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6805__A1 _7111_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1616 _7096_/Q VGND VGND VPWR VPWR hold259/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6805__B2 _7110_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1627 _7506_/Q VGND VGND VPWR VPWR hold247/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5074_ _5081_/A _5074_/B _5387_/C _5091_/A VGND VGND VPWR VPWR _5074_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1638 hold253/X VGND VGND VPWR VPWR _4435_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1649 _5609_/X VGND VGND VPWR VPWR hold274/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3550__B hold22/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4025_ _4025_/A _4025_/B VGND VGND VPWR VPWR _4025_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4138__S _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4292__A1 _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_189_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5758__A _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5976_ _5985_/A1 _5976_/A1 _5982_/S VGND VGND VPWR VPWR _5976_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_177_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6584__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4927_ _4927_/A _4927_/B _4927_/C VGND VGND VPWR VPWR _4930_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_176_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7646_ _7646_/CLK _7646_/D _6780_/B VGND VGND VPWR VPWR _7646_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4858_ _4856_/A _5072_/B _5058_/D VGND VGND VPWR VPWR _4858_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_117_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6336__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3809_ _7313_/Q _3521_/X _3804_/X _3806_/X _3808_/X VGND VGND VPWR VPWR _3809_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5544__A1 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7577_ _7577_/CLK hold9/X fanout584/X VGND VGND VPWR VPWR _7577_/Q sky130_fd_sc_hd__dfrtp_4
X_4789_ _5387_/C _4790_/C VGND VGND VPWR VPWR _4789_/Y sky130_fd_sc_hd__nand2_2
X_6528_ _7570_/Q _6424_/X _6526_/X _6527_/X VGND VGND VPWR VPWR _6528_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_160_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4844__A_N _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7176_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6459_ _7351_/Q _6459_/B _6459_/C VGND VGND VPWR VPWR _6459_/X sky130_fd_sc_hd__and3_1
XANTENNA__4259__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2840 hold2840/A VGND VGND VPWR VPWR hold2840/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2851 hold2851/A VGND VGND VPWR VPWR hold2851/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2862 _7000_/Q VGND VGND VPWR VPWR _4321_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2873 hold2873/A VGND VGND VPWR VPWR _4377_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2884 _7464_/Q VGND VGND VPWR VPWR hold2884/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5075__A3 _4709_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6272__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2895 _7630_/Q VGND VGND VPWR VPWR _6783_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7076__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6575__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_183_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3281_A _6895_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3546__B1 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output266_A _7229_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__A1 input45/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6263__A2 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4274__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5471__B1 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5830_ hold22/X _5866_/B _5830_/C _5992_/D VGND VGND VPWR VPWR _5838_/S sky130_fd_sc_hd__and4_4
XANTENNA_clkbuf_0_mgmt_gpio_in[4]_A mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_174_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5761_ _5896_/A0 _5761_/A1 _5766_/S VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7500_ _7572_/CLK _7500_/D fanout596/X VGND VGND VPWR VPWR _7500_/Q sky130_fd_sc_hd__dfrtp_4
X_4712_ _4753_/C _4767_/B VGND VGND VPWR VPWR _4712_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3785__B1 _3675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3529__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5692_ _5953_/A1 _5692_/A1 _5694_/S VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6318__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7431_ _7569_/CLK _7431_/D fanout593/X VGND VGND VPWR VPWR _7431_/Q sky130_fd_sc_hd__dfstp_2
X_4643_ _4675_/A _4675_/B _4643_/C _4645_/D VGND VGND VPWR VPWR _4643_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__5526__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4421__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7362_ _7366_/CLK _7362_/D fanout579/X VGND VGND VPWR VPWR _7362_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4574_ _5058_/D _4888_/B _5282_/A _4805_/B VGND VGND VPWR VPWR _4574_/X sky130_fd_sc_hd__and4_2
Xhold702 hold702/A VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold713 hold713/A VGND VGND VPWR VPWR _7424_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3545__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold724 hold724/A VGND VGND VPWR VPWR hold724/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6313_ _7193_/Q _6072_/B _6120_/B _6379_/B1 _7188_/Q VGND VGND VPWR VPWR _6313_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold735 _5934_/X VGND VGND VPWR VPWR _7523_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3525_ hold22/A _5875_/A _5830_/C VGND VGND VPWR VPWR _3525_/X sky130_fd_sc_hd__and3_4
Xhold746 _4308_/X VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7293_ _7366_/CLK _7293_/D fanout579/X VGND VGND VPWR VPWR _7293_/Q sky130_fd_sc_hd__dfrtp_4
Xmax_cap454 _4743_/Y VGND VGND VPWR VPWR _5061_/B sky130_fd_sc_hd__buf_4
Xhold757 hold757/A VGND VGND VPWR VPWR hold757/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold768 hold768/A VGND VGND VPWR VPWR _7419_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold779 hold779/A VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6244_ _7525_/Q _6112_/D _6119_/B _6136_/B _6144_/C VGND VGND VPWR VPWR _6244_/X
+ sky130_fd_sc_hd__a41o_1
X_3456_ _4429_/B _3456_/B VGND VGND VPWR VPWR _3456_/X sky130_fd_sc_hd__and2b_1
Xhold2103 hold147/X VGND VGND VPWR VPWR _5844_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2114 hold474/X VGND VGND VPWR VPWR _5885_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6175_ _7322_/Q _6082_/X _6099_/X _7354_/Q _6174_/X VGND VGND VPWR VPWR _6175_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2125 hold162/X VGND VGND VPWR VPWR _5916_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3561__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2136 _7121_/Q VGND VGND VPWR VPWR hold2136/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1402 _4187_/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2147 hold2147/A VGND VGND VPWR VPWR _4472_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2158 _7097_/Q VGND VGND VPWR VPWR hold169/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1413 hold1413/A VGND VGND VPWR VPWR _5968_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5126_ _4428_/B _4557_/Y _5125_/Y _4967_/Y VGND VGND VPWR VPWR _7202_/D sky130_fd_sc_hd__a22oi_1
Xhold1424 _5716_/X VGND VGND VPWR VPWR hold194/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2169 _4210_/X VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4376__B _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1435 hold201/X VGND VGND VPWR VPWR _5725_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6254__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1446 _3537_/A VGND VGND VPWR VPWR _3569_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1457 _5649_/X VGND VGND VPWR VPWR hold178/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1468 _3931_/D VGND VGND VPWR VPWR _5596_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_5057_ _5199_/C _5058_/C VGND VGND VPWR VPWR _5202_/C sky130_fd_sc_hd__nand2_1
Xhold1479 hold28/X VGND VGND VPWR VPWR _7446_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ _6910_/Q _6908_/Q VGND VGND VPWR VPWR _4008_/Y sky130_fd_sc_hd__nand2_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5959_ _5959_/A0 _5986_/A1 _5964_/S VGND VGND VPWR VPWR _5959_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5000__B _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6309__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7629_ _7630_/CLK _7629_/D VGND VGND VPWR VPWR _7629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3791__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6190__B2 _6189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input164_A wb_rstn_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6493__A2 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_117_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2670 hold765/X VGND VGND VPWR VPWR _4357_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input25_A mask_rev_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6245__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2681 hold767/X VGND VGND VPWR VPWR _5817_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2692 _7427_/Q VGND VGND VPWR VPWR hold761/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__buf_12
XANTENNA__4256__A1 _4256_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_187_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1980 hold452/X VGND VGND VPWR VPWR _4477_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1991 hold549/X VGND VGND VPWR VPWR _5815_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_86_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4559__A2 _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5756__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5220__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6705__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3646__A _4449_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4241__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6181__A1 _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _3706_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6720__A3 _6771_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4290_ _4425_/A _6780_/B VGND VGND VPWR VPWR _4302_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6484__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5692__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4495__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5800__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6931_ _7601_/CLK _6931_/D fanout567/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5995__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4924__B _4929_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4416__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6862_ _6865_/A _6869_/B VGND VGND VPWR VPWR _6862_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5813_ _5813_/A0 _5840_/A1 _5820_/S VGND VGND VPWR VPWR _5813_/X sky130_fd_sc_hd__mux2_1
X_6793_ _6824_/C _6793_/A2 _7107_/Q VGND VGND VPWR VPWR _6798_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5744_ _5744_/A0 _5987_/A1 _5748_/S VGND VGND VPWR VPWR _5744_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5675_ _5954_/A1 _5675_/A1 _5676_/S VGND VGND VPWR VPWR _5675_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_72_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7264_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3556__A hold36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7414_ _7478_/CLK _7414_/D fanout581/X VGND VGND VPWR VPWR _7414_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4151__S _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6172__A1 _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4626_ _4805_/B _4626_/B VGND VGND VPWR VPWR _4733_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_115_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6172__B2 _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold510 hold510/A VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5380__C1 _5451_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7345_ _7537_/CLK _7345_/D fanout577/X VGND VGND VPWR VPWR _7345_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold521 hold521/A VGND VGND VPWR VPWR _7231_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4557_ hold10/A _7107_/Q VGND VGND VPWR VPWR _4557_/Y sky130_fd_sc_hd__nor2_1
Xhold532 hold532/A VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_130_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold543 hold543/A VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold554 hold554/A VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold565 hold565/A VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3508_ _5590_/A _5992_/C _3931_/D VGND VGND VPWR VPWR _3508_/X sky130_fd_sc_hd__and3_4
X_7276_ _7577_/CLK _7276_/D fanout583/X VGND VGND VPWR VPWR _7276_/Q sky130_fd_sc_hd__dfrtp_1
X_4488_ _5950_/A1 _4488_/A1 _4490_/S VGND VGND VPWR VPWR _4488_/X sky130_fd_sc_hd__mux2_1
Xhold576 hold576/A VGND VGND VPWR VPWR hold576/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold587 hold587/A VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold598 hold598/A VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6227_ _7332_/Q _6136_/B _6116_/A _6084_/X _7372_/Q VGND VGND VPWR VPWR _6227_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6475__A2 _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3439_ _7330_/Q VGND VGND VPWR VPWR _3439_/Y sky130_fd_sc_hd__inv_2
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _7377_/Q _6089_/X _6379_/B1 _7393_/Q VGND VGND VPWR VPWR _6158_/X sky130_fd_sc_hd__a22o_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 hold1210/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 hold3059/X VGND VGND VPWR VPWR hold3060/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_10_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7070_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6227__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1232 _5777_/X VGND VGND VPWR VPWR _7383_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1243 _5621_/X VGND VGND VPWR VPWR _5622_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
X_5109_ _5118_/A _5453_/B _5113_/B VGND VGND VPWR VPWR _5111_/A sky130_fd_sc_hd__and3_1
XANTENNA__4238__A1 _5896_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1254 hold3064/X VGND VGND VPWR VPWR hold3065/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6089_ _6119_/A _6106_/B _6116_/C VGND VGND VPWR VPWR _6089_/X sky130_fd_sc_hd__and3_4
Xhold1265 hold3143/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_169_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1276 hold3113/X VGND VGND VPWR VPWR hold3114/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1287 hold3092/X VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 hold3102/X VGND VGND VPWR VPWR hold3103/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5986__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk _7267_/CLK VGND VGND VPWR VPWR _7566_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5738__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_192_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4410__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6163__A1 _7449_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6163__B2 _7505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3913__B _3913_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5674__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4477__A1 _5852_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4564_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6806_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3190 _7624_/Q VGND VGND VPWR VPWR _6726_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6811_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6803_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6218__A2 _6121_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7091__RESET_B fanout605/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4229__A1 hold61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6769__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_176_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4236__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5729__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4401__A1 _5714_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3790_ _7175_/Q _5866_/B _4521_/B _3789_/X VGND VGND VPWR VPWR _3790_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_82_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5460_ _4952_/B _5453_/C _5457_/Y _5459_/X VGND VGND VPWR VPWR _5460_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4411_ _4411_/A0 _4410_/X _4423_/S VGND VGND VPWR VPWR _4411_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5391_ _4601_/Y _4703_/Y _4744_/Y _4844_/Y _4798_/Y VGND VGND VPWR VPWR _5476_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_111_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7130_ _7395_/CLK _7130_/D fanout598/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfstp_2
X_4342_ hold43/X _4342_/A1 _4345_/S VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__mux2_1
X_7061_ _7268_/CLK _7061_/D _6873_/A VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfrtp_4
X_4273_ _4273_/A0 _5583_/A0 _4276_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
X_6012_ _4117_/Y _6010_/Y _6011_/X _6006_/A _6012_/B2 VGND VGND VPWR VPWR _7585_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3542__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

