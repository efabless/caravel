magic
tech sky130A
magscale 1 2
timestamp 1636991847
<< metal1 >>
rect 284662 995256 284668 995308
rect 284720 995296 284726 995308
rect 288986 995296 288992 995308
rect 284720 995268 288992 995296
rect 284720 995256 284726 995268
rect 288986 995256 288992 995268
rect 289044 995256 289050 995308
rect 538122 995256 538128 995308
rect 538180 995296 538186 995308
rect 539870 995296 539876 995308
rect 538180 995268 539876 995296
rect 538180 995256 538186 995268
rect 539870 995256 539876 995268
rect 539928 995256 539934 995308
rect 130286 995188 130292 995240
rect 130344 995228 130350 995240
rect 134610 995228 134616 995240
rect 130344 995200 134616 995228
rect 130344 995188 130350 995200
rect 134610 995188 134616 995200
rect 134668 995188 134674 995240
rect 526898 995188 526904 995240
rect 526956 995228 526962 995240
rect 531222 995228 531228 995240
rect 526956 995200 531228 995228
rect 526956 995188 526962 995200
rect 531222 995188 531228 995200
rect 531280 995188 531286 995240
rect 143258 995024 143264 995036
rect 142092 994996 143264 995024
rect 78858 994856 78864 994908
rect 78916 994896 78922 994908
rect 83182 994896 83188 994908
rect 78916 994868 83188 994896
rect 78916 994856 78922 994868
rect 83182 994856 83188 994868
rect 83240 994856 83246 994908
rect 83274 994856 83280 994908
rect 83332 994896 83338 994908
rect 133966 994896 133972 994908
rect 83332 994868 133972 994896
rect 83332 994856 83338 994868
rect 133966 994856 133972 994868
rect 134024 994896 134030 994908
rect 135162 994896 135168 994908
rect 134024 994868 135168 994896
rect 134024 994856 134030 994868
rect 135162 994856 135168 994868
rect 135220 994856 135226 994908
rect 135254 994856 135260 994908
rect 135312 994896 135318 994908
rect 142092 994896 142120 994996
rect 143258 994984 143264 994996
rect 143316 994984 143322 995036
rect 390756 994936 390968 994964
rect 135312 994868 142120 994896
rect 135312 994856 135318 994868
rect 186682 994856 186688 994908
rect 186740 994896 186746 994908
rect 194686 994896 194692 994908
rect 186740 994868 194692 994896
rect 186740 994856 186746 994868
rect 194686 994856 194692 994868
rect 194744 994856 194750 994908
rect 233694 994856 233700 994908
rect 233752 994896 233758 994908
rect 237466 994896 237472 994908
rect 233752 994868 237472 994896
rect 233752 994856 233758 994868
rect 237466 994856 237472 994868
rect 237524 994856 237530 994908
rect 288342 994896 288348 994908
rect 238726 994868 288348 994896
rect 79502 994788 79508 994840
rect 79560 994828 79566 994840
rect 130930 994828 130936 994840
rect 79560 994800 130936 994828
rect 79560 994788 79566 994800
rect 130930 994788 130936 994800
rect 130988 994828 130994 994840
rect 182358 994828 182364 994840
rect 130988 994800 182364 994828
rect 130988 994788 130994 994800
rect 182358 994788 182364 994800
rect 182416 994828 182422 994840
rect 183462 994828 183468 994840
rect 182416 994800 183468 994828
rect 182416 994788 182422 994800
rect 183462 994788 183468 994800
rect 183520 994788 183526 994840
rect 185394 994788 185400 994840
rect 185452 994828 185458 994840
rect 236730 994828 236736 994840
rect 185452 994800 236736 994828
rect 185452 994788 185458 994800
rect 236730 994788 236736 994800
rect 236788 994828 236794 994840
rect 238726 994828 238754 994868
rect 288342 994856 288348 994868
rect 288400 994856 288406 994908
rect 289630 994856 289636 994908
rect 289688 994896 289694 994908
rect 297634 994896 297640 994908
rect 289688 994868 297640 994896
rect 289688 994856 289694 994868
rect 297634 994856 297640 994868
rect 297692 994856 297698 994908
rect 295794 994828 295800 994840
rect 236788 994800 238754 994828
rect 248386 994800 295800 994828
rect 236788 994788 236794 994800
rect 89990 994720 89996 994772
rect 90048 994760 90054 994772
rect 141418 994760 141424 994772
rect 90048 994732 141424 994760
rect 90048 994720 90054 994732
rect 141418 994720 141424 994732
rect 141476 994760 141482 994772
rect 192846 994760 192852 994772
rect 141476 994732 192852 994760
rect 141476 994720 141482 994732
rect 192846 994720 192852 994732
rect 192904 994760 192910 994772
rect 244182 994760 244188 994772
rect 192904 994732 244188 994760
rect 192904 994720 192910 994732
rect 244182 994720 244188 994732
rect 244240 994760 244246 994772
rect 248386 994760 248414 994800
rect 295794 994788 295800 994800
rect 295852 994828 295858 994840
rect 390756 994828 390784 994936
rect 390940 994896 390968 994936
rect 390940 994868 391060 994896
rect 295852 994800 390784 994828
rect 391032 994828 391060 994868
rect 391474 994856 391480 994908
rect 391532 994896 391538 994908
rect 399478 994896 399484 994908
rect 391532 994868 399484 994896
rect 391532 994856 391538 994868
rect 399478 994856 399484 994868
rect 399536 994856 399542 994908
rect 480438 994856 480444 994908
rect 480496 994896 480502 994908
rect 488442 994896 488448 994908
rect 480496 994868 488448 994896
rect 480496 994856 480502 994868
rect 488442 994856 488448 994868
rect 488500 994856 488506 994908
rect 531866 994856 531872 994908
rect 531924 994896 531930 994908
rect 538122 994896 538128 994908
rect 531924 994868 538128 994896
rect 531924 994856 531930 994868
rect 538122 994856 538128 994868
rect 538180 994856 538186 994908
rect 633618 994856 633624 994908
rect 633676 994896 633682 994908
rect 641622 994896 641628 994908
rect 633676 994868 641628 994896
rect 633676 994856 633682 994868
rect 641622 994856 641628 994868
rect 641680 994856 641686 994908
rect 397638 994828 397644 994840
rect 391032 994800 397644 994828
rect 295852 994788 295858 994800
rect 397638 994788 397644 994800
rect 397696 994828 397702 994840
rect 486602 994828 486608 994840
rect 397696 994800 486608 994828
rect 397696 994788 397702 994800
rect 486602 994788 486608 994800
rect 486660 994828 486666 994840
rect 538030 994828 538036 994840
rect 486660 994800 538036 994828
rect 486660 994788 486666 994800
rect 538030 994788 538036 994800
rect 538088 994828 538094 994840
rect 639782 994828 639788 994840
rect 538088 994800 639788 994828
rect 538088 994788 538094 994800
rect 639782 994788 639788 994800
rect 639840 994788 639846 994840
rect 244240 994732 248414 994760
rect 244240 994720 244246 994732
rect 288618 994720 288624 994772
rect 288676 994760 288682 994772
rect 288986 994760 288992 994772
rect 288676 994732 288992 994760
rect 288676 994720 288682 994732
rect 288986 994720 288992 994732
rect 289044 994760 289050 994772
rect 386506 994760 386512 994772
rect 289044 994732 386512 994760
rect 289044 994720 289050 994732
rect 386506 994720 386512 994732
rect 386564 994760 386570 994772
rect 390646 994760 390652 994772
rect 386564 994732 390652 994760
rect 386564 994720 386570 994732
rect 390646 994720 390652 994732
rect 390704 994720 390710 994772
rect 476114 994760 476120 994772
rect 390848 994732 476120 994760
rect 83182 994652 83188 994704
rect 83240 994692 83246 994704
rect 130286 994692 130292 994704
rect 83240 994664 130292 994692
rect 83240 994652 83246 994664
rect 130286 994652 130292 994664
rect 130344 994692 130350 994704
rect 181714 994692 181720 994704
rect 130344 994664 181720 994692
rect 130344 994652 130350 994664
rect 181714 994652 181720 994664
rect 181772 994692 181778 994704
rect 186038 994692 186044 994704
rect 181772 994664 186044 994692
rect 181772 994652 181778 994664
rect 186038 994652 186044 994664
rect 186096 994692 186102 994704
rect 233050 994692 233056 994704
rect 186096 994664 233056 994692
rect 186096 994652 186102 994664
rect 233050 994652 233056 994664
rect 233108 994692 233114 994704
rect 237374 994692 237380 994704
rect 233108 994664 237380 994692
rect 233108 994652 233114 994664
rect 237374 994652 237380 994664
rect 237432 994652 237438 994704
rect 237466 994652 237472 994704
rect 237524 994692 237530 994704
rect 285306 994692 285312 994704
rect 237524 994664 285312 994692
rect 237524 994652 237530 994664
rect 285306 994652 285312 994664
rect 285364 994692 285370 994704
rect 333238 994692 333244 994704
rect 285364 994664 333244 994692
rect 285364 994652 285370 994664
rect 333238 994652 333244 994664
rect 333296 994692 333302 994704
rect 387150 994692 387156 994704
rect 333296 994664 387156 994692
rect 333296 994652 333302 994664
rect 387150 994652 387156 994664
rect 387208 994692 387214 994704
rect 390848 994692 390876 994732
rect 476114 994720 476120 994732
rect 476172 994760 476178 994772
rect 527542 994760 527548 994772
rect 476172 994732 527548 994760
rect 476172 994720 476178 994732
rect 527542 994720 527548 994732
rect 527600 994760 527606 994772
rect 528278 994760 528284 994772
rect 527600 994732 528284 994760
rect 527600 994720 527606 994732
rect 528278 994720 528284 994732
rect 528336 994720 528342 994772
rect 531222 994720 531228 994772
rect 531280 994760 531286 994772
rect 632330 994760 632336 994772
rect 531280 994732 632336 994760
rect 531280 994720 531286 994732
rect 632330 994720 632336 994732
rect 632388 994720 632394 994772
rect 387208 994664 390876 994692
rect 387208 994652 387214 994664
rect 390922 994652 390928 994704
rect 390980 994692 390986 994704
rect 475470 994692 475476 994704
rect 390980 994664 475476 994692
rect 390980 994652 390986 994664
rect 475470 994652 475476 994664
rect 475528 994692 475534 994704
rect 479794 994692 479800 994704
rect 475528 994664 479800 994692
rect 475528 994652 475534 994664
rect 479794 994652 479800 994664
rect 479852 994692 479858 994704
rect 526898 994692 526904 994704
rect 479852 994664 526904 994692
rect 479852 994652 479858 994664
rect 526898 994652 526904 994664
rect 526956 994692 526962 994704
rect 628650 994692 628656 994704
rect 526956 994664 628656 994692
rect 526956 994652 526962 994664
rect 628650 994652 628656 994664
rect 628708 994692 628714 994704
rect 632974 994692 632980 994704
rect 628708 994664 632980 994692
rect 628708 994652 628714 994664
rect 632974 994652 632980 994664
rect 633032 994652 633038 994704
rect 83826 994584 83832 994636
rect 83884 994624 83890 994636
rect 91830 994624 91836 994636
rect 83884 994596 91836 994624
rect 83884 994584 83890 994596
rect 91830 994584 91836 994596
rect 91888 994584 91894 994636
rect 183462 994584 183468 994636
rect 183520 994624 183526 994636
rect 233694 994624 233700 994636
rect 183520 994596 233700 994624
rect 183520 994584 183526 994596
rect 233694 994584 233700 994596
rect 233752 994584 233758 994636
rect 237392 994624 237420 994652
rect 288618 994624 288624 994636
rect 237392 994596 288624 994624
rect 288618 994584 288624 994596
rect 288676 994584 288682 994636
rect 390186 994624 390192 994636
rect 296686 994596 390192 994624
rect 135162 994516 135168 994568
rect 135220 994556 135226 994568
rect 185394 994556 185400 994568
rect 135220 994528 185400 994556
rect 135220 994516 135226 994528
rect 185394 994516 185400 994528
rect 185452 994516 185458 994568
rect 238018 994516 238024 994568
rect 238076 994556 238082 994568
rect 246022 994556 246028 994568
rect 238076 994528 246028 994556
rect 238076 994516 238082 994528
rect 246022 994516 246028 994528
rect 246080 994516 246086 994568
rect 288342 994516 288348 994568
rect 288400 994556 288406 994568
rect 296686 994556 296714 994596
rect 390186 994584 390192 994596
rect 390244 994624 390250 994636
rect 479150 994624 479156 994636
rect 390244 994596 479156 994624
rect 390244 994584 390250 994596
rect 479150 994584 479156 994596
rect 479208 994624 479214 994636
rect 479208 994596 480254 994624
rect 479208 994584 479214 994596
rect 288400 994528 296714 994556
rect 480226 994556 480254 994596
rect 528278 994584 528284 994636
rect 528336 994624 528342 994636
rect 629294 994624 629300 994636
rect 528336 994596 629300 994624
rect 528336 994584 528342 994596
rect 629294 994584 629300 994596
rect 629352 994584 629358 994636
rect 530578 994556 530584 994568
rect 480226 994528 530584 994556
rect 288400 994516 288406 994528
rect 530578 994516 530584 994528
rect 530636 994556 530642 994568
rect 531222 994556 531228 994568
rect 530636 994528 531228 994556
rect 530636 994516 530642 994528
rect 531222 994516 531228 994528
rect 531280 994516 531286 994568
rect 43622 994380 43628 994432
rect 43680 994420 43686 994432
rect 78858 994420 78864 994432
rect 43680 994392 78864 994420
rect 43680 994380 43686 994392
rect 78858 994380 78864 994392
rect 78916 994380 78922 994432
rect 639782 994380 639788 994432
rect 639840 994420 639846 994432
rect 674190 994420 674196 994432
rect 639840 994392 674196 994420
rect 639840 994380 639846 994392
rect 674190 994380 674196 994392
rect 674248 994380 674254 994432
rect 43438 994312 43444 994364
rect 43496 994352 43502 994364
rect 79502 994352 79508 994364
rect 43496 994324 79508 994352
rect 43496 994312 43502 994324
rect 79502 994312 79508 994324
rect 79560 994312 79566 994364
rect 632330 994312 632336 994364
rect 632388 994352 632394 994364
rect 674282 994352 674288 994364
rect 632388 994324 674288 994352
rect 632388 994312 632394 994324
rect 674282 994312 674288 994324
rect 674340 994312 674346 994364
rect 43530 994244 43536 994296
rect 43588 994284 43594 994296
rect 82538 994284 82544 994296
rect 43588 994256 82544 994284
rect 43588 994244 43594 994256
rect 82538 994244 82544 994256
rect 82596 994284 82602 994296
rect 83274 994284 83280 994296
rect 82596 994256 83280 994284
rect 82596 994244 82602 994256
rect 83274 994244 83280 994256
rect 83332 994244 83338 994296
rect 632974 994244 632980 994296
rect 633032 994284 633038 994296
rect 674374 994284 674380 994296
rect 633032 994256 674380 994284
rect 633032 994244 633038 994256
rect 674374 994244 674380 994256
rect 674432 994244 674438 994296
rect 42334 994176 42340 994228
rect 42392 994216 42398 994228
rect 89990 994216 89996 994228
rect 42392 994188 89996 994216
rect 42392 994176 42398 994188
rect 89990 994176 89996 994188
rect 90048 994176 90054 994228
rect 629294 994176 629300 994228
rect 629352 994216 629358 994228
rect 675110 994216 675116 994228
rect 629352 994188 675116 994216
rect 629352 994176 629358 994188
rect 675110 994176 675116 994188
rect 675168 994176 675174 994228
rect 580534 994088 580540 994140
rect 580592 994128 580598 994140
rect 674098 994128 674104 994140
rect 580592 994100 674104 994128
rect 580592 994088 580598 994100
rect 674098 994088 674104 994100
rect 674156 994088 674162 994140
rect 41782 967920 41788 967972
rect 41840 967960 41846 967972
rect 42426 967960 42432 967972
rect 41840 967932 42432 967960
rect 41840 967920 41846 967932
rect 42426 967920 42432 967932
rect 42484 967920 42490 967972
rect 674374 967376 674380 967428
rect 674432 967416 674438 967428
rect 675202 967416 675208 967428
rect 674432 967388 675208 967416
rect 674432 967376 674438 967388
rect 675202 967376 675208 967388
rect 675260 967376 675266 967428
rect 675202 965268 675208 965320
rect 675260 965308 675266 965320
rect 675386 965308 675392 965320
rect 675260 965280 675392 965308
rect 675260 965268 675266 965280
rect 675386 965268 675392 965280
rect 675444 965268 675450 965320
rect 674282 964112 674288 964164
rect 674340 964152 674346 964164
rect 675294 964152 675300 964164
rect 674340 964124 675300 964152
rect 674340 964112 674346 964124
rect 675294 964112 675300 964124
rect 675352 964112 675358 964164
rect 41782 961324 41788 961376
rect 41840 961364 41846 961376
rect 42334 961364 42340 961376
rect 41840 961336 42340 961364
rect 41840 961324 41846 961336
rect 42334 961324 42340 961336
rect 42392 961364 42398 961376
rect 43622 961364 43628 961376
rect 42392 961336 43628 961364
rect 42392 961324 42398 961336
rect 43622 961324 43628 961336
rect 43680 961324 43686 961376
rect 674926 960644 674932 960696
rect 674984 960684 674990 960696
rect 675386 960684 675392 960696
rect 674984 960656 675392 960684
rect 674984 960644 674990 960656
rect 675386 960644 675392 960656
rect 675444 960644 675450 960696
rect 675202 960168 675208 960220
rect 675260 960168 675266 960220
rect 675220 960016 675248 960168
rect 675202 959964 675208 960016
rect 675260 959964 675266 960016
rect 42242 959012 42248 959064
rect 42300 959052 42306 959064
rect 42610 959052 42616 959064
rect 42300 959024 42616 959052
rect 42300 959012 42306 959024
rect 42610 959012 42616 959024
rect 42668 959052 42674 959064
rect 43530 959052 43536 959064
rect 42668 959024 43536 959052
rect 42668 959012 42674 959024
rect 43530 959012 43536 959024
rect 43588 959012 43594 959064
rect 41782 957652 41788 957704
rect 41840 957692 41846 957704
rect 43438 957692 43444 957704
rect 41840 957664 43444 957692
rect 41840 957652 41846 957664
rect 43438 957652 43444 957664
rect 43496 957652 43502 957704
rect 42426 957448 42432 957500
rect 42484 957448 42490 957500
rect 42444 957296 42472 957448
rect 42426 957244 42432 957296
rect 42484 957244 42490 957296
rect 674190 953300 674196 953352
rect 674248 953340 674254 953352
rect 675110 953340 675116 953352
rect 674248 953312 675116 953340
rect 674248 953300 674254 953312
rect 675110 953300 675116 953312
rect 675168 953340 675174 953352
rect 675570 953340 675576 953352
rect 675168 953312 675576 953340
rect 675168 953300 675174 953312
rect 675570 953300 675576 953312
rect 675628 953300 675634 953352
rect 675018 875780 675024 875832
rect 675076 875820 675082 875832
rect 675386 875820 675392 875832
rect 675076 875792 675392 875820
rect 675076 875780 675082 875792
rect 675386 875780 675392 875792
rect 675444 875780 675450 875832
rect 674834 874488 674840 874540
rect 674892 874528 674898 874540
rect 675202 874528 675208 874540
rect 674892 874500 675208 874528
rect 674892 874488 674898 874500
rect 675202 874488 675208 874500
rect 675260 874528 675266 874540
rect 675386 874528 675392 874540
rect 675260 874500 675392 874528
rect 675260 874488 675266 874500
rect 675386 874488 675392 874500
rect 675444 874488 675450 874540
rect 675018 871632 675024 871684
rect 675076 871672 675082 871684
rect 675386 871672 675392 871684
rect 675076 871644 675392 871672
rect 675076 871632 675082 871644
rect 675386 871632 675392 871644
rect 675444 871632 675450 871684
rect 674926 864084 674932 864136
rect 674984 864124 674990 864136
rect 675110 864124 675116 864136
rect 674984 864096 675116 864124
rect 674984 864084 674990 864096
rect 675110 864084 675116 864096
rect 675168 864124 675174 864136
rect 675386 864124 675392 864136
rect 675168 864096 675392 864124
rect 675168 864084 675174 864096
rect 675386 864084 675392 864096
rect 675444 864084 675450 864136
rect 675294 818320 675300 818372
rect 675352 818360 675358 818372
rect 677502 818360 677508 818372
rect 675352 818332 677508 818360
rect 675352 818320 675358 818332
rect 677502 818320 677508 818332
rect 677560 818320 677566 818372
rect 41782 799552 41788 799604
rect 41840 799592 41846 799604
rect 42334 799592 42340 799604
rect 41840 799564 42340 799592
rect 41840 799552 41846 799564
rect 42334 799552 42340 799564
rect 42392 799552 42398 799604
rect 41782 797716 41788 797768
rect 41840 797756 41846 797768
rect 42426 797756 42432 797768
rect 41840 797728 42432 797756
rect 41840 797716 41846 797728
rect 42426 797716 42432 797728
rect 42484 797756 42490 797768
rect 42610 797756 42616 797768
rect 42484 797728 42616 797756
rect 42484 797716 42490 797728
rect 42610 797716 42616 797728
rect 42668 797716 42674 797768
rect 41782 792548 41788 792600
rect 41840 792588 41846 792600
rect 42334 792588 42340 792600
rect 41840 792560 42340 792588
rect 41840 792548 41846 792560
rect 42334 792548 42340 792560
rect 42392 792548 42398 792600
rect 41782 791936 41788 791988
rect 41840 791976 41846 791988
rect 42518 791976 42524 791988
rect 41840 791948 42524 791976
rect 41840 791936 41846 791948
rect 42518 791936 42524 791948
rect 42576 791936 42582 791988
rect 41782 787244 41788 787296
rect 41840 787284 41846 787296
rect 42518 787284 42524 787296
rect 41840 787256 42524 787284
rect 41840 787244 41846 787256
rect 42518 787244 42524 787256
rect 42576 787244 42582 787296
rect 41782 786632 41788 786684
rect 41840 786672 41846 786684
rect 42334 786672 42340 786684
rect 41840 786644 42340 786672
rect 41840 786632 41846 786644
rect 42334 786632 42340 786644
rect 42392 786632 42398 786684
rect 675202 786564 675208 786616
rect 675260 786604 675266 786616
rect 675386 786604 675392 786616
rect 675260 786576 675392 786604
rect 675260 786564 675266 786576
rect 675386 786564 675392 786576
rect 675444 786564 675450 786616
rect 674834 785272 674840 785324
rect 674892 785312 674898 785324
rect 675386 785312 675392 785324
rect 674892 785284 675392 785312
rect 674892 785272 674898 785284
rect 675386 785272 675392 785284
rect 675444 785272 675450 785324
rect 675018 783232 675024 783284
rect 675076 783272 675082 783284
rect 675386 783272 675392 783284
rect 675076 783244 675392 783272
rect 675076 783232 675082 783244
rect 675386 783232 675392 783244
rect 675444 783232 675450 783284
rect 675202 782688 675208 782740
rect 675260 782728 675266 782740
rect 675386 782728 675392 782740
rect 675260 782700 675392 782728
rect 675260 782688 675266 782700
rect 675386 782688 675392 782700
rect 675444 782688 675450 782740
rect 675202 780988 675208 781040
rect 675260 781028 675266 781040
rect 675386 781028 675392 781040
rect 675260 781000 675392 781028
rect 675260 780988 675266 781000
rect 675386 780988 675392 781000
rect 675444 780988 675450 781040
rect 674926 775004 674932 775056
rect 674984 775044 674990 775056
rect 675386 775044 675392 775056
rect 674984 775016 675392 775044
rect 674984 775004 674990 775016
rect 675386 775004 675392 775016
rect 675444 775004 675450 775056
rect 675202 773984 675208 774036
rect 675260 774024 675266 774036
rect 675386 774024 675392 774036
rect 675260 773996 675392 774024
rect 675260 773984 675266 773996
rect 675386 773984 675392 773996
rect 675444 773984 675450 774036
rect 41782 756372 41788 756424
rect 41840 756412 41846 756424
rect 42702 756412 42708 756424
rect 41840 756384 42708 756412
rect 41840 756372 41846 756384
rect 42702 756372 42708 756384
rect 42760 756372 42766 756424
rect 41782 755352 41788 755404
rect 41840 755392 41846 755404
rect 42426 755392 42432 755404
rect 41840 755364 42432 755392
rect 41840 755352 41846 755364
rect 42426 755352 42432 755364
rect 42484 755392 42490 755404
rect 42610 755392 42616 755404
rect 42484 755364 42616 755392
rect 42484 755352 42490 755364
rect 42610 755352 42616 755364
rect 42668 755352 42674 755404
rect 41782 749368 41788 749420
rect 41840 749408 41846 749420
rect 42702 749408 42708 749420
rect 41840 749380 42708 749408
rect 41840 749368 41846 749380
rect 42702 749368 42708 749380
rect 42760 749368 42766 749420
rect 41782 747668 41788 747720
rect 41840 747708 41846 747720
rect 42334 747708 42340 747720
rect 41840 747680 42340 747708
rect 41840 747668 41846 747680
rect 42334 747668 42340 747680
rect 42392 747668 42398 747720
rect 41782 745084 41788 745136
rect 41840 745124 41846 745136
rect 42518 745124 42524 745136
rect 41840 745096 42524 745124
rect 41840 745084 41846 745096
rect 42518 745084 42524 745096
rect 42576 745084 42582 745136
rect 41782 743792 41788 743844
rect 41840 743832 41846 743844
rect 42334 743832 42340 743844
rect 41840 743804 42340 743832
rect 41840 743792 41846 743804
rect 42334 743792 42340 743804
rect 42392 743792 42398 743844
rect 675110 741004 675116 741056
rect 675168 741044 675174 741056
rect 675570 741044 675576 741056
rect 675168 741016 675576 741044
rect 675168 741004 675174 741016
rect 675570 741004 675576 741016
rect 675628 741004 675634 741056
rect 674834 740324 674840 740376
rect 674892 740364 674898 740376
rect 675202 740364 675208 740376
rect 674892 740336 675208 740364
rect 674892 740324 674898 740336
rect 675202 740324 675208 740336
rect 675260 740364 675266 740376
rect 675386 740364 675392 740376
rect 675260 740336 675392 740364
rect 675260 740324 675266 740336
rect 675386 740324 675392 740336
rect 675444 740324 675450 740376
rect 675018 737264 675024 737316
rect 675076 737304 675082 737316
rect 675386 737304 675392 737316
rect 675076 737276 675392 737304
rect 675076 737264 675082 737276
rect 675386 737264 675392 737276
rect 675444 737264 675450 737316
rect 675110 736992 675116 737044
rect 675168 737032 675174 737044
rect 675386 737032 675392 737044
rect 675168 737004 675392 737032
rect 675168 736992 675174 737004
rect 675386 736992 675392 737004
rect 675444 736992 675450 737044
rect 674834 735972 674840 736024
rect 674892 736012 674898 736024
rect 675386 736012 675392 736024
rect 674892 735984 675392 736012
rect 674892 735972 674898 735984
rect 675386 735972 675392 735984
rect 675444 735972 675450 736024
rect 674926 729920 674932 729972
rect 674984 729960 674990 729972
rect 675386 729960 675392 729972
rect 674984 729932 675392 729960
rect 674984 729920 674990 729932
rect 675386 729920 675392 729932
rect 675444 729920 675450 729972
rect 674834 729036 674840 729088
rect 674892 729076 674898 729088
rect 675386 729076 675392 729088
rect 674892 729048 675392 729076
rect 674892 729036 674898 729048
rect 675386 729036 675392 729048
rect 675444 729036 675450 729088
rect 675294 726656 675300 726708
rect 675352 726656 675358 726708
rect 675312 726504 675340 726656
rect 674926 726452 674932 726504
rect 674984 726492 674990 726504
rect 675202 726492 675208 726504
rect 674984 726464 675208 726492
rect 674984 726452 674990 726464
rect 675202 726452 675208 726464
rect 675260 726452 675266 726504
rect 675294 726452 675300 726504
rect 675352 726452 675358 726504
rect 41782 713124 41788 713176
rect 41840 713164 41846 713176
rect 42426 713164 42432 713176
rect 41840 713136 42432 713164
rect 41840 713124 41846 713136
rect 42426 713124 42432 713136
rect 42484 713124 42490 713176
rect 41782 711696 41788 711748
rect 41840 711736 41846 711748
rect 42610 711736 42616 711748
rect 41840 711708 42616 711736
rect 41840 711696 41846 711708
rect 42610 711696 42616 711708
rect 42668 711696 42674 711748
rect 41782 706188 41788 706240
rect 41840 706228 41846 706240
rect 42426 706228 42432 706240
rect 41840 706200 42432 706228
rect 41840 706188 41846 706200
rect 42426 706188 42432 706200
rect 42484 706188 42490 706240
rect 42334 705780 42340 705832
rect 42392 705780 42398 705832
rect 42352 705560 42380 705780
rect 41782 705508 41788 705560
rect 41840 705548 41846 705560
rect 42334 705548 42340 705560
rect 41840 705520 42340 705548
rect 41840 705508 41846 705520
rect 42334 705508 42340 705520
rect 42392 705508 42398 705560
rect 42242 705168 42248 705220
rect 42300 705168 42306 705220
rect 41782 704896 41788 704948
rect 41840 704936 41846 704948
rect 42260 704936 42288 705168
rect 42518 704936 42524 704948
rect 41840 704908 42524 704936
rect 41840 704896 41846 704908
rect 42518 704896 42524 704908
rect 42576 704896 42582 704948
rect 41782 700816 41788 700868
rect 41840 700856 41846 700868
rect 42702 700856 42708 700868
rect 41840 700828 42708 700856
rect 41840 700816 41846 700828
rect 42260 700528 42288 700828
rect 42702 700816 42708 700828
rect 42760 700816 42766 700868
rect 42242 700476 42248 700528
rect 42300 700476 42306 700528
rect 674926 698980 674932 699032
rect 674984 699020 674990 699032
rect 675386 699020 675392 699032
rect 674984 698992 675392 699020
rect 674984 698980 674990 698992
rect 675386 698980 675392 698992
rect 675444 698980 675450 699032
rect 674926 696192 674932 696244
rect 674984 696192 674990 696244
rect 674944 696040 674972 696192
rect 674926 695988 674932 696040
rect 674984 695988 674990 696040
rect 675018 695920 675024 695972
rect 675076 695960 675082 695972
rect 675386 695960 675392 695972
rect 675076 695932 675392 695960
rect 675076 695920 675082 695932
rect 675386 695920 675392 695932
rect 675444 695920 675450 695972
rect 674926 695308 674932 695360
rect 674984 695348 674990 695360
rect 675386 695348 675392 695360
rect 674984 695320 675392 695348
rect 674984 695308 674990 695320
rect 675386 695308 675392 695320
rect 675444 695308 675450 695360
rect 674834 693200 674840 693252
rect 674892 693240 674898 693252
rect 675386 693240 675392 693252
rect 674892 693212 675392 693240
rect 674892 693200 674898 693212
rect 675386 693200 675392 693212
rect 675444 693200 675450 693252
rect 675018 692044 675024 692096
rect 675076 692084 675082 692096
rect 675386 692084 675392 692096
rect 675076 692056 675392 692084
rect 675076 692044 675082 692056
rect 675386 692044 675392 692056
rect 675444 692044 675450 692096
rect 675202 691636 675208 691688
rect 675260 691676 675266 691688
rect 675386 691676 675392 691688
rect 675260 691648 675392 691676
rect 675260 691636 675266 691648
rect 675386 691636 675392 691648
rect 675444 691636 675450 691688
rect 675294 691568 675300 691620
rect 675352 691568 675358 691620
rect 675312 691416 675340 691568
rect 675294 691364 675300 691416
rect 675352 691364 675358 691416
rect 675110 685176 675116 685228
rect 675168 685216 675174 685228
rect 675386 685216 675392 685228
rect 675168 685188 675392 685216
rect 675168 685176 675174 685188
rect 675386 685176 675392 685188
rect 675444 685176 675450 685228
rect 675202 684020 675208 684072
rect 675260 684060 675266 684072
rect 675386 684060 675392 684072
rect 675260 684032 675392 684060
rect 675260 684020 675266 684032
rect 675386 684020 675392 684032
rect 675444 684020 675450 684072
rect 675110 674160 675116 674212
rect 675168 674160 675174 674212
rect 675128 674008 675156 674160
rect 675110 673956 675116 674008
rect 675168 673956 675174 674008
rect 675018 671372 675024 671424
rect 675076 671412 675082 671424
rect 675202 671412 675208 671424
rect 675076 671384 675208 671412
rect 675076 671372 675082 671384
rect 675202 671372 675208 671384
rect 675260 671372 675266 671424
rect 41782 669944 41788 669996
rect 41840 669984 41846 669996
rect 42426 669984 42432 669996
rect 41840 669956 42432 669984
rect 41840 669944 41846 669956
rect 42426 669944 42432 669956
rect 42484 669944 42490 669996
rect 41782 668516 41788 668568
rect 41840 668556 41846 668568
rect 42610 668556 42616 668568
rect 41840 668528 42616 668556
rect 41840 668516 41846 668528
rect 42610 668516 42616 668528
rect 42668 668516 42674 668568
rect 42426 663116 42432 663128
rect 41800 663088 42432 663116
rect 41800 663060 41828 663088
rect 42426 663076 42432 663088
rect 42484 663076 42490 663128
rect 41782 663008 41788 663060
rect 41840 663008 41846 663060
rect 42242 663008 42248 663060
rect 42300 663048 42306 663060
rect 42300 663020 42472 663048
rect 42300 663008 42306 663020
rect 42444 662856 42472 663020
rect 42426 662804 42432 662856
rect 42484 662804 42490 662856
rect 41782 660764 41788 660816
rect 41840 660804 41846 660816
rect 42426 660804 42432 660816
rect 41840 660776 42432 660804
rect 41840 660764 41846 660776
rect 42426 660764 42432 660776
rect 42484 660764 42490 660816
rect 41782 658656 41788 658708
rect 41840 658696 41846 658708
rect 42334 658696 42340 658708
rect 41840 658668 42340 658696
rect 41840 658656 41846 658668
rect 42334 658656 42340 658668
rect 42392 658696 42398 658708
rect 42702 658696 42708 658708
rect 42392 658668 42708 658696
rect 42392 658656 42398 658668
rect 42702 658656 42708 658668
rect 42760 658656 42766 658708
rect 675110 651380 675116 651432
rect 675168 651420 675174 651432
rect 675386 651420 675392 651432
rect 675168 651392 675392 651420
rect 675168 651380 675174 651392
rect 675386 651380 675392 651392
rect 675444 651380 675450 651432
rect 674926 650088 674932 650140
rect 674984 650128 674990 650140
rect 675386 650128 675392 650140
rect 674984 650100 675392 650128
rect 674984 650088 674990 650100
rect 675386 650088 675392 650100
rect 675444 650088 675450 650140
rect 674834 647980 674840 648032
rect 674892 648020 674898 648032
rect 675386 648020 675392 648032
rect 674892 647992 675392 648020
rect 674892 647980 674898 647992
rect 675386 647980 675392 647992
rect 675444 647980 675450 648032
rect 675110 647436 675116 647488
rect 675168 647476 675174 647488
rect 675386 647476 675392 647488
rect 675168 647448 675392 647476
rect 675168 647436 675174 647448
rect 675386 647436 675392 647448
rect 675444 647436 675450 647488
rect 675202 645736 675208 645788
rect 675260 645776 675266 645788
rect 675386 645776 675392 645788
rect 675260 645748 675392 645776
rect 675260 645736 675266 645748
rect 675386 645736 675392 645748
rect 675444 645736 675450 645788
rect 675018 639752 675024 639804
rect 675076 639792 675082 639804
rect 675386 639792 675392 639804
rect 675076 639764 675392 639792
rect 675076 639752 675082 639764
rect 675386 639752 675392 639764
rect 675444 639752 675450 639804
rect 675202 638800 675208 638852
rect 675260 638840 675266 638852
rect 675386 638840 675392 638852
rect 675260 638812 675392 638840
rect 675260 638800 675266 638812
rect 675386 638800 675392 638812
rect 675444 638800 675450 638852
rect 41966 625064 41972 625116
rect 42024 625104 42030 625116
rect 42610 625104 42616 625116
rect 42024 625076 42616 625104
rect 42024 625064 42030 625076
rect 42610 625064 42616 625076
rect 42668 625064 42674 625116
rect 41782 618468 41788 618520
rect 41840 618508 41846 618520
rect 42426 618508 42432 618520
rect 41840 618480 42432 618508
rect 41840 618468 41846 618480
rect 42426 618468 42432 618480
rect 42484 618468 42490 618520
rect 42242 614932 42248 614984
rect 42300 614972 42306 614984
rect 42702 614972 42708 614984
rect 42300 614944 42708 614972
rect 42300 614932 42306 614944
rect 42702 614932 42708 614944
rect 42760 614932 42766 614984
rect 41782 613844 41788 613896
rect 41840 613884 41846 613896
rect 42334 613884 42340 613896
rect 41840 613856 42340 613884
rect 41840 613844 41846 613856
rect 42334 613844 42340 613856
rect 42392 613844 42398 613896
rect 42518 605820 42524 605872
rect 42576 605860 42582 605872
rect 42702 605860 42708 605872
rect 42576 605832 42708 605860
rect 42576 605820 42582 605832
rect 42702 605820 42708 605832
rect 42760 605820 42766 605872
rect 675110 605752 675116 605804
rect 675168 605792 675174 605804
rect 675570 605792 675576 605804
rect 675168 605764 675576 605792
rect 675168 605752 675174 605764
rect 675570 605752 675576 605764
rect 675628 605752 675634 605804
rect 674926 605480 674932 605532
rect 674984 605520 674990 605532
rect 675386 605520 675392 605532
rect 674984 605492 675392 605520
rect 674984 605480 674990 605492
rect 675386 605480 675392 605492
rect 675444 605480 675450 605532
rect 674834 602352 674840 602404
rect 674892 602392 674898 602404
rect 674892 602364 674972 602392
rect 674892 602352 674898 602364
rect 674944 602132 674972 602364
rect 674926 602080 674932 602132
rect 674984 602120 674990 602132
rect 675386 602120 675392 602132
rect 674984 602092 675392 602120
rect 674984 602080 674990 602092
rect 675386 602080 675392 602092
rect 675444 602080 675450 602132
rect 675110 601808 675116 601860
rect 675168 601848 675174 601860
rect 675386 601848 675392 601860
rect 675168 601820 675392 601848
rect 675168 601808 675174 601820
rect 675386 601808 675392 601820
rect 675444 601808 675450 601860
rect 675202 600788 675208 600840
rect 675260 600828 675266 600840
rect 675386 600828 675392 600840
rect 675260 600800 675392 600828
rect 675260 600788 675266 600800
rect 675386 600788 675392 600800
rect 675444 600788 675450 600840
rect 675018 594668 675024 594720
rect 675076 594708 675082 594720
rect 675386 594708 675392 594720
rect 675076 594680 675392 594708
rect 675076 594668 675082 594680
rect 675386 594668 675392 594680
rect 675444 594668 675450 594720
rect 675202 593784 675208 593836
rect 675260 593824 675266 593836
rect 675386 593824 675392 593836
rect 675260 593796 675392 593824
rect 675260 593784 675266 593796
rect 675386 593784 675392 593796
rect 675444 593784 675450 593836
rect 41782 583516 41788 583568
rect 41840 583556 41846 583568
rect 42426 583556 42432 583568
rect 41840 583528 42432 583556
rect 41840 583516 41846 583528
rect 42426 583516 42432 583528
rect 42484 583516 42490 583568
rect 41782 581816 41788 581868
rect 41840 581856 41846 581868
rect 42518 581856 42524 581868
rect 41840 581828 42524 581856
rect 41840 581816 41846 581828
rect 42518 581816 42524 581828
rect 42576 581816 42582 581868
rect 41782 576444 41788 576496
rect 41840 576484 41846 576496
rect 42426 576484 42432 576496
rect 41840 576456 42432 576484
rect 41840 576444 41846 576456
rect 42426 576444 42432 576456
rect 42484 576444 42490 576496
rect 42242 576240 42248 576292
rect 42300 576280 42306 576292
rect 42702 576280 42708 576292
rect 42300 576252 42708 576280
rect 42300 576240 42306 576252
rect 42702 576240 42708 576252
rect 42760 576240 42766 576292
rect 41782 574336 41788 574388
rect 41840 574376 41846 574388
rect 42426 574376 42432 574388
rect 41840 574348 42432 574376
rect 41840 574336 41846 574348
rect 42426 574336 42432 574348
rect 42484 574376 42490 574388
rect 42610 574376 42616 574388
rect 42484 574348 42616 574376
rect 42484 574336 42490 574348
rect 42610 574336 42616 574348
rect 42668 574336 42674 574388
rect 41782 571616 41788 571668
rect 41840 571656 41846 571668
rect 42610 571656 42616 571668
rect 41840 571628 42616 571656
rect 41840 571616 41846 571628
rect 42610 571616 42616 571628
rect 42668 571616 42674 571668
rect 675110 561484 675116 561536
rect 675168 561524 675174 561536
rect 675386 561524 675392 561536
rect 675168 561496 675392 561524
rect 675168 561484 675174 561496
rect 675386 561484 675392 561496
rect 675444 561484 675450 561536
rect 674834 560940 674840 560992
rect 674892 560980 674898 560992
rect 675386 560980 675392 560992
rect 674892 560952 675392 560980
rect 674892 560940 674898 560952
rect 675386 560940 675392 560952
rect 675444 560940 675450 560992
rect 674926 557812 674932 557864
rect 674984 557852 674990 557864
rect 675386 557852 675392 557864
rect 674984 557824 675392 557852
rect 674984 557812 674990 557824
rect 675386 557812 675392 557824
rect 675444 557812 675450 557864
rect 675110 557132 675116 557184
rect 675168 557172 675174 557184
rect 675386 557172 675392 557184
rect 675168 557144 675392 557172
rect 675168 557132 675174 557144
rect 675386 557132 675392 557144
rect 675444 557132 675450 557184
rect 675202 555568 675208 555620
rect 675260 555608 675266 555620
rect 675386 555608 675392 555620
rect 675260 555580 675392 555608
rect 675260 555568 675266 555580
rect 675386 555568 675392 555580
rect 675444 555568 675450 555620
rect 675018 550468 675024 550520
rect 675076 550508 675082 550520
rect 675386 550508 675392 550520
rect 675076 550480 675392 550508
rect 675076 550468 675082 550480
rect 675386 550468 675392 550480
rect 675444 550468 675450 550520
rect 41782 539112 41788 539164
rect 41840 539152 41846 539164
rect 42518 539152 42524 539164
rect 41840 539124 42524 539152
rect 41840 539112 41846 539124
rect 42518 539112 42524 539124
rect 42576 539112 42582 539164
rect 41782 532108 41788 532160
rect 41840 532148 41846 532160
rect 42426 532148 42432 532160
rect 41840 532120 42432 532148
rect 41840 532108 41846 532120
rect 42426 532108 42432 532120
rect 42484 532108 42490 532160
rect 41966 528436 41972 528488
rect 42024 528476 42030 528488
rect 42702 528476 42708 528488
rect 42024 528448 42708 528476
rect 42024 528436 42030 528448
rect 42702 528436 42708 528448
rect 42760 528436 42766 528488
rect 675294 503888 675300 503940
rect 675352 503928 675358 503940
rect 677422 503928 677428 503940
rect 675352 503900 677428 503928
rect 675352 503888 675358 503900
rect 677422 503888 677428 503900
rect 677480 503888 677486 503940
rect 674098 427796 674104 427848
rect 674156 427836 674162 427848
rect 677442 427836 677448 427848
rect 674156 427808 677448 427836
rect 674156 427796 674162 427808
rect 677442 427796 677448 427808
rect 677500 427796 677506 427848
rect 41782 412904 41788 412956
rect 41840 412944 41846 412956
rect 42334 412944 42340 412956
rect 41840 412916 42340 412944
rect 41840 412904 41846 412916
rect 42334 412904 42340 412916
rect 42392 412904 42398 412956
rect 41782 410932 41788 410984
rect 41840 410972 41846 410984
rect 42610 410972 42616 410984
rect 41840 410944 42616 410972
rect 41840 410932 41846 410944
rect 42610 410932 42616 410944
rect 42668 410932 42674 410984
rect 41782 405764 41788 405816
rect 41840 405804 41846 405816
rect 42334 405804 42340 405816
rect 41840 405776 42340 405804
rect 41840 405764 41846 405776
rect 42334 405764 42340 405776
rect 42392 405764 42398 405816
rect 41782 404472 41788 404524
rect 41840 404512 41846 404524
rect 42426 404512 42432 404524
rect 41840 404484 42432 404512
rect 41840 404472 41846 404484
rect 42426 404472 42432 404484
rect 42484 404472 42490 404524
rect 41782 400392 41788 400444
rect 41840 400432 41846 400444
rect 42426 400432 42432 400444
rect 41840 400404 42432 400432
rect 41840 400392 41846 400404
rect 42426 400392 42432 400404
rect 42484 400432 42490 400444
rect 42702 400432 42708 400444
rect 42484 400404 42708 400432
rect 42484 400392 42490 400404
rect 42702 400392 42708 400404
rect 42760 400392 42766 400444
rect 674834 383732 674840 383784
rect 674892 383772 674898 383784
rect 675386 383772 675392 383784
rect 674892 383744 675392 383772
rect 674892 383732 674898 383744
rect 675386 383732 675392 383744
rect 675444 383732 675450 383784
rect 675018 379788 675024 379840
rect 675076 379828 675082 379840
rect 675386 379828 675392 379840
rect 675076 379800 675392 379828
rect 675076 379788 675082 379800
rect 675386 379788 675392 379800
rect 675444 379788 675450 379840
rect 674834 378360 674840 378412
rect 674892 378400 674898 378412
rect 675386 378400 675392 378412
rect 674892 378372 675392 378400
rect 674892 378360 674898 378372
rect 675386 378360 675392 378372
rect 675444 378360 675450 378412
rect 674834 371424 674840 371476
rect 674892 371464 674898 371476
rect 675386 371464 675392 371476
rect 674892 371436 675392 371464
rect 674892 371424 674898 371436
rect 675386 371424 675392 371436
rect 675444 371424 675450 371476
rect 41782 369520 41788 369572
rect 41840 369560 41846 369572
rect 42334 369560 42340 369572
rect 41840 369532 42340 369560
rect 41840 369520 41846 369532
rect 42334 369520 42340 369532
rect 42392 369520 42398 369572
rect 41782 368636 41788 368688
rect 41840 368676 41846 368688
rect 42610 368676 42616 368688
rect 41840 368648 42616 368676
rect 41840 368636 41846 368648
rect 42610 368636 42616 368648
rect 42668 368636 42674 368688
rect 41782 362584 41788 362636
rect 41840 362624 41846 362636
rect 42334 362624 42340 362636
rect 41840 362596 42340 362624
rect 41840 362584 41846 362596
rect 42334 362584 42340 362596
rect 42392 362584 42398 362636
rect 41782 360340 41788 360392
rect 41840 360380 41846 360392
rect 42518 360380 42524 360392
rect 41840 360352 42524 360380
rect 41840 360340 41846 360352
rect 42518 360340 42524 360352
rect 42576 360380 42582 360392
rect 42702 360380 42708 360392
rect 42576 360352 42708 360380
rect 42576 360340 42582 360352
rect 42702 360340 42708 360352
rect 42760 360340 42766 360392
rect 41782 357212 41788 357264
rect 41840 357252 41846 357264
rect 42426 357252 42432 357264
rect 41840 357224 42432 357252
rect 41840 357212 41846 357224
rect 42260 357060 42288 357224
rect 42426 357212 42432 357224
rect 42484 357212 42490 357264
rect 42242 357008 42248 357060
rect 42300 357008 42306 357060
rect 675110 338784 675116 338836
rect 675168 338824 675174 338836
rect 675386 338824 675392 338836
rect 675168 338796 675392 338824
rect 675168 338784 675174 338796
rect 675386 338784 675392 338796
rect 675444 338784 675450 338836
rect 674926 337492 674932 337544
rect 674984 337532 674990 337544
rect 675386 337532 675392 337544
rect 674984 337504 675392 337532
rect 674984 337492 674990 337504
rect 675386 337492 675392 337504
rect 675444 337492 675450 337544
rect 675018 335384 675024 335436
rect 675076 335424 675082 335436
rect 675202 335424 675208 335436
rect 675076 335396 675208 335424
rect 675076 335384 675082 335396
rect 675202 335384 675208 335396
rect 675260 335424 675266 335436
rect 675386 335424 675392 335436
rect 675260 335396 675392 335424
rect 675260 335384 675266 335396
rect 675386 335384 675392 335396
rect 675444 335384 675450 335436
rect 675018 334228 675024 334280
rect 675076 334268 675082 334280
rect 675386 334268 675392 334280
rect 675076 334240 675392 334268
rect 675076 334228 675082 334240
rect 675386 334228 675392 334240
rect 675444 334228 675450 334280
rect 674834 328040 674840 328092
rect 674892 328080 674898 328092
rect 675110 328080 675116 328092
rect 674892 328052 675116 328080
rect 674892 328040 674898 328052
rect 675110 328040 675116 328052
rect 675168 328080 675174 328092
rect 675386 328080 675392 328092
rect 675168 328052 675392 328080
rect 675168 328040 675174 328052
rect 675386 328040 675392 328052
rect 675444 328040 675450 328092
rect 41782 326340 41788 326392
rect 41840 326380 41846 326392
rect 42426 326380 42432 326392
rect 41840 326352 42432 326380
rect 41840 326340 41846 326352
rect 42426 326340 42432 326352
rect 42484 326340 42490 326392
rect 41782 325116 41788 325168
rect 41840 325156 41846 325168
rect 42518 325156 42524 325168
rect 41840 325128 42524 325156
rect 41840 325116 41846 325128
rect 42518 325116 42524 325128
rect 42576 325116 42582 325168
rect 41782 319404 41788 319456
rect 41840 319444 41846 319456
rect 42426 319444 42432 319456
rect 41840 319416 42432 319444
rect 41840 319404 41846 319416
rect 42426 319404 42432 319416
rect 42484 319404 42490 319456
rect 41782 318724 41788 318776
rect 41840 318764 41846 318776
rect 42334 318764 42340 318776
rect 41840 318736 42340 318764
rect 41840 318724 41846 318736
rect 42334 318724 42340 318736
rect 42392 318724 42398 318776
rect 41782 318112 41788 318164
rect 41840 318152 41846 318164
rect 42702 318152 42708 318164
rect 41840 318124 42708 318152
rect 41840 318112 41846 318124
rect 42702 318112 42708 318124
rect 42760 318112 42766 318164
rect 41782 313488 41788 313540
rect 41840 313528 41846 313540
rect 42334 313528 42340 313540
rect 41840 313500 42340 313528
rect 41840 313488 41846 313500
rect 42334 313488 42340 313500
rect 42392 313488 42398 313540
rect 675018 294108 675024 294160
rect 675076 294148 675082 294160
rect 675386 294148 675392 294160
rect 675076 294120 675392 294148
rect 675076 294108 675082 294120
rect 675386 294108 675392 294120
rect 675444 294108 675450 294160
rect 674926 293224 674932 293276
rect 674984 293264 674990 293276
rect 675386 293264 675392 293276
rect 674984 293236 675392 293264
rect 674984 293224 674990 293236
rect 675386 293224 675392 293236
rect 675444 293224 675450 293276
rect 674926 289484 674932 289536
rect 674984 289524 674990 289536
rect 675110 289524 675116 289536
rect 674984 289496 675116 289524
rect 674984 289484 674990 289496
rect 675110 289484 675116 289496
rect 675168 289524 675174 289536
rect 675386 289524 675392 289536
rect 675168 289496 675392 289524
rect 675168 289484 675174 289496
rect 675386 289484 675392 289496
rect 675444 289484 675450 289536
rect 675018 288600 675024 288652
rect 675076 288640 675082 288652
rect 675294 288640 675300 288652
rect 675076 288612 675300 288640
rect 675076 288600 675082 288612
rect 675294 288600 675300 288612
rect 675352 288600 675358 288652
rect 41782 283160 41788 283212
rect 41840 283200 41846 283212
rect 42426 283200 42432 283212
rect 41840 283172 42432 283200
rect 41840 283160 41846 283172
rect 42426 283160 42432 283172
rect 42484 283160 42490 283212
rect 674834 282276 674840 282328
rect 674892 282316 674898 282328
rect 675386 282316 675392 282328
rect 674892 282288 675392 282316
rect 674892 282276 674898 282288
rect 675386 282276 675392 282288
rect 675444 282276 675450 282328
rect 41782 282072 41788 282124
rect 41840 282112 41846 282124
rect 42518 282112 42524 282124
rect 41840 282084 42524 282112
rect 41840 282072 41846 282084
rect 42518 282072 42524 282084
rect 42576 282072 42582 282124
rect 675202 281188 675208 281240
rect 675260 281228 675266 281240
rect 675386 281228 675392 281240
rect 675260 281200 675392 281228
rect 675260 281188 675266 281200
rect 675386 281188 675392 281200
rect 675444 281188 675450 281240
rect 41782 276156 41788 276208
rect 41840 276196 41846 276208
rect 42426 276196 42432 276208
rect 41840 276168 42432 276196
rect 41840 276156 41846 276168
rect 42426 276156 42432 276168
rect 42484 276156 42490 276208
rect 41782 274524 41788 274576
rect 41840 274564 41846 274576
rect 42334 274564 42340 274576
rect 41840 274536 42340 274564
rect 41840 274524 41846 274536
rect 42334 274524 42340 274536
rect 42392 274524 42398 274576
rect 41782 273912 41788 273964
rect 41840 273952 41846 273964
rect 42610 273952 42616 273964
rect 41840 273924 42616 273952
rect 41840 273912 41846 273924
rect 42610 273912 42616 273924
rect 42668 273912 42674 273964
rect 41782 270580 41788 270632
rect 41840 270620 41846 270632
rect 42334 270620 42340 270632
rect 41840 270592 42340 270620
rect 41840 270580 41846 270592
rect 42334 270580 42340 270592
rect 42392 270580 42398 270632
rect 675110 248752 675116 248804
rect 675168 248792 675174 248804
rect 675386 248792 675392 248804
rect 675168 248764 675392 248792
rect 675168 248752 675174 248764
rect 675386 248752 675392 248764
rect 675444 248752 675450 248804
rect 675018 247460 675024 247512
rect 675076 247500 675082 247512
rect 675386 247500 675392 247512
rect 675076 247472 675392 247500
rect 675076 247460 675082 247472
rect 675386 247460 675392 247472
rect 675444 247460 675450 247512
rect 674926 244468 674932 244520
rect 674984 244508 674990 244520
rect 675386 244508 675392 244520
rect 674984 244480 675392 244508
rect 674984 244468 674990 244480
rect 675386 244468 675392 244480
rect 675444 244468 675450 244520
rect 41782 239912 41788 239964
rect 41840 239952 41846 239964
rect 42426 239952 42432 239964
rect 41840 239924 42432 239952
rect 41840 239912 41846 239924
rect 42426 239912 42432 239924
rect 42484 239912 42490 239964
rect 41782 238484 41788 238536
rect 41840 238524 41846 238536
rect 42518 238524 42524 238536
rect 41840 238496 42524 238524
rect 41840 238484 41846 238496
rect 42518 238484 42524 238496
rect 42576 238484 42582 238536
rect 674834 237668 674840 237720
rect 674892 237708 674898 237720
rect 675386 237708 675392 237720
rect 674892 237680 675392 237708
rect 674892 237668 674898 237680
rect 675386 237668 675392 237680
rect 675444 237668 675450 237720
rect 675202 236240 675208 236292
rect 675260 236280 675266 236292
rect 675386 236280 675392 236292
rect 675260 236252 675392 236280
rect 675260 236240 675266 236252
rect 675386 236240 675392 236252
rect 675444 236240 675450 236292
rect 41782 232976 41788 233028
rect 41840 233016 41846 233028
rect 42426 233016 42432 233028
rect 41840 232988 42432 233016
rect 41840 232976 41846 232988
rect 42426 232976 42432 232988
rect 42484 232976 42490 233028
rect 41782 232364 41788 232416
rect 41840 232404 41846 232416
rect 42334 232404 42340 232416
rect 41840 232376 42340 232404
rect 41840 232364 41846 232376
rect 42334 232364 42340 232376
rect 42392 232364 42398 232416
rect 41782 231684 41788 231736
rect 41840 231724 41846 231736
rect 42610 231724 42616 231736
rect 41840 231696 42616 231724
rect 41840 231684 41846 231696
rect 42610 231684 42616 231696
rect 42668 231684 42674 231736
rect 41782 227060 41788 227112
rect 41840 227100 41846 227112
rect 42334 227100 42340 227112
rect 41840 227072 42340 227100
rect 41840 227060 41846 227072
rect 42334 227060 42340 227072
rect 42392 227060 42398 227112
rect 675110 203464 675116 203516
rect 675168 203504 675174 203516
rect 675294 203504 675300 203516
rect 675168 203476 675300 203504
rect 675168 203464 675174 203476
rect 675294 203464 675300 203476
rect 675352 203464 675358 203516
rect 675018 202308 675024 202360
rect 675076 202348 675082 202360
rect 675386 202348 675392 202360
rect 675076 202320 675392 202348
rect 675076 202308 675082 202320
rect 675386 202308 675392 202320
rect 675444 202308 675450 202360
rect 674926 200200 674932 200252
rect 674984 200240 674990 200252
rect 675386 200240 675392 200252
rect 674984 200212 675392 200240
rect 674984 200200 674990 200212
rect 675386 200200 675392 200212
rect 675444 200200 675450 200252
rect 675202 199248 675208 199300
rect 675260 199248 675266 199300
rect 675220 199096 675248 199248
rect 675202 199044 675208 199096
rect 675260 199044 675266 199096
rect 41782 196732 41788 196784
rect 41840 196772 41846 196784
rect 42702 196772 42708 196784
rect 41840 196744 42708 196772
rect 41840 196732 41846 196744
rect 42702 196732 42708 196744
rect 42760 196732 42766 196784
rect 41782 195304 41788 195356
rect 41840 195344 41846 195356
rect 42426 195344 42432 195356
rect 41840 195316 42432 195344
rect 41840 195304 41846 195316
rect 42426 195304 42432 195316
rect 42484 195304 42490 195356
rect 675202 191904 675208 191956
rect 675260 191944 675266 191956
rect 675386 191944 675392 191956
rect 675260 191916 675392 191944
rect 675260 191904 675266 191916
rect 675386 191904 675392 191916
rect 675444 191904 675450 191956
rect 41782 189796 41788 189848
rect 41840 189836 41846 189848
rect 42702 189836 42708 189848
rect 41840 189808 42708 189836
rect 41840 189796 41846 189808
rect 42702 189796 42708 189808
rect 42760 189796 42766 189848
rect 41782 188096 41788 188148
rect 41840 188136 41846 188148
rect 42334 188136 42340 188148
rect 41840 188108 42340 188136
rect 41840 188096 41846 188108
rect 42334 188096 42340 188108
rect 42392 188096 42398 188148
rect 41782 187552 41788 187604
rect 41840 187592 41846 187604
rect 42518 187592 42524 187604
rect 41840 187564 42524 187592
rect 41840 187552 41846 187564
rect 42518 187552 42524 187564
rect 42576 187552 42582 187604
rect 41782 184152 41788 184204
rect 41840 184192 41846 184204
rect 42334 184192 42340 184204
rect 41840 184164 42340 184192
rect 41840 184152 41846 184164
rect 42334 184152 42340 184164
rect 42392 184152 42398 184204
rect 675294 158720 675300 158772
rect 675352 158720 675358 158772
rect 675110 158516 675116 158568
rect 675168 158556 675174 158568
rect 675312 158556 675340 158720
rect 675168 158528 675340 158556
rect 675168 158516 675174 158528
rect 674834 157292 674840 157344
rect 674892 157332 674898 157344
rect 675018 157332 675024 157344
rect 674892 157304 675024 157332
rect 674892 157292 674898 157304
rect 675018 157292 675024 157304
rect 675076 157332 675082 157344
rect 675386 157332 675392 157344
rect 675076 157304 675392 157332
rect 675076 157292 675082 157304
rect 675386 157292 675392 157304
rect 675444 157292 675450 157344
rect 674926 155184 674932 155236
rect 674984 155224 674990 155236
rect 675386 155224 675392 155236
rect 674984 155196 675392 155224
rect 674984 155184 674990 155196
rect 675386 155184 675392 155196
rect 675444 155184 675450 155236
rect 675018 147092 675024 147144
rect 675076 147132 675082 147144
rect 675202 147132 675208 147144
rect 675076 147104 675208 147132
rect 675076 147092 675082 147104
rect 675202 147092 675208 147104
rect 675260 147132 675266 147144
rect 675386 147132 675392 147144
rect 675260 147104 675392 147132
rect 675260 147092 675266 147104
rect 675386 147092 675392 147104
rect 675444 147092 675450 147144
rect 675018 113092 675024 113144
rect 675076 113132 675082 113144
rect 675386 113132 675392 113144
rect 675076 113104 675392 113132
rect 675076 113092 675082 113104
rect 675386 113092 675392 113104
rect 675444 113092 675450 113144
rect 674834 112480 674840 112532
rect 674892 112520 674898 112532
rect 675386 112520 675392 112532
rect 674892 112492 675392 112520
rect 674892 112480 674898 112492
rect 675386 112480 675392 112492
rect 675444 112480 675450 112532
rect 674926 109080 674932 109132
rect 674984 109120 674990 109132
rect 675386 109120 675392 109132
rect 674984 109092 675392 109120
rect 674984 109080 674990 109092
rect 675386 109080 675392 109092
rect 675444 109080 675450 109132
rect 675018 108808 675024 108860
rect 675076 108848 675082 108860
rect 675386 108848 675392 108860
rect 675076 108820 675392 108848
rect 675076 108808 675082 108820
rect 675386 108808 675392 108820
rect 675444 108808 675450 108860
rect 675202 107788 675208 107840
rect 675260 107828 675266 107840
rect 675386 107828 675392 107840
rect 675260 107800 675392 107828
rect 675260 107788 675266 107800
rect 675386 107788 675392 107800
rect 675444 107788 675450 107840
rect 675202 102008 675208 102060
rect 675260 102008 675266 102060
rect 675220 101844 675248 102008
rect 675294 101844 675300 101856
rect 675220 101816 675300 101844
rect 675294 101804 675300 101816
rect 675352 101804 675358 101856
rect 527450 43156 527456 43208
rect 527508 43196 527514 43208
rect 527508 43168 528014 43196
rect 527508 43156 527514 43168
rect 523770 43088 523776 43140
rect 523828 43128 523834 43140
rect 523828 43100 527946 43128
rect 523828 43088 523834 43100
rect 516134 43020 516140 43072
rect 516192 43060 516198 43072
rect 516192 43032 527878 43060
rect 516192 43020 516198 43032
rect 459646 42952 459652 43004
rect 459704 42992 459710 43004
rect 467650 42992 467656 43004
rect 459704 42964 467656 42992
rect 459704 42952 459710 42964
rect 467650 42952 467656 42964
rect 467708 42952 467714 43004
rect 415302 42884 415308 42936
rect 415360 42924 415366 42936
rect 467834 42924 467840 42936
rect 415360 42896 467840 42924
rect 415360 42884 415366 42896
rect 467834 42884 467840 42896
rect 467892 42884 467898 42936
rect 473262 42884 473268 42936
rect 473320 42924 473326 42936
rect 526806 42924 526812 42936
rect 473320 42896 526812 42924
rect 473320 42884 473326 42896
rect 526806 42884 526812 42896
rect 526864 42884 526870 42936
rect 411070 42816 411076 42868
rect 411128 42856 411134 42868
rect 419718 42856 419724 42868
rect 411128 42828 419724 42856
rect 411128 42816 411134 42828
rect 419718 42816 419724 42828
rect 419776 42816 419782 42868
rect 461486 42856 461492 42868
rect 451246 42828 461492 42856
rect 195974 42760 195980 42772
rect 186138 42732 195980 42760
rect 42150 42428 42156 42480
rect 42208 42468 42214 42480
rect 147674 42468 147680 42480
rect 42208 42440 147680 42468
rect 42208 42428 42214 42440
rect 147674 42428 147680 42440
rect 147732 42428 147738 42480
rect 42058 42360 42064 42412
rect 42116 42400 42122 42412
rect 186138 42400 186166 42732
rect 195974 42720 195980 42732
rect 196032 42720 196038 42772
rect 295242 42748 295248 42800
rect 295300 42788 295306 42800
rect 303246 42788 303252 42800
rect 295300 42760 303252 42788
rect 295300 42748 295306 42760
rect 303246 42748 303252 42760
rect 303304 42748 303310 42800
rect 350074 42748 350080 42800
rect 350132 42788 350138 42800
rect 358078 42788 358084 42800
rect 350132 42760 358084 42788
rect 350132 42748 350138 42760
rect 358078 42748 358084 42760
rect 358136 42748 358142 42800
rect 360562 42748 360568 42800
rect 360620 42788 360626 42800
rect 406746 42788 406752 42800
rect 360620 42760 406752 42788
rect 360620 42748 360626 42760
rect 406746 42748 406752 42760
rect 406804 42788 406810 42800
rect 451246 42788 451274 42828
rect 461486 42816 461492 42828
rect 461544 42856 461550 42868
rect 516134 42856 516140 42868
rect 461544 42828 516140 42856
rect 461544 42816 461550 42828
rect 516134 42816 516140 42828
rect 516192 42816 516198 42868
rect 406804 42760 451274 42788
rect 406804 42748 406810 42760
rect 467834 42748 467840 42800
rect 467892 42788 467898 42800
rect 468938 42788 468944 42800
rect 467892 42760 468944 42788
rect 467892 42748 467898 42760
rect 468938 42748 468944 42760
rect 468996 42788 469002 42800
rect 523770 42788 523776 42800
rect 468996 42760 523776 42788
rect 468996 42748 469002 42760
rect 523770 42748 523776 42760
rect 523828 42748 523834 42800
rect 307570 42720 307576 42732
rect 200086 42692 307576 42720
rect 199010 42652 199016 42664
rect 42116 42372 186166 42400
rect 186246 42624 199016 42652
rect 42116 42360 42122 42372
rect 88794 42252 88800 42304
rect 88852 42292 88858 42304
rect 186246 42292 186274 42624
rect 199010 42612 199016 42624
rect 199068 42652 199074 42664
rect 200086 42652 200114 42692
rect 307570 42680 307576 42692
rect 307628 42720 307634 42732
rect 362402 42720 362408 42732
rect 307628 42692 362408 42720
rect 307628 42680 307634 42692
rect 362402 42680 362408 42692
rect 362460 42720 362466 42732
rect 417234 42720 417240 42732
rect 362460 42692 417240 42720
rect 362460 42680 362466 42692
rect 417234 42680 417240 42692
rect 417292 42720 417298 42732
rect 471974 42720 471980 42732
rect 417292 42692 471980 42720
rect 417292 42680 417298 42692
rect 471974 42680 471980 42692
rect 472032 42720 472038 42732
rect 473262 42720 473268 42732
rect 472032 42692 473268 42720
rect 472032 42680 472038 42692
rect 473262 42680 473268 42692
rect 473320 42680 473326 42732
rect 514478 42680 514484 42732
rect 514536 42720 514542 42732
rect 522482 42720 522488 42732
rect 514536 42692 522488 42720
rect 514536 42680 514542 42692
rect 522482 42680 522488 42692
rect 522540 42680 522546 42732
rect 199068 42624 200114 42652
rect 199068 42612 199074 42624
rect 200850 42612 200856 42664
rect 200908 42652 200914 42664
rect 241330 42652 241336 42664
rect 200908 42624 241336 42652
rect 200908 42612 200914 42624
rect 241330 42612 241336 42624
rect 241388 42652 241394 42664
rect 297726 42652 297732 42664
rect 241388 42624 297732 42652
rect 241388 42612 241394 42624
rect 297726 42612 297732 42624
rect 297784 42652 297790 42664
rect 300762 42652 300768 42664
rect 297784 42624 300768 42652
rect 297784 42612 297790 42624
rect 300762 42612 300768 42624
rect 300820 42652 300826 42664
rect 305086 42652 305092 42664
rect 300820 42624 305092 42652
rect 300820 42612 300826 42624
rect 305086 42612 305092 42624
rect 305144 42612 305150 42664
rect 309410 42612 309416 42664
rect 309468 42652 309474 42664
rect 352558 42652 352564 42664
rect 309468 42624 352564 42652
rect 309468 42612 309474 42624
rect 352558 42612 352564 42624
rect 352616 42652 352622 42664
rect 355594 42652 355600 42664
rect 352616 42624 355600 42652
rect 352616 42612 352622 42624
rect 355594 42612 355600 42624
rect 355652 42652 355658 42664
rect 359918 42652 359924 42664
rect 355652 42624 359924 42652
rect 355652 42612 355658 42624
rect 359918 42612 359924 42624
rect 359976 42612 359982 42664
rect 364242 42612 364248 42664
rect 364300 42652 364306 42664
rect 407390 42652 407396 42664
rect 364300 42624 407396 42652
rect 364300 42612 364306 42624
rect 407390 42612 407396 42624
rect 407448 42652 407454 42664
rect 410426 42652 410432 42664
rect 407448 42624 410432 42652
rect 407448 42612 407454 42624
rect 410426 42612 410432 42624
rect 410484 42612 410490 42664
rect 416038 42612 416044 42664
rect 416096 42652 416102 42664
rect 419074 42652 419080 42664
rect 416096 42624 419080 42652
rect 416096 42612 416102 42624
rect 419074 42612 419080 42624
rect 419132 42652 419138 42664
rect 462130 42652 462136 42664
rect 419132 42624 462136 42652
rect 419132 42612 419138 42624
rect 462130 42612 462136 42624
rect 462188 42652 462194 42664
rect 465166 42652 465172 42664
rect 462188 42624 465172 42652
rect 462188 42612 462194 42624
rect 465166 42612 465172 42624
rect 465224 42612 465230 42664
rect 470778 42612 470784 42664
rect 470836 42652 470842 42664
rect 473814 42652 473820 42664
rect 470836 42624 473820 42652
rect 470836 42612 470842 42624
rect 473814 42612 473820 42624
rect 473872 42652 473878 42664
rect 516962 42652 516968 42664
rect 473872 42624 516968 42652
rect 473872 42612 473878 42624
rect 516962 42612 516968 42624
rect 517020 42652 517026 42664
rect 519998 42652 520004 42664
rect 517020 42624 520004 42652
rect 517020 42612 517026 42624
rect 519998 42612 520004 42624
rect 520056 42612 520062 42664
rect 188522 42544 188528 42596
rect 188580 42584 188586 42596
rect 192846 42584 192852 42596
rect 188580 42556 192852 42584
rect 188580 42544 188586 42556
rect 192846 42544 192852 42556
rect 192904 42584 192910 42596
rect 201494 42584 201500 42596
rect 192904 42556 201500 42584
rect 192904 42544 192910 42556
rect 201494 42544 201500 42556
rect 201552 42584 201558 42596
rect 297082 42584 297088 42596
rect 201552 42556 297088 42584
rect 201552 42544 201558 42556
rect 297082 42544 297088 42556
rect 297140 42584 297146 42596
rect 299566 42584 299572 42596
rect 297140 42556 299572 42584
rect 297140 42544 297146 42556
rect 299566 42544 299572 42556
rect 299624 42584 299630 42596
rect 305730 42584 305736 42596
rect 299624 42556 305736 42584
rect 299624 42544 299630 42556
rect 305730 42544 305736 42556
rect 305788 42584 305794 42596
rect 351914 42584 351920 42596
rect 305788 42556 351920 42584
rect 305788 42544 305794 42556
rect 351914 42544 351920 42556
rect 351972 42584 351978 42596
rect 354398 42584 354404 42596
rect 351972 42556 354404 42584
rect 351972 42544 351978 42556
rect 354398 42544 354404 42556
rect 354456 42584 354462 42596
rect 360562 42584 360568 42596
rect 354456 42556 360568 42584
rect 354456 42544 354462 42556
rect 360562 42544 360568 42556
rect 360620 42544 360626 42596
rect 404906 42544 404912 42596
rect 404964 42584 404970 42596
rect 412910 42584 412916 42596
rect 404964 42556 412916 42584
rect 404964 42544 404970 42556
rect 412910 42544 412916 42556
rect 412968 42544 412974 42596
rect 413554 42544 413560 42596
rect 413612 42584 413618 42596
rect 417878 42584 417884 42596
rect 413612 42556 417884 42584
rect 413612 42544 413618 42556
rect 417878 42544 417884 42556
rect 417936 42584 417942 42596
rect 468294 42584 468300 42596
rect 417936 42556 468300 42584
rect 417936 42544 417942 42556
rect 468294 42544 468300 42556
rect 468352 42584 468358 42596
rect 472618 42584 472624 42596
rect 468352 42556 472624 42584
rect 468352 42544 468358 42556
rect 472618 42544 472624 42556
rect 472676 42584 472682 42596
rect 523126 42584 523132 42596
rect 472676 42556 523132 42584
rect 472676 42544 472682 42556
rect 523126 42544 523132 42556
rect 523184 42584 523190 42596
rect 527450 42584 527456 42596
rect 523184 42556 527456 42584
rect 523184 42544 523190 42556
rect 527450 42544 527456 42556
rect 527508 42544 527514 42596
rect 199654 42476 199660 42528
rect 199712 42516 199718 42528
rect 303890 42516 303896 42528
rect 199712 42488 303896 42516
rect 199712 42476 199718 42488
rect 303890 42476 303896 42488
rect 303948 42516 303954 42528
rect 308214 42516 308220 42528
rect 303948 42488 308220 42516
rect 303948 42476 303954 42488
rect 308214 42476 308220 42488
rect 308272 42516 308278 42528
rect 358722 42516 358728 42528
rect 308272 42488 358728 42516
rect 308272 42476 308278 42488
rect 358722 42476 358728 42488
rect 358780 42516 358786 42528
rect 363046 42516 363052 42528
rect 358780 42488 363052 42516
rect 358780 42476 358786 42488
rect 363046 42476 363052 42488
rect 363104 42516 363110 42528
rect 413572 42516 413600 42544
rect 363104 42488 413600 42516
rect 363104 42476 363110 42488
rect 465810 42476 465816 42528
rect 465868 42516 465874 42528
rect 474458 42516 474464 42528
rect 465868 42488 474464 42516
rect 465868 42476 465874 42488
rect 474458 42476 474464 42488
rect 474516 42476 474522 42528
rect 527850 42460 527878 43032
rect 527918 42528 527946 43100
rect 527986 42596 528014 43168
rect 527986 42568 530996 42596
rect 527918 42500 530928 42528
rect 188522 42448 188528 42460
rect 88852 42264 186274 42292
rect 186450 42420 188528 42448
rect 88852 42252 88858 42264
rect 42242 42100 42248 42152
rect 42300 42140 42306 42152
rect 140958 42140 140964 42152
rect 42300 42112 140964 42140
rect 42300 42100 42306 42112
rect 140958 42100 140964 42112
rect 141016 42100 141022 42152
rect 42334 42032 42340 42084
rect 42392 42072 42398 42084
rect 145098 42072 145104 42084
rect 42392 42044 145104 42072
rect 42392 42032 42398 42044
rect 145098 42032 145104 42044
rect 145156 42032 145162 42084
rect 147674 42048 147680 42100
rect 147732 42088 147738 42100
rect 186450 42088 186478 42420
rect 188522 42408 188528 42420
rect 188580 42408 188586 42460
rect 195974 42408 195980 42460
rect 196032 42448 196038 42460
rect 304534 42448 304540 42460
rect 196032 42420 304540 42448
rect 196032 42408 196038 42420
rect 304534 42408 304540 42420
rect 304592 42448 304598 42460
rect 359366 42448 359372 42460
rect 304592 42420 359372 42448
rect 304592 42408 304598 42420
rect 359366 42408 359372 42420
rect 359424 42448 359430 42460
rect 414198 42448 414204 42460
rect 359424 42420 414204 42448
rect 359424 42408 359430 42420
rect 414198 42408 414204 42420
rect 414256 42448 414262 42460
rect 415302 42448 415308 42460
rect 414256 42420 415308 42448
rect 414256 42408 414262 42420
rect 415302 42408 415308 42420
rect 415360 42408 415366 42460
rect 527850 42432 530860 42460
rect 186682 42340 186688 42392
rect 186740 42380 186746 42392
rect 194686 42380 194692 42392
rect 186740 42352 194692 42380
rect 186740 42340 186746 42352
rect 194686 42340 194692 42352
rect 194744 42340 194750 42392
rect 409230 42340 409236 42392
rect 409288 42380 409294 42392
rect 412266 42380 412272 42392
rect 409288 42352 412272 42380
rect 409288 42340 409294 42352
rect 412266 42340 412272 42352
rect 412324 42380 412330 42392
rect 415394 42380 415400 42392
rect 412324 42352 415400 42380
rect 412324 42340 412330 42352
rect 415394 42340 415400 42352
rect 415452 42340 415458 42392
rect 518802 42340 518808 42392
rect 518860 42380 518866 42392
rect 524966 42380 524972 42392
rect 518860 42352 524972 42380
rect 518860 42340 518866 42352
rect 524966 42340 524972 42352
rect 525024 42340 525030 42392
rect 147732 42060 186478 42088
rect 238464 42096 253268 42124
rect 147732 42048 147738 42060
rect 198458 41896 198464 41948
rect 198516 41936 198522 41948
rect 200114 41936 200120 41948
rect 198516 41908 200120 41936
rect 198516 41896 198522 41908
rect 200114 41896 200120 41908
rect 200172 41896 200178 41948
rect 186130 41828 186136 41880
rect 186188 41868 186194 41880
rect 195238 41868 195244 41880
rect 186188 41840 195244 41868
rect 186188 41828 186194 41840
rect 195238 41828 195244 41840
rect 195296 41868 195302 41880
rect 199562 41868 199568 41880
rect 195296 41840 199568 41868
rect 195296 41828 195302 41840
rect 199562 41828 199568 41840
rect 199620 41828 199626 41880
rect 189258 41760 189264 41812
rect 189316 41800 189322 41812
rect 191098 41800 191104 41812
rect 189316 41772 191104 41800
rect 189316 41760 189322 41772
rect 191098 41760 191104 41772
rect 191156 41800 191162 41812
rect 192294 41800 192300 41812
rect 191156 41772 192300 41800
rect 191156 41760 191162 41772
rect 192294 41760 192300 41772
rect 192352 41800 192358 41812
rect 193582 41800 193588 41812
rect 192352 41772 193588 41800
rect 192352 41760 192358 41772
rect 193582 41760 193588 41772
rect 193640 41800 193646 41812
rect 196434 41800 196440 41812
rect 193640 41772 196440 41800
rect 193640 41760 193646 41772
rect 196434 41760 196440 41772
rect 196492 41760 196498 41812
rect 143074 41420 143080 41472
rect 143132 41460 143138 41472
rect 143132 41432 144684 41460
rect 143132 41420 143138 41432
rect 144656 41404 144684 41432
rect 145098 41420 145104 41472
rect 145156 41460 145162 41472
rect 186130 41460 186136 41472
rect 145156 41432 186136 41460
rect 145156 41420 145162 41432
rect 186130 41420 186136 41432
rect 186188 41420 186194 41472
rect 186286 41432 202552 41460
rect 144638 41352 144644 41404
rect 144696 41392 144702 41404
rect 186286 41392 186314 41432
rect 144696 41364 186314 41392
rect 202524 41392 202552 41432
rect 238464 41392 238492 42096
rect 202524 41364 238492 41392
rect 253240 41392 253268 42096
rect 469674 41964 469680 42016
rect 469732 42004 469738 42016
rect 470686 42004 470692 42016
rect 469732 41976 470692 42004
rect 469732 41964 469738 41976
rect 470686 41964 470692 41976
rect 470744 41964 470750 42016
rect 305270 41896 305276 41948
rect 305328 41936 305334 41948
rect 306282 41936 306288 41948
rect 305328 41908 306288 41936
rect 305328 41896 305334 41908
rect 306282 41896 306288 41908
rect 306340 41936 306346 41948
rect 308674 41936 308680 41948
rect 306340 41908 308680 41936
rect 306340 41896 306346 41908
rect 308674 41896 308680 41908
rect 308732 41896 308738 41948
rect 464154 41828 464160 41880
rect 464212 41868 464218 41880
rect 467190 41868 467196 41880
rect 464212 41840 467196 41868
rect 464212 41828 464218 41840
rect 467190 41828 467196 41840
rect 467248 41868 467254 41880
rect 470042 41868 470048 41880
rect 467248 41840 470048 41868
rect 467248 41828 467254 41840
rect 470042 41828 470048 41840
rect 470100 41828 470106 41880
rect 360010 41760 360016 41812
rect 360068 41800 360074 41812
rect 361114 41800 361120 41812
rect 360068 41772 361120 41800
rect 360068 41760 360074 41772
rect 361114 41760 361120 41772
rect 361172 41800 361178 41812
rect 363506 41800 363512 41812
rect 361172 41772 363512 41800
rect 361172 41760 361178 41772
rect 363506 41760 363512 41772
rect 363564 41760 363570 41812
rect 410518 41760 410524 41812
rect 410576 41800 410582 41812
rect 411530 41800 411536 41812
rect 410576 41772 411536 41800
rect 410576 41760 410582 41772
rect 411530 41760 411536 41772
rect 411588 41800 411594 41812
rect 414842 41800 414848 41812
rect 411588 41772 414848 41800
rect 411588 41760 411594 41772
rect 414842 41760 414848 41772
rect 414900 41800 414906 41812
rect 415854 41800 415860 41812
rect 414900 41772 415860 41800
rect 414900 41760 414906 41772
rect 415854 41760 415860 41772
rect 415912 41760 415918 41812
rect 465350 41760 465356 41812
rect 465408 41800 465414 41812
rect 466362 41800 466368 41812
rect 465408 41772 466368 41800
rect 465408 41760 465414 41772
rect 466362 41760 466368 41772
rect 466420 41800 466426 41812
rect 469398 41800 469404 41812
rect 466420 41772 469404 41800
rect 466420 41760 466426 41772
rect 469398 41760 469404 41772
rect 469456 41760 469462 41812
rect 520090 41760 520096 41812
rect 520148 41800 520154 41812
rect 521194 41800 521200 41812
rect 520148 41772 521200 41800
rect 520148 41760 520154 41772
rect 521194 41760 521200 41772
rect 521252 41800 521258 41812
rect 524230 41800 524236 41812
rect 521252 41772 524236 41800
rect 521252 41760 521258 41772
rect 524230 41760 524236 41772
rect 524288 41800 524294 41812
rect 525518 41800 525524 41812
rect 524288 41772 525524 41800
rect 524288 41760 524294 41772
rect 525518 41760 525524 41772
rect 525576 41800 525582 41812
rect 527910 41800 527916 41812
rect 525576 41772 527916 41800
rect 525576 41760 525582 41772
rect 527910 41760 527916 41772
rect 527968 41760 527974 41812
rect 294852 41432 311142 41460
rect 294852 41392 294880 41432
rect 253240 41364 294880 41392
rect 311114 41392 311142 41432
rect 349632 41432 365944 41460
rect 349632 41392 349660 41432
rect 311114 41364 349660 41392
rect 365916 41392 365944 41432
rect 404464 41432 420776 41460
rect 404464 41392 404492 41432
rect 365916 41364 404492 41392
rect 420748 41392 420776 41432
rect 459246 41432 475516 41460
rect 459246 41392 459274 41432
rect 420748 41364 459274 41392
rect 475488 41392 475516 41432
rect 514036 41432 530748 41460
rect 514036 41392 514064 41432
rect 475488 41364 514064 41392
rect 144696 41352 144702 41364
rect 530720 40892 530748 41432
rect 530832 40960 530860 42432
rect 530900 41028 530928 42500
rect 530968 41096 530996 42568
rect 675018 41096 675024 41108
rect 530968 41068 675024 41096
rect 675018 41056 675024 41068
rect 675076 41056 675082 41108
rect 674926 41028 674932 41040
rect 530900 41000 674932 41028
rect 674926 40988 674932 41000
rect 674984 40988 674990 41040
rect 675110 40960 675116 40972
rect 530832 40932 675116 40960
rect 675110 40920 675116 40932
rect 675168 40920 675174 40972
rect 572714 40892 572720 40904
rect 530720 40864 572720 40892
rect 572714 40852 572720 40864
rect 572772 40852 572778 40904
rect 572714 40672 572720 40724
rect 572772 40712 572778 40724
rect 674834 40712 674840 40724
rect 572772 40684 674840 40712
rect 572772 40672 572778 40684
rect 674834 40672 674840 40684
rect 674892 40672 674898 40724
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143074 40100 143080 40112
rect 141048 40072 143080 40100
rect 141048 40060 141054 40072
rect 142586 39950 142614 40072
rect 143074 40060 143080 40072
rect 143132 40060 143138 40112
<< via1 >>
rect 284668 995256 284720 995308
rect 288992 995256 289044 995308
rect 538128 995256 538180 995308
rect 539876 995256 539928 995308
rect 130292 995188 130344 995240
rect 134616 995188 134668 995240
rect 526904 995188 526956 995240
rect 531228 995188 531280 995240
rect 78864 994856 78916 994908
rect 83188 994856 83240 994908
rect 83280 994856 83332 994908
rect 133972 994856 134024 994908
rect 135168 994856 135220 994908
rect 135260 994856 135312 994908
rect 143264 994984 143316 995036
rect 186688 994856 186740 994908
rect 194692 994856 194744 994908
rect 233700 994856 233752 994908
rect 237472 994856 237524 994908
rect 79508 994788 79560 994840
rect 130936 994788 130988 994840
rect 182364 994788 182416 994840
rect 183468 994788 183520 994840
rect 185400 994788 185452 994840
rect 236736 994788 236788 994840
rect 288348 994856 288400 994908
rect 289636 994856 289688 994908
rect 297640 994856 297692 994908
rect 89996 994720 90048 994772
rect 141424 994720 141476 994772
rect 192852 994720 192904 994772
rect 244188 994720 244240 994772
rect 295800 994788 295852 994840
rect 391480 994856 391532 994908
rect 399484 994856 399536 994908
rect 480444 994856 480496 994908
rect 488448 994856 488500 994908
rect 531872 994856 531924 994908
rect 538128 994856 538180 994908
rect 633624 994856 633676 994908
rect 641628 994856 641680 994908
rect 397644 994788 397696 994840
rect 486608 994788 486660 994840
rect 538036 994788 538088 994840
rect 639788 994788 639840 994840
rect 288624 994720 288676 994772
rect 288992 994720 289044 994772
rect 386512 994720 386564 994772
rect 390652 994720 390704 994772
rect 83188 994652 83240 994704
rect 130292 994652 130344 994704
rect 181720 994652 181772 994704
rect 186044 994652 186096 994704
rect 233056 994652 233108 994704
rect 237380 994652 237432 994704
rect 237472 994652 237524 994704
rect 285312 994652 285364 994704
rect 333244 994652 333296 994704
rect 387156 994652 387208 994704
rect 476120 994720 476172 994772
rect 527548 994720 527600 994772
rect 528284 994720 528336 994772
rect 531228 994720 531280 994772
rect 632336 994720 632388 994772
rect 390928 994652 390980 994704
rect 475476 994652 475528 994704
rect 479800 994652 479852 994704
rect 526904 994652 526956 994704
rect 628656 994652 628708 994704
rect 632980 994652 633032 994704
rect 83832 994584 83884 994636
rect 91836 994584 91888 994636
rect 183468 994584 183520 994636
rect 233700 994584 233752 994636
rect 288624 994584 288676 994636
rect 135168 994516 135220 994568
rect 185400 994516 185452 994568
rect 238024 994516 238076 994568
rect 246028 994516 246080 994568
rect 288348 994516 288400 994568
rect 390192 994584 390244 994636
rect 479156 994584 479208 994636
rect 528284 994584 528336 994636
rect 629300 994584 629352 994636
rect 530584 994516 530636 994568
rect 531228 994516 531280 994568
rect 43628 994380 43680 994432
rect 78864 994380 78916 994432
rect 639788 994380 639840 994432
rect 674196 994380 674248 994432
rect 43444 994312 43496 994364
rect 79508 994312 79560 994364
rect 632336 994312 632388 994364
rect 674288 994312 674340 994364
rect 43536 994244 43588 994296
rect 82544 994244 82596 994296
rect 83280 994244 83332 994296
rect 632980 994244 633032 994296
rect 674380 994244 674432 994296
rect 42340 994176 42392 994228
rect 89996 994176 90048 994228
rect 629300 994176 629352 994228
rect 675116 994176 675168 994228
rect 580540 994088 580592 994140
rect 674104 994088 674156 994140
rect 41788 967920 41840 967972
rect 42432 967920 42484 967972
rect 674380 967376 674432 967428
rect 675208 967376 675260 967428
rect 675208 965268 675260 965320
rect 675392 965268 675444 965320
rect 674288 964112 674340 964164
rect 675300 964112 675352 964164
rect 41788 961324 41840 961376
rect 42340 961324 42392 961376
rect 43628 961324 43680 961376
rect 674932 960644 674984 960696
rect 675392 960644 675444 960696
rect 675208 960168 675260 960220
rect 675208 959964 675260 960016
rect 42248 959012 42300 959064
rect 42616 959012 42668 959064
rect 43536 959012 43588 959064
rect 41788 957652 41840 957704
rect 43444 957652 43496 957704
rect 42432 957448 42484 957500
rect 42432 957244 42484 957296
rect 674196 953300 674248 953352
rect 675116 953300 675168 953352
rect 675576 953300 675628 953352
rect 675024 875780 675076 875832
rect 675392 875780 675444 875832
rect 674840 874488 674892 874540
rect 675208 874488 675260 874540
rect 675392 874488 675444 874540
rect 675024 871632 675076 871684
rect 675392 871632 675444 871684
rect 674932 864084 674984 864136
rect 675116 864084 675168 864136
rect 675392 864084 675444 864136
rect 675300 818320 675352 818372
rect 677508 818320 677560 818372
rect 41788 799552 41840 799604
rect 42340 799552 42392 799604
rect 41788 797716 41840 797768
rect 42432 797716 42484 797768
rect 42616 797716 42668 797768
rect 41788 792548 41840 792600
rect 42340 792548 42392 792600
rect 41788 791936 41840 791988
rect 42524 791936 42576 791988
rect 41788 787244 41840 787296
rect 42524 787244 42576 787296
rect 41788 786632 41840 786684
rect 42340 786632 42392 786684
rect 675208 786564 675260 786616
rect 675392 786564 675444 786616
rect 674840 785272 674892 785324
rect 675392 785272 675444 785324
rect 675024 783232 675076 783284
rect 675392 783232 675444 783284
rect 675208 782688 675260 782740
rect 675392 782688 675444 782740
rect 675208 780988 675260 781040
rect 675392 780988 675444 781040
rect 674932 775004 674984 775056
rect 675392 775004 675444 775056
rect 675208 773984 675260 774036
rect 675392 773984 675444 774036
rect 41788 756372 41840 756424
rect 42708 756372 42760 756424
rect 41788 755352 41840 755404
rect 42432 755352 42484 755404
rect 42616 755352 42668 755404
rect 41788 749368 41840 749420
rect 42708 749368 42760 749420
rect 41788 747668 41840 747720
rect 42340 747668 42392 747720
rect 41788 745084 41840 745136
rect 42524 745084 42576 745136
rect 41788 743792 41840 743844
rect 42340 743792 42392 743844
rect 675116 741004 675168 741056
rect 675576 741004 675628 741056
rect 674840 740324 674892 740376
rect 675208 740324 675260 740376
rect 675392 740324 675444 740376
rect 675024 737264 675076 737316
rect 675392 737264 675444 737316
rect 675116 736992 675168 737044
rect 675392 736992 675444 737044
rect 674840 735972 674892 736024
rect 675392 735972 675444 736024
rect 674932 729920 674984 729972
rect 675392 729920 675444 729972
rect 674840 729036 674892 729088
rect 675392 729036 675444 729088
rect 675300 726656 675352 726708
rect 674932 726452 674984 726504
rect 675208 726452 675260 726504
rect 675300 726452 675352 726504
rect 41788 713124 41840 713176
rect 42432 713124 42484 713176
rect 41788 711696 41840 711748
rect 42616 711696 42668 711748
rect 41788 706188 41840 706240
rect 42432 706188 42484 706240
rect 42340 705780 42392 705832
rect 41788 705508 41840 705560
rect 42340 705508 42392 705560
rect 42248 705168 42300 705220
rect 41788 704896 41840 704948
rect 42524 704896 42576 704948
rect 41788 700816 41840 700868
rect 42708 700816 42760 700868
rect 42248 700476 42300 700528
rect 674932 698980 674984 699032
rect 675392 698980 675444 699032
rect 674932 696192 674984 696244
rect 674932 695988 674984 696040
rect 675024 695920 675076 695972
rect 675392 695920 675444 695972
rect 674932 695308 674984 695360
rect 675392 695308 675444 695360
rect 674840 693200 674892 693252
rect 675392 693200 675444 693252
rect 675024 692044 675076 692096
rect 675392 692044 675444 692096
rect 675208 691636 675260 691688
rect 675392 691636 675444 691688
rect 675300 691568 675352 691620
rect 675300 691364 675352 691416
rect 675116 685176 675168 685228
rect 675392 685176 675444 685228
rect 675208 684020 675260 684072
rect 675392 684020 675444 684072
rect 675116 674160 675168 674212
rect 675116 673956 675168 674008
rect 675024 671372 675076 671424
rect 675208 671372 675260 671424
rect 41788 669944 41840 669996
rect 42432 669944 42484 669996
rect 41788 668516 41840 668568
rect 42616 668516 42668 668568
rect 42432 663076 42484 663128
rect 41788 663008 41840 663060
rect 42248 663008 42300 663060
rect 42432 662804 42484 662856
rect 41788 660764 41840 660816
rect 42432 660764 42484 660816
rect 41788 658656 41840 658708
rect 42340 658656 42392 658708
rect 42708 658656 42760 658708
rect 675116 651380 675168 651432
rect 675392 651380 675444 651432
rect 674932 650088 674984 650140
rect 675392 650088 675444 650140
rect 674840 647980 674892 648032
rect 675392 647980 675444 648032
rect 675116 647436 675168 647488
rect 675392 647436 675444 647488
rect 675208 645736 675260 645788
rect 675392 645736 675444 645788
rect 675024 639752 675076 639804
rect 675392 639752 675444 639804
rect 675208 638800 675260 638852
rect 675392 638800 675444 638852
rect 41972 625064 42024 625116
rect 42616 625064 42668 625116
rect 41788 618468 41840 618520
rect 42432 618468 42484 618520
rect 42248 614932 42300 614984
rect 42708 614932 42760 614984
rect 41788 613844 41840 613896
rect 42340 613844 42392 613896
rect 42524 605820 42576 605872
rect 42708 605820 42760 605872
rect 675116 605752 675168 605804
rect 675576 605752 675628 605804
rect 674932 605480 674984 605532
rect 675392 605480 675444 605532
rect 674840 602352 674892 602404
rect 674932 602080 674984 602132
rect 675392 602080 675444 602132
rect 675116 601808 675168 601860
rect 675392 601808 675444 601860
rect 675208 600788 675260 600840
rect 675392 600788 675444 600840
rect 675024 594668 675076 594720
rect 675392 594668 675444 594720
rect 675208 593784 675260 593836
rect 675392 593784 675444 593836
rect 41788 583516 41840 583568
rect 42432 583516 42484 583568
rect 41788 581816 41840 581868
rect 42524 581816 42576 581868
rect 41788 576444 41840 576496
rect 42432 576444 42484 576496
rect 42248 576240 42300 576292
rect 42708 576240 42760 576292
rect 41788 574336 41840 574388
rect 42432 574336 42484 574388
rect 42616 574336 42668 574388
rect 41788 571616 41840 571668
rect 42616 571616 42668 571668
rect 675116 561484 675168 561536
rect 675392 561484 675444 561536
rect 674840 560940 674892 560992
rect 675392 560940 675444 560992
rect 674932 557812 674984 557864
rect 675392 557812 675444 557864
rect 675116 557132 675168 557184
rect 675392 557132 675444 557184
rect 675208 555568 675260 555620
rect 675392 555568 675444 555620
rect 675024 550468 675076 550520
rect 675392 550468 675444 550520
rect 41788 539112 41840 539164
rect 42524 539112 42576 539164
rect 41788 532108 41840 532160
rect 42432 532108 42484 532160
rect 41972 528436 42024 528488
rect 42708 528436 42760 528488
rect 675300 503888 675352 503940
rect 677428 503888 677480 503940
rect 674104 427796 674156 427848
rect 677448 427796 677500 427848
rect 41788 412904 41840 412956
rect 42340 412904 42392 412956
rect 41788 410932 41840 410984
rect 42616 410932 42668 410984
rect 41788 405764 41840 405816
rect 42340 405764 42392 405816
rect 41788 404472 41840 404524
rect 42432 404472 42484 404524
rect 41788 400392 41840 400444
rect 42432 400392 42484 400444
rect 42708 400392 42760 400444
rect 674840 383732 674892 383784
rect 675392 383732 675444 383784
rect 675024 379788 675076 379840
rect 675392 379788 675444 379840
rect 674840 378360 674892 378412
rect 675392 378360 675444 378412
rect 674840 371424 674892 371476
rect 675392 371424 675444 371476
rect 41788 369520 41840 369572
rect 42340 369520 42392 369572
rect 41788 368636 41840 368688
rect 42616 368636 42668 368688
rect 41788 362584 41840 362636
rect 42340 362584 42392 362636
rect 41788 360340 41840 360392
rect 42524 360340 42576 360392
rect 42708 360340 42760 360392
rect 41788 357212 41840 357264
rect 42432 357212 42484 357264
rect 42248 357008 42300 357060
rect 675116 338784 675168 338836
rect 675392 338784 675444 338836
rect 674932 337492 674984 337544
rect 675392 337492 675444 337544
rect 675024 335384 675076 335436
rect 675208 335384 675260 335436
rect 675392 335384 675444 335436
rect 675024 334228 675076 334280
rect 675392 334228 675444 334280
rect 674840 328040 674892 328092
rect 675116 328040 675168 328092
rect 675392 328040 675444 328092
rect 41788 326340 41840 326392
rect 42432 326340 42484 326392
rect 41788 325116 41840 325168
rect 42524 325116 42576 325168
rect 41788 319404 41840 319456
rect 42432 319404 42484 319456
rect 41788 318724 41840 318776
rect 42340 318724 42392 318776
rect 41788 318112 41840 318164
rect 42708 318112 42760 318164
rect 41788 313488 41840 313540
rect 42340 313488 42392 313540
rect 675024 294108 675076 294160
rect 675392 294108 675444 294160
rect 674932 293224 674984 293276
rect 675392 293224 675444 293276
rect 674932 289484 674984 289536
rect 675116 289484 675168 289536
rect 675392 289484 675444 289536
rect 675024 288600 675076 288652
rect 675300 288600 675352 288652
rect 41788 283160 41840 283212
rect 42432 283160 42484 283212
rect 674840 282276 674892 282328
rect 675392 282276 675444 282328
rect 41788 282072 41840 282124
rect 42524 282072 42576 282124
rect 675208 281188 675260 281240
rect 675392 281188 675444 281240
rect 41788 276156 41840 276208
rect 42432 276156 42484 276208
rect 41788 274524 41840 274576
rect 42340 274524 42392 274576
rect 41788 273912 41840 273964
rect 42616 273912 42668 273964
rect 41788 270580 41840 270632
rect 42340 270580 42392 270632
rect 675116 248752 675168 248804
rect 675392 248752 675444 248804
rect 675024 247460 675076 247512
rect 675392 247460 675444 247512
rect 674932 244468 674984 244520
rect 675392 244468 675444 244520
rect 41788 239912 41840 239964
rect 42432 239912 42484 239964
rect 41788 238484 41840 238536
rect 42524 238484 42576 238536
rect 674840 237668 674892 237720
rect 675392 237668 675444 237720
rect 675208 236240 675260 236292
rect 675392 236240 675444 236292
rect 41788 232976 41840 233028
rect 42432 232976 42484 233028
rect 41788 232364 41840 232416
rect 42340 232364 42392 232416
rect 41788 231684 41840 231736
rect 42616 231684 42668 231736
rect 41788 227060 41840 227112
rect 42340 227060 42392 227112
rect 675116 203464 675168 203516
rect 675300 203464 675352 203516
rect 675024 202308 675076 202360
rect 675392 202308 675444 202360
rect 674932 200200 674984 200252
rect 675392 200200 675444 200252
rect 675208 199248 675260 199300
rect 675208 199044 675260 199096
rect 41788 196732 41840 196784
rect 42708 196732 42760 196784
rect 41788 195304 41840 195356
rect 42432 195304 42484 195356
rect 675208 191904 675260 191956
rect 675392 191904 675444 191956
rect 41788 189796 41840 189848
rect 42708 189796 42760 189848
rect 41788 188096 41840 188148
rect 42340 188096 42392 188148
rect 41788 187552 41840 187604
rect 42524 187552 42576 187604
rect 41788 184152 41840 184204
rect 42340 184152 42392 184204
rect 675300 158720 675352 158772
rect 675116 158516 675168 158568
rect 674840 157292 674892 157344
rect 675024 157292 675076 157344
rect 675392 157292 675444 157344
rect 674932 155184 674984 155236
rect 675392 155184 675444 155236
rect 675024 147092 675076 147144
rect 675208 147092 675260 147144
rect 675392 147092 675444 147144
rect 675024 113092 675076 113144
rect 675392 113092 675444 113144
rect 674840 112480 674892 112532
rect 675392 112480 675444 112532
rect 674932 109080 674984 109132
rect 675392 109080 675444 109132
rect 675024 108808 675076 108860
rect 675392 108808 675444 108860
rect 675208 107788 675260 107840
rect 675392 107788 675444 107840
rect 675208 102008 675260 102060
rect 675300 101804 675352 101856
rect 527456 43156 527508 43208
rect 523776 43088 523828 43140
rect 516140 43020 516192 43072
rect 459652 42952 459704 43004
rect 467656 42952 467708 43004
rect 415308 42884 415360 42936
rect 467840 42884 467892 42936
rect 473268 42884 473320 42936
rect 526812 42884 526864 42936
rect 411076 42816 411128 42868
rect 419724 42816 419776 42868
rect 42156 42428 42208 42480
rect 147680 42428 147732 42480
rect 42064 42360 42116 42412
rect 195980 42720 196032 42772
rect 295248 42748 295300 42800
rect 303252 42748 303304 42800
rect 350080 42748 350132 42800
rect 358084 42748 358136 42800
rect 360568 42748 360620 42800
rect 406752 42748 406804 42800
rect 461492 42816 461544 42868
rect 516140 42816 516192 42868
rect 467840 42748 467892 42800
rect 468944 42748 468996 42800
rect 523776 42748 523828 42800
rect 88800 42252 88852 42304
rect 199016 42612 199068 42664
rect 307576 42680 307628 42732
rect 362408 42680 362460 42732
rect 417240 42680 417292 42732
rect 471980 42680 472032 42732
rect 473268 42680 473320 42732
rect 514484 42680 514536 42732
rect 522488 42680 522540 42732
rect 200856 42612 200908 42664
rect 241336 42612 241388 42664
rect 297732 42612 297784 42664
rect 300768 42612 300820 42664
rect 305092 42612 305144 42664
rect 309416 42612 309468 42664
rect 352564 42612 352616 42664
rect 355600 42612 355652 42664
rect 359924 42612 359976 42664
rect 364248 42612 364300 42664
rect 407396 42612 407448 42664
rect 410432 42612 410484 42664
rect 416044 42612 416096 42664
rect 419080 42612 419132 42664
rect 462136 42612 462188 42664
rect 465172 42612 465224 42664
rect 470784 42612 470836 42664
rect 473820 42612 473872 42664
rect 516968 42612 517020 42664
rect 520004 42612 520056 42664
rect 188528 42544 188580 42596
rect 192852 42544 192904 42596
rect 201500 42544 201552 42596
rect 297088 42544 297140 42596
rect 299572 42544 299624 42596
rect 305736 42544 305788 42596
rect 351920 42544 351972 42596
rect 354404 42544 354456 42596
rect 360568 42544 360620 42596
rect 404912 42544 404964 42596
rect 412916 42544 412968 42596
rect 413560 42544 413612 42596
rect 417884 42544 417936 42596
rect 468300 42544 468352 42596
rect 472624 42544 472676 42596
rect 523132 42544 523184 42596
rect 527456 42544 527508 42596
rect 199660 42476 199712 42528
rect 303896 42476 303948 42528
rect 308220 42476 308272 42528
rect 358728 42476 358780 42528
rect 363052 42476 363104 42528
rect 465816 42476 465868 42528
rect 474464 42476 474516 42528
rect 42248 42100 42300 42152
rect 140964 42100 141016 42152
rect 42340 42032 42392 42084
rect 145104 42032 145156 42084
rect 147680 42048 147732 42100
rect 188528 42408 188580 42460
rect 195980 42408 196032 42460
rect 304540 42408 304592 42460
rect 359372 42408 359424 42460
rect 414204 42408 414256 42460
rect 415308 42408 415360 42460
rect 186688 42340 186740 42392
rect 194692 42340 194744 42392
rect 409236 42340 409288 42392
rect 412272 42340 412324 42392
rect 415400 42340 415452 42392
rect 518808 42340 518860 42392
rect 524972 42340 525024 42392
rect 198464 41896 198516 41948
rect 200120 41896 200172 41948
rect 186136 41828 186188 41880
rect 195244 41828 195296 41880
rect 199568 41828 199620 41880
rect 189264 41760 189316 41812
rect 191104 41760 191156 41812
rect 192300 41760 192352 41812
rect 193588 41760 193640 41812
rect 196440 41760 196492 41812
rect 143080 41420 143132 41472
rect 145104 41420 145156 41472
rect 186136 41420 186188 41472
rect 144644 41352 144696 41404
rect 469680 41964 469732 42016
rect 470692 41964 470744 42016
rect 305276 41896 305328 41948
rect 306288 41896 306340 41948
rect 308680 41896 308732 41948
rect 464160 41828 464212 41880
rect 467196 41828 467248 41880
rect 470048 41828 470100 41880
rect 360016 41760 360068 41812
rect 361120 41760 361172 41812
rect 363512 41760 363564 41812
rect 410524 41760 410576 41812
rect 411536 41760 411588 41812
rect 414848 41760 414900 41812
rect 415860 41760 415912 41812
rect 465356 41760 465408 41812
rect 466368 41760 466420 41812
rect 469404 41760 469456 41812
rect 520096 41760 520148 41812
rect 521200 41760 521252 41812
rect 524236 41760 524288 41812
rect 525524 41760 525576 41812
rect 527916 41760 527968 41812
rect 675024 41056 675076 41108
rect 674932 40988 674984 41040
rect 675116 40920 675168 40972
rect 572720 40852 572772 40904
rect 572720 40672 572772 40724
rect 674840 40672 674892 40724
rect 140996 40060 141048 40112
rect 143080 40060 143132 40112
<< metal2 >>
rect 333242 997928 333298 997937
rect 333242 997863 333298 997872
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 78876 994914 78904 995452
rect 78864 994908 78916 994914
rect 78864 994850 78916 994856
rect 78876 994438 78904 994850
rect 79520 994846 79548 995452
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 79508 994840 79560 994846
rect 79508 994782 79560 994788
rect 43628 994432 43680 994438
rect 43628 994374 43680 994380
rect 78864 994432 78916 994438
rect 78864 994374 78916 994380
rect 43444 994364 43496 994370
rect 43444 994306 43496 994312
rect 42340 994228 42392 994234
rect 42340 994170 42392 994176
rect 42352 982574 42380 994170
rect 42352 982546 42472 982574
rect 41722 969870 41920 969898
rect 41892 969354 41920 969870
rect 41892 969326 42288 969354
rect 41713 969217 42193 969273
rect 41722 968035 41828 968063
rect 41800 967978 41828 968035
rect 41788 967972 41840 967978
rect 41788 967914 41840 967920
rect 41713 967377 42193 967433
rect 41713 966733 42193 966789
rect 41713 965537 42193 965593
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 41713 963053 42193 963109
rect 41713 962501 42193 962557
rect 42260 962010 42288 969326
rect 42444 967978 42472 982546
rect 42432 967972 42484 967978
rect 42432 967914 42484 967920
rect 41800 961982 42288 962010
rect 41800 961894 41828 961982
rect 41722 961866 41828 961894
rect 41788 961376 41840 961382
rect 41788 961318 41840 961324
rect 42340 961376 42392 961382
rect 42340 961318 42392 961324
rect 41800 961255 41828 961318
rect 41722 961227 41828 961255
rect 41722 960583 41920 960611
rect 41892 960514 41920 960583
rect 41892 960486 42288 960514
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 42260 959070 42288 960486
rect 42248 959064 42300 959070
rect 42248 959006 42300 959012
rect 41713 958729 42193 958785
rect 41713 958177 42193 958233
rect 41788 957704 41840 957710
rect 41788 957646 41840 957652
rect 41800 957575 41828 957646
rect 41722 957547 41828 957575
rect 42352 957386 42380 961318
rect 42444 957506 42472 967914
rect 42616 959064 42668 959070
rect 42616 959006 42668 959012
rect 42432 957500 42484 957506
rect 42432 957442 42484 957448
rect 41800 957358 42564 957386
rect 41800 956931 41828 957358
rect 42432 957296 42484 957302
rect 42432 957238 42484 957244
rect 41722 956903 41828 956931
rect 41713 956337 42193 956393
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 41418 881920 41474 881929
rect 41418 881855 41474 881864
rect 41432 880025 41460 881855
rect 41418 880016 41474 880025
rect 41418 879951 41474 879960
rect 42246 880016 42302 880025
rect 42246 879951 42302 879960
rect 41722 800075 41828 800103
rect 41800 799610 41828 800075
rect 41788 799604 41840 799610
rect 41788 799546 41840 799552
rect 41713 799417 42193 799473
rect 41722 798238 41828 798266
rect 41800 797774 41828 798238
rect 41788 797768 41840 797774
rect 41788 797710 41840 797716
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41788 792600 41840 792606
rect 41788 792542 41840 792548
rect 41800 792099 41828 792542
rect 41722 792071 41828 792099
rect 41788 791988 41840 791994
rect 41788 791930 41840 791936
rect 41800 791466 41828 791930
rect 41722 791438 41828 791466
rect 42260 790922 42288 879951
rect 42340 799604 42392 799610
rect 42340 799546 42392 799552
rect 42352 792606 42380 799546
rect 42444 797774 42472 957238
rect 42432 797768 42484 797774
rect 42432 797710 42484 797716
rect 42340 792600 42392 792606
rect 42340 792542 42392 792548
rect 42536 791994 42564 957358
rect 42628 881929 42656 959006
rect 43456 957710 43484 994306
rect 43536 994296 43588 994302
rect 43536 994238 43588 994244
rect 43548 959070 43576 994238
rect 43640 961382 43668 994374
rect 79520 994370 79548 994782
rect 79508 994364 79560 994370
rect 79508 994306 79560 994312
rect 82556 994302 82584 995452
rect 83200 994914 83228 995452
rect 83188 994908 83240 994914
rect 83188 994850 83240 994856
rect 83280 994908 83332 994914
rect 83280 994850 83332 994856
rect 83200 994710 83228 994850
rect 83188 994704 83240 994710
rect 83188 994646 83240 994652
rect 83292 994302 83320 994850
rect 83844 994642 83872 995452
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 90008 994778 90036 995452
rect 91217 995407 91273 995887
rect 89996 994772 90048 994778
rect 89996 994714 90048 994720
rect 83832 994636 83884 994642
rect 83832 994578 83884 994584
rect 82544 994296 82596 994302
rect 82544 994238 82596 994244
rect 83280 994296 83332 994302
rect 83280 994238 83332 994244
rect 90008 994234 90036 994714
rect 91848 994642 91876 995452
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 130304 995246 130332 995452
rect 130292 995240 130344 995246
rect 130292 995182 130344 995188
rect 130304 994710 130332 995182
rect 130948 994846 130976 995452
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 133984 994914 134012 995452
rect 134628 995246 134656 995452
rect 134616 995240 134668 995246
rect 134616 995182 134668 995188
rect 135272 994914 135300 995452
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 133972 994908 134024 994914
rect 133972 994850 134024 994856
rect 135168 994908 135220 994914
rect 135168 994850 135220 994856
rect 135260 994908 135312 994914
rect 135260 994850 135312 994856
rect 130936 994840 130988 994846
rect 130936 994782 130988 994788
rect 130292 994704 130344 994710
rect 130292 994646 130344 994652
rect 91836 994636 91888 994642
rect 91836 994578 91888 994584
rect 135180 994574 135208 994850
rect 141436 994778 141464 995452
rect 142617 995407 142673 995887
rect 143276 995042 143304 995452
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 181717 995438 181760 995466
rect 182361 995438 182404 995466
rect 143264 995036 143316 995042
rect 143264 994978 143316 994984
rect 141424 994772 141476 994778
rect 141424 994714 141476 994720
rect 181732 994710 181760 995438
rect 182376 994846 182404 995438
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 185397 995438 185440 995466
rect 186041 995438 186084 995466
rect 186685 995438 186728 995466
rect 185412 994846 185440 995438
rect 182364 994840 182416 994846
rect 182364 994782 182416 994788
rect 183468 994840 183520 994846
rect 183468 994782 183520 994788
rect 185400 994840 185452 994846
rect 185400 994782 185452 994788
rect 181720 994704 181772 994710
rect 181720 994646 181772 994652
rect 183480 994642 183508 994782
rect 183468 994636 183520 994642
rect 183468 994578 183520 994584
rect 185412 994574 185440 994782
rect 186056 994710 186084 995438
rect 186700 994914 186728 995438
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 192849 995438 192892 995466
rect 186688 994908 186740 994914
rect 186688 994850 186740 994856
rect 192864 994778 192892 995438
rect 194017 995407 194073 995887
rect 194689 995438 194732 995466
rect 194704 994914 194732 995438
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 233068 995438 233117 995466
rect 233712 995438 233761 995466
rect 194692 994908 194744 994914
rect 194692 994850 194744 994856
rect 192852 994772 192904 994778
rect 192852 994714 192904 994720
rect 233068 994710 233096 995438
rect 233712 994914 233740 995438
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 236748 995438 236797 995466
rect 237392 995438 237441 995466
rect 238036 995438 238085 995466
rect 233700 994908 233752 994914
rect 233700 994850 233752 994856
rect 186044 994704 186096 994710
rect 186044 994646 186096 994652
rect 233056 994704 233108 994710
rect 233056 994646 233108 994652
rect 233712 994642 233740 994850
rect 236748 994846 236776 995438
rect 236736 994840 236788 994846
rect 236736 994782 236788 994788
rect 237392 994710 237420 995438
rect 237472 994908 237524 994914
rect 237472 994850 237524 994856
rect 237484 994710 237512 994850
rect 237380 994704 237432 994710
rect 237380 994646 237432 994652
rect 237472 994704 237524 994710
rect 237472 994646 237524 994652
rect 233700 994636 233752 994642
rect 233700 994578 233752 994584
rect 238036 994574 238064 995438
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 244200 995438 244249 995466
rect 244200 994778 244228 995438
rect 245417 995407 245473 995887
rect 246040 995438 246089 995466
rect 244188 994772 244240 994778
rect 244188 994714 244240 994720
rect 246040 994574 246068 995438
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 284680 995314 284708 995452
rect 284668 995308 284720 995314
rect 284668 995250 284720 995256
rect 285324 994710 285352 995452
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 288360 994914 288388 995452
rect 289004 995314 289032 995452
rect 288992 995308 289044 995314
rect 288992 995250 289044 995256
rect 288348 994908 288400 994914
rect 288348 994850 288400 994856
rect 285312 994704 285364 994710
rect 285312 994646 285364 994652
rect 288360 994574 288388 994850
rect 289004 994778 289032 995250
rect 289648 994914 289676 995452
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 289636 994908 289688 994914
rect 289636 994850 289688 994856
rect 295812 994846 295840 995452
rect 297017 995407 297073 995887
rect 297652 994914 297680 995452
rect 297640 994908 297692 994914
rect 297640 994850 297692 994856
rect 295800 994840 295852 994846
rect 295800 994782 295852 994788
rect 288624 994772 288676 994778
rect 288624 994714 288676 994720
rect 288992 994772 289044 994778
rect 288992 994714 289044 994720
rect 288636 994642 288664 994714
rect 333256 994710 333284 997863
rect 580630 997858 580686 997867
rect 580630 997793 580686 997802
rect 580644 996234 580672 997793
rect 580552 996206 580672 996234
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 386524 994778 386552 995452
rect 386512 994772 386564 994778
rect 386512 994714 386564 994720
rect 387168 994710 387196 995452
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 333244 994704 333296 994710
rect 333244 994646 333296 994652
rect 387156 994704 387208 994710
rect 387156 994646 387208 994652
rect 390204 994642 390232 995452
rect 390664 995438 390862 995466
rect 390664 994778 390692 995438
rect 391492 994914 391520 995452
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 391480 994908 391532 994914
rect 391480 994850 391532 994856
rect 397656 994846 397684 995452
rect 398817 995407 398873 995887
rect 399496 994914 399524 995452
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 399484 994908 399536 994914
rect 399484 994850 399536 994856
rect 397644 994840 397696 994846
rect 397644 994782 397696 994788
rect 390652 994772 390704 994778
rect 390704 994720 390968 994726
rect 390652 994714 390968 994720
rect 390664 994710 390968 994714
rect 475488 994710 475516 995452
rect 476132 994778 476160 995452
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 476120 994772 476172 994778
rect 476120 994714 476172 994720
rect 390664 994704 390980 994710
rect 390664 994698 390928 994704
rect 390928 994646 390980 994652
rect 475476 994704 475528 994710
rect 475476 994646 475528 994652
rect 479168 994642 479196 995452
rect 479812 994710 479840 995452
rect 480456 994914 480484 995452
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 480444 994908 480496 994914
rect 480444 994850 480496 994856
rect 486620 994846 486648 995452
rect 487817 995407 487873 995887
rect 488460 994914 488488 995452
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 526916 995246 526944 995452
rect 526904 995240 526956 995246
rect 526904 995182 526956 995188
rect 488448 994908 488500 994914
rect 488448 994850 488500 994856
rect 486608 994840 486660 994846
rect 486608 994782 486660 994788
rect 526916 994710 526944 995182
rect 527560 994778 527588 995452
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 527548 994772 527600 994778
rect 527548 994714 527600 994720
rect 528284 994772 528336 994778
rect 528284 994714 528336 994720
rect 479800 994704 479852 994710
rect 479800 994646 479852 994652
rect 526904 994704 526956 994710
rect 526904 994646 526956 994652
rect 528296 994642 528324 994714
rect 288624 994636 288676 994642
rect 288624 994578 288676 994584
rect 390192 994636 390244 994642
rect 390192 994578 390244 994584
rect 479156 994636 479208 994642
rect 479156 994578 479208 994584
rect 528284 994636 528336 994642
rect 528284 994578 528336 994584
rect 530596 994574 530624 995452
rect 531240 995246 531268 995452
rect 531228 995240 531280 995246
rect 531228 995182 531280 995188
rect 531884 994914 531912 995452
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 531872 994908 531924 994914
rect 531872 994850 531924 994856
rect 538048 994846 538076 995452
rect 539217 995407 539273 995887
rect 539888 995314 539916 995452
rect 538128 995308 538180 995314
rect 538128 995250 538180 995256
rect 539876 995308 539928 995314
rect 539876 995250 539928 995256
rect 538140 994914 538168 995250
rect 538128 994908 538180 994914
rect 538128 994850 538180 994856
rect 538036 994840 538088 994846
rect 538036 994782 538088 994788
rect 531228 994772 531280 994778
rect 531228 994714 531280 994720
rect 531240 994574 531268 994714
rect 135168 994568 135220 994574
rect 135168 994510 135220 994516
rect 185400 994568 185452 994574
rect 185400 994510 185452 994516
rect 238024 994568 238076 994574
rect 238024 994510 238076 994516
rect 246028 994568 246080 994574
rect 246028 994510 246080 994516
rect 288348 994568 288400 994574
rect 288348 994510 288400 994516
rect 530584 994568 530636 994574
rect 530584 994510 530636 994516
rect 531228 994568 531280 994574
rect 531228 994510 531280 994516
rect 89996 994228 90048 994234
rect 89996 994170 90048 994176
rect 580552 994146 580580 996206
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 628668 995438 628717 995466
rect 629312 995438 629361 995466
rect 628668 994710 628696 995438
rect 628656 994704 628708 994710
rect 628656 994646 628708 994652
rect 629312 994642 629340 995438
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 632348 995438 632397 995466
rect 632992 995438 633041 995466
rect 633636 995438 633685 995466
rect 632348 994778 632376 995438
rect 632336 994772 632388 994778
rect 632336 994714 632388 994720
rect 629300 994636 629352 994642
rect 629300 994578 629352 994584
rect 629312 994234 629340 994578
rect 632348 994370 632376 994714
rect 632992 994710 633020 995438
rect 633636 994914 633664 995438
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 639800 995438 639849 995466
rect 633624 994908 633676 994914
rect 633624 994850 633676 994856
rect 639800 994846 639828 995438
rect 641017 995407 641073 995887
rect 641640 995438 641689 995466
rect 641640 994914 641668 995438
rect 641628 994908 641680 994914
rect 641628 994850 641680 994856
rect 639788 994840 639840 994846
rect 639788 994782 639840 994788
rect 632980 994704 633032 994710
rect 632980 994646 633032 994652
rect 632336 994364 632388 994370
rect 632336 994306 632388 994312
rect 632992 994302 633020 994646
rect 639800 994438 639828 994782
rect 639788 994432 639840 994438
rect 639788 994374 639840 994380
rect 674196 994432 674248 994438
rect 674196 994374 674248 994380
rect 632980 994296 633032 994302
rect 632980 994238 633032 994244
rect 629300 994228 629352 994234
rect 629300 994170 629352 994176
rect 580540 994140 580592 994146
rect 580540 994082 580592 994088
rect 674104 994140 674156 994146
rect 674104 994082 674156 994088
rect 43628 961376 43680 961382
rect 43628 961318 43680 961324
rect 43536 959064 43588 959070
rect 43536 959006 43588 959012
rect 43444 957704 43496 957710
rect 43444 957646 43496 957652
rect 42614 881920 42670 881929
rect 42614 881855 42670 881864
rect 42616 797768 42668 797774
rect 42616 797710 42668 797716
rect 42524 791988 42576 791994
rect 42524 791930 42576 791936
rect 41892 790894 42288 790922
rect 41892 790806 41920 790894
rect 41722 790778 41920 790806
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 41722 787746 41828 787774
rect 41800 787302 41828 787746
rect 41788 787296 41840 787302
rect 41788 787238 41840 787244
rect 41722 787106 41828 787134
rect 41800 786690 41828 787106
rect 41788 786684 41840 786690
rect 41788 786626 41840 786632
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 41722 756894 41828 756922
rect 41800 756430 41828 756894
rect 41788 756424 41840 756430
rect 41788 756366 41840 756372
rect 41713 756217 42193 756273
rect 41788 755404 41840 755410
rect 41788 755346 41840 755352
rect 41800 755063 41828 755346
rect 41722 755035 41828 755063
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41788 749420 41840 749426
rect 41788 749362 41840 749368
rect 41800 748898 41828 749362
rect 41722 748870 41828 748898
rect 41722 748227 41828 748255
rect 41800 747726 41828 748227
rect 41788 747720 41840 747726
rect 41788 747662 41840 747668
rect 41722 747583 41828 747611
rect 41800 747130 41828 747583
rect 42260 747130 42288 790894
rect 42536 789374 42564 791930
rect 42352 789346 42564 789374
rect 42352 786690 42380 789346
rect 42524 787296 42576 787302
rect 42524 787238 42576 787244
rect 42340 786684 42392 786690
rect 42340 786626 42392 786632
rect 42352 747726 42380 786626
rect 42432 755404 42484 755410
rect 42432 755346 42484 755352
rect 42340 747720 42392 747726
rect 42340 747662 42392 747668
rect 41800 747102 42288 747130
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41788 745136 41840 745142
rect 41788 745078 41840 745084
rect 41800 744575 41828 745078
rect 41722 744547 41828 744575
rect 41722 743903 41828 743931
rect 41800 743850 41828 743903
rect 41788 743844 41840 743850
rect 41788 743786 41840 743792
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 41722 713675 41828 713703
rect 41800 713182 41828 713675
rect 41788 713176 41840 713182
rect 41788 713118 41840 713124
rect 41713 713017 42193 713073
rect 41722 711835 41828 711863
rect 41800 711754 41828 711835
rect 41788 711748 41840 711754
rect 41788 711690 41840 711696
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41788 706240 41840 706246
rect 41788 706182 41840 706188
rect 41800 705699 41828 706182
rect 41722 705671 41828 705699
rect 41788 705560 41840 705566
rect 41788 705502 41840 705508
rect 41800 705055 41828 705502
rect 42260 705226 42288 747102
rect 42352 743850 42380 747662
rect 42340 743844 42392 743850
rect 42340 743786 42392 743792
rect 42352 705838 42380 743786
rect 42444 731414 42472 755346
rect 42536 745142 42564 787238
rect 42628 755410 42656 797710
rect 42708 756424 42760 756430
rect 42708 756366 42760 756372
rect 42616 755404 42668 755410
rect 42616 755346 42668 755352
rect 42720 749426 42748 756366
rect 42708 749420 42760 749426
rect 42708 749362 42760 749368
rect 42524 745136 42576 745142
rect 42524 745078 42576 745084
rect 42536 741074 42564 745078
rect 42536 741046 42748 741074
rect 42444 731386 42656 731414
rect 42432 713176 42484 713182
rect 42432 713118 42484 713124
rect 42444 706246 42472 713118
rect 42628 711754 42656 731386
rect 42616 711748 42668 711754
rect 42616 711690 42668 711696
rect 42432 706240 42484 706246
rect 42432 706182 42484 706188
rect 42340 705832 42392 705838
rect 42340 705774 42392 705780
rect 42340 705560 42392 705566
rect 42340 705502 42392 705508
rect 42248 705220 42300 705226
rect 42248 705162 42300 705168
rect 41722 705027 41828 705055
rect 41788 704948 41840 704954
rect 41788 704890 41840 704896
rect 41800 704416 41828 704890
rect 41722 704388 41828 704416
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 42352 702434 42380 705502
rect 42524 704948 42576 704954
rect 42524 704890 42576 704896
rect 42260 702406 42380 702434
rect 41713 701977 42193 702033
rect 41722 701347 41828 701375
rect 41800 700874 41828 701347
rect 41788 700868 41840 700874
rect 41788 700810 41840 700816
rect 41722 700706 41828 700734
rect 41800 700618 41828 700706
rect 42260 700618 42288 702406
rect 41800 700590 42380 700618
rect 42248 700528 42300 700534
rect 42248 700470 42300 700476
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41722 670475 41828 670503
rect 41800 670002 41828 670475
rect 41788 669996 41840 670002
rect 41788 669938 41840 669944
rect 41713 669817 42193 669873
rect 41722 668630 41828 668658
rect 41800 668574 41828 668630
rect 41788 668568 41840 668574
rect 41788 668510 41840 668516
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 42260 663066 42288 700470
rect 41788 663060 41840 663066
rect 41788 663002 41840 663008
rect 42248 663060 42300 663066
rect 42248 663002 42300 663008
rect 41800 662499 41828 663002
rect 41722 662471 41828 662499
rect 41722 661830 41920 661858
rect 41892 661722 41920 661830
rect 42352 661722 42380 700590
rect 42432 669996 42484 670002
rect 42432 669938 42484 669944
rect 42444 663134 42472 669938
rect 42432 663128 42484 663134
rect 42432 663070 42484 663076
rect 42432 662856 42484 662862
rect 42432 662798 42484 662804
rect 41892 661694 42380 661722
rect 41722 661183 41828 661211
rect 41800 660822 41828 661183
rect 41788 660816 41840 660822
rect 41788 660758 41840 660764
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41788 658708 41840 658714
rect 41788 658650 41840 658656
rect 41800 658186 41828 658650
rect 41722 658158 41828 658186
rect 41722 657498 41828 657526
rect 41800 657370 41828 657498
rect 42260 657370 42288 661694
rect 42444 661042 42472 662798
rect 42352 661014 42472 661042
rect 42352 658714 42380 661014
rect 42536 660906 42564 704890
rect 42628 668574 42656 711690
rect 42720 700874 42748 741046
rect 42708 700868 42760 700874
rect 42708 700810 42760 700816
rect 42616 668568 42668 668574
rect 42616 668510 42668 668516
rect 42444 660878 42564 660906
rect 42444 660822 42472 660878
rect 42432 660816 42484 660822
rect 42432 660758 42484 660764
rect 42340 658708 42392 658714
rect 42340 658650 42392 658656
rect 41800 657342 42288 657370
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 42260 654134 42288 657342
rect 42260 654106 42380 654134
rect 41722 627286 41828 627314
rect 41800 627178 41828 627286
rect 41800 627150 42288 627178
rect 41713 626617 42193 626673
rect 41722 625435 42012 625463
rect 41984 625122 42012 625435
rect 41972 625116 42024 625122
rect 41972 625058 42024 625064
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 42260 619426 42288 627150
rect 41800 619398 42288 619426
rect 41800 619290 41828 619398
rect 41722 619262 41828 619290
rect 42352 619154 42380 654106
rect 41800 619126 42380 619154
rect 41800 618655 41828 619126
rect 41722 618627 41828 618655
rect 41788 618520 41840 618526
rect 41788 618462 41840 618468
rect 41800 618011 41828 618462
rect 41722 617983 41828 618011
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 42260 614990 42288 615021
rect 42248 614984 42300 614990
rect 42110 614940 42248 614968
rect 42248 614926 42300 614932
rect 42248 614925 42288 614926
rect 41722 614303 41828 614331
rect 41800 613902 41828 614303
rect 41788 613896 41840 613902
rect 41788 613838 41840 613844
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 41722 584075 41828 584103
rect 41800 583574 41828 584075
rect 41788 583568 41840 583574
rect 41788 583510 41840 583516
rect 41713 583417 42193 583473
rect 41722 582235 41828 582263
rect 41800 581874 41828 582235
rect 41788 581868 41840 581874
rect 41788 581810 41840 581816
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41788 576496 41840 576502
rect 41788 576438 41840 576444
rect 41800 576099 41828 576438
rect 42260 576298 42288 614925
rect 42352 613902 42380 619126
rect 42444 618526 42472 660758
rect 42628 625122 42656 668510
rect 42708 658708 42760 658714
rect 42708 658650 42760 658656
rect 42616 625116 42668 625122
rect 42616 625058 42668 625064
rect 42432 618520 42484 618526
rect 42432 618462 42484 618468
rect 42340 613896 42392 613902
rect 42340 613838 42392 613844
rect 42248 576292 42300 576298
rect 42248 576234 42300 576240
rect 42352 576099 42380 613838
rect 42444 610586 42472 618462
rect 42628 610858 42656 625058
rect 42720 614990 42748 658650
rect 42708 614984 42760 614990
rect 42708 614926 42760 614932
rect 42628 610830 42748 610858
rect 42444 610558 42656 610586
rect 42524 605872 42576 605878
rect 42524 605814 42576 605820
rect 42432 583568 42484 583574
rect 42432 583510 42484 583516
rect 42444 576502 42472 583510
rect 42536 581874 42564 605814
rect 42524 581868 42576 581874
rect 42524 581810 42576 581816
rect 42432 576496 42484 576502
rect 42432 576438 42484 576444
rect 41722 576071 41828 576099
rect 42260 576071 42380 576099
rect 41722 575427 41920 575455
rect 41892 575362 41920 575427
rect 42260 575362 42288 576071
rect 41892 575334 42288 575362
rect 41722 574790 41828 574818
rect 41800 574394 41828 574790
rect 41788 574388 41840 574394
rect 41788 574330 41840 574336
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41722 571747 41828 571775
rect 41800 571674 41828 571747
rect 41788 571668 41840 571674
rect 41788 571610 41840 571616
rect 41722 571098 41920 571126
rect 41892 571010 41920 571098
rect 42260 571010 42288 575334
rect 42432 574388 42484 574394
rect 42432 574330 42484 574336
rect 41892 570982 42288 571010
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 42260 557534 42288 570982
rect 42260 557506 42380 557534
rect 41722 540875 42288 540903
rect 41713 540217 42193 540273
rect 41788 539164 41840 539170
rect 41788 539106 41840 539112
rect 41800 539050 41828 539106
rect 41722 539022 41828 539050
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 42260 533338 42288 540875
rect 41800 533310 42288 533338
rect 41800 532899 41828 533310
rect 41722 532871 41828 532899
rect 42352 532794 42380 557506
rect 41800 532766 42380 532794
rect 41800 532250 41828 532766
rect 41722 532222 41828 532250
rect 41788 532160 41840 532166
rect 41788 532102 41840 532108
rect 41800 531611 41828 532102
rect 41722 531583 41828 531611
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41778 528546 42012 528574
rect 41984 528494 42012 528546
rect 41972 528488 42024 528494
rect 41972 528430 42024 528436
rect 41722 527903 41920 527931
rect 41892 527490 41920 527903
rect 42260 527490 42288 532766
rect 42444 532166 42472 574330
rect 42536 539170 42564 581810
rect 42628 574394 42656 610558
rect 42720 605878 42748 610830
rect 42708 605872 42760 605878
rect 42708 605814 42760 605820
rect 42708 576292 42760 576298
rect 42708 576234 42760 576240
rect 42616 574388 42668 574394
rect 42616 574330 42668 574336
rect 42720 574274 42748 576234
rect 42628 574246 42748 574274
rect 42628 571674 42656 574246
rect 42616 571668 42668 571674
rect 42616 571610 42668 571616
rect 42524 539164 42576 539170
rect 42524 539106 42576 539112
rect 42432 532160 42484 532166
rect 42432 532102 42484 532108
rect 41892 527462 42288 527490
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41722 413275 41828 413303
rect 41800 412962 41828 413275
rect 41788 412956 41840 412962
rect 41788 412898 41840 412904
rect 41713 412617 42193 412673
rect 41722 411434 41828 411462
rect 41800 410990 41828 411434
rect 41788 410984 41840 410990
rect 41788 410926 41840 410932
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 41788 405816 41840 405822
rect 41788 405758 41840 405764
rect 41800 405299 41828 405758
rect 41722 405271 41828 405299
rect 42260 404818 42288 527462
rect 42340 412956 42392 412962
rect 42340 412898 42392 412904
rect 42352 405822 42380 412898
rect 42340 405816 42392 405822
rect 42340 405758 42392 405764
rect 41892 404790 42288 404818
rect 41892 404652 41920 404790
rect 41722 404624 41920 404652
rect 41788 404524 41840 404530
rect 41788 404466 41840 404472
rect 41800 404002 41828 404466
rect 41722 403974 41828 404002
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41722 400947 41828 400975
rect 41800 400450 41828 400947
rect 41788 400444 41840 400450
rect 41788 400386 41840 400392
rect 41722 400302 41828 400330
rect 41800 400194 41828 400302
rect 42260 400194 42288 404790
rect 42444 404530 42472 532102
rect 42536 422294 42564 539106
rect 42628 538214 42656 571610
rect 42628 538186 42748 538214
rect 42720 528494 42748 538186
rect 42708 528488 42760 528494
rect 42708 528430 42760 528436
rect 42536 422266 42656 422294
rect 42628 410990 42656 422266
rect 42616 410984 42668 410990
rect 42616 410926 42668 410932
rect 42432 404524 42484 404530
rect 42432 404466 42484 404472
rect 42444 402974 42472 404466
rect 42444 402946 42564 402974
rect 42432 400444 42484 400450
rect 42432 400386 42484 400392
rect 41800 400166 42288 400194
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41722 370075 41828 370103
rect 41800 369578 41828 370075
rect 41788 369572 41840 369578
rect 41788 369514 41840 369520
rect 41713 369417 42193 369473
rect 41788 368688 41840 368694
rect 41788 368630 41840 368636
rect 41800 368263 41828 368630
rect 41722 368235 41828 368263
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41788 362636 41840 362642
rect 41788 362578 41840 362584
rect 41800 362094 41828 362578
rect 42260 362386 42288 400166
rect 42340 369572 42392 369578
rect 42340 369514 42392 369520
rect 42352 362642 42380 369514
rect 42340 362636 42392 362642
rect 42340 362578 42392 362584
rect 42260 362358 42380 362386
rect 41722 362066 41828 362094
rect 42352 361570 42380 362358
rect 41892 361542 42380 361570
rect 41892 361464 41920 361542
rect 41722 361436 41920 361464
rect 41722 360783 41828 360811
rect 41800 360398 41828 360783
rect 41788 360392 41840 360398
rect 41788 360334 41840 360340
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41722 357734 41828 357762
rect 41800 357270 41828 357734
rect 41788 357264 41840 357270
rect 41788 357206 41840 357212
rect 42260 357131 42288 361542
rect 42444 357270 42472 400386
rect 42536 360398 42564 402946
rect 42628 368694 42656 410926
rect 42720 400450 42748 528430
rect 674116 427854 674144 994082
rect 674208 953358 674236 994374
rect 674288 994364 674340 994370
rect 674288 994306 674340 994312
rect 674300 964170 674328 994306
rect 674380 994296 674432 994302
rect 674380 994238 674432 994244
rect 674392 967434 674420 994238
rect 675116 994228 675168 994234
rect 675116 994170 675168 994176
rect 675128 982574 675156 994170
rect 675128 982546 675340 982574
rect 674380 967428 674432 967434
rect 674380 967370 674432 967376
rect 675208 967428 675260 967434
rect 675208 967370 675260 967376
rect 675220 965326 675248 967370
rect 675208 965320 675260 965326
rect 675036 965268 675208 965274
rect 675036 965262 675260 965268
rect 675036 965246 675248 965262
rect 674288 964164 674340 964170
rect 674288 964106 674340 964112
rect 675036 963254 675064 965246
rect 675312 964253 675340 982546
rect 675407 966695 675887 966751
rect 675407 966051 675887 966107
rect 675407 965407 675887 965463
rect 675392 965320 675444 965326
rect 675392 965262 675444 965268
rect 675404 964883 675432 965262
rect 675220 964225 675418 964253
rect 675036 963226 675156 963254
rect 674932 960696 674984 960702
rect 674932 960638 674984 960644
rect 674196 953352 674248 953358
rect 674196 953294 674248 953300
rect 674840 874540 674892 874546
rect 674840 874482 674892 874488
rect 674852 785330 674880 874482
rect 674944 871706 674972 960638
rect 675128 960106 675156 963226
rect 675220 960226 675248 964225
rect 675300 964164 675352 964170
rect 675300 964106 675352 964112
rect 675312 961194 675340 964106
rect 675407 963567 675887 963623
rect 675407 963015 675887 963071
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 675312 961180 675418 961194
rect 675312 961166 675432 961180
rect 675404 960702 675432 961166
rect 675392 960696 675444 960702
rect 675392 960638 675444 960644
rect 675208 960220 675260 960226
rect 675208 960162 675260 960168
rect 675404 960106 675432 960559
rect 675128 960078 675432 960106
rect 675128 953594 675156 960078
rect 675208 960016 675260 960022
rect 675208 959958 675260 959964
rect 675036 953566 675156 953594
rect 675036 875838 675064 953566
rect 675116 953352 675168 953358
rect 675116 953294 675168 953300
rect 675024 875832 675076 875838
rect 675024 875774 675076 875780
rect 674944 871690 675064 871706
rect 674944 871684 675076 871690
rect 674944 871678 675024 871684
rect 675024 871626 675076 871632
rect 674932 864136 674984 864142
rect 674932 864078 674984 864084
rect 674840 785324 674892 785330
rect 674840 785266 674892 785272
rect 674852 740382 674880 785266
rect 674944 775062 674972 864078
rect 675036 783290 675064 871626
rect 675128 864142 675156 953294
rect 675220 874546 675248 959958
rect 675312 959901 675418 959929
rect 675312 951810 675340 959901
rect 675407 959243 675887 959299
rect 675407 958691 675887 958747
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 675407 956207 675887 956263
rect 675407 955011 675887 955067
rect 675407 954367 675887 954423
rect 675404 953594 675432 953751
rect 675404 953566 675616 953594
rect 675588 953358 675616 953566
rect 675576 953352 675628 953358
rect 675576 953294 675628 953300
rect 675407 952527 675887 952583
rect 675404 951810 675432 951932
rect 675312 951782 675432 951810
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675392 875832 675444 875838
rect 675392 875774 675444 875780
rect 675404 875242 675432 875774
rect 675312 875214 675432 875242
rect 675208 874540 675260 874546
rect 675208 874482 675260 874488
rect 675312 871298 675340 875214
rect 675404 874546 675432 875039
rect 675392 874540 675444 874546
rect 675392 874482 675444 874488
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675404 871690 675432 872003
rect 675392 871684 675444 871690
rect 675392 871626 675444 871632
rect 675404 871298 675432 871359
rect 675220 871270 675432 871298
rect 675116 864136 675168 864142
rect 675116 864078 675168 864084
rect 675220 786622 675248 871270
rect 675404 870210 675432 870740
rect 675312 870182 675432 870210
rect 675312 862730 675340 870182
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675404 864142 675432 864551
rect 675392 864136 675444 864142
rect 675392 864078 675444 864084
rect 675407 863327 675887 863383
rect 675312 862702 675418 862730
rect 677506 818408 677562 818417
rect 675300 818372 675352 818378
rect 677506 818343 677508 818352
rect 675300 818314 675352 818320
rect 677560 818343 677562 818352
rect 677508 818314 677560 818320
rect 675208 786616 675260 786622
rect 675208 786558 675260 786564
rect 675024 783284 675076 783290
rect 675024 783226 675076 783232
rect 674932 775056 674984 775062
rect 674932 774998 674984 775004
rect 674840 740376 674892 740382
rect 674840 740318 674892 740324
rect 674840 736024 674892 736030
rect 674840 735966 674892 735972
rect 674852 729094 674880 735966
rect 674944 729978 674972 774998
rect 675036 737322 675064 783226
rect 675220 782746 675248 786558
rect 675208 782740 675260 782746
rect 675208 782682 675260 782688
rect 675220 782626 675248 782682
rect 675128 782598 675248 782626
rect 675128 741062 675156 782598
rect 675208 781040 675260 781046
rect 675208 780982 675260 780988
rect 675220 774042 675248 780982
rect 675208 774036 675260 774042
rect 675208 773978 675260 773984
rect 675116 741056 675168 741062
rect 675116 740998 675168 741004
rect 675024 737316 675076 737322
rect 675024 737258 675076 737264
rect 674932 729972 674984 729978
rect 674932 729914 674984 729920
rect 674840 729088 674892 729094
rect 674840 729030 674892 729036
rect 674944 726510 674972 729914
rect 674932 726504 674984 726510
rect 674932 726446 674984 726452
rect 674932 699032 674984 699038
rect 674932 698974 674984 698980
rect 674944 696250 674972 698974
rect 674932 696244 674984 696250
rect 674932 696186 674984 696192
rect 675036 696130 675064 737258
rect 675128 737050 675156 740998
rect 675208 740376 675260 740382
rect 675208 740318 675260 740324
rect 675116 737044 675168 737050
rect 675116 736986 675168 736992
rect 674852 696102 675064 696130
rect 674852 693258 674880 696102
rect 674932 696040 674984 696046
rect 675128 695994 675156 736986
rect 675220 726594 675248 740318
rect 675312 726714 675340 818314
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675392 786616 675444 786622
rect 675392 786558 675444 786564
rect 675404 786483 675432 786558
rect 675404 785330 675432 785839
rect 675392 785324 675444 785330
rect 675392 785266 675444 785272
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675392 783284 675444 783290
rect 675392 783226 675444 783232
rect 675404 782803 675432 783226
rect 675392 782740 675444 782746
rect 675392 782682 675444 782688
rect 675404 782159 675432 782682
rect 675404 781046 675432 781524
rect 675392 781040 675444 781046
rect 675392 780982 675444 780988
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675404 775062 675432 775351
rect 675392 775056 675444 775062
rect 675392 774998 675444 775004
rect 675407 774127 675887 774183
rect 675392 774036 675444 774042
rect 675392 773978 675444 773984
rect 675404 773500 675432 773978
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 675404 741074 675432 741483
rect 675404 741062 675616 741074
rect 675404 741056 675628 741062
rect 675404 741046 675576 741056
rect 675576 740998 675628 741004
rect 675404 740382 675432 740860
rect 675392 740376 675444 740382
rect 675392 740318 675444 740324
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675404 737322 675432 737803
rect 675392 737316 675444 737322
rect 675392 737258 675444 737264
rect 675404 737050 675432 737159
rect 675392 737044 675444 737050
rect 675392 736986 675444 736992
rect 675404 736030 675432 736508
rect 675392 736024 675444 736030
rect 675392 735966 675444 735972
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675404 729978 675432 730351
rect 675392 729972 675444 729978
rect 675392 729914 675444 729920
rect 675407 729127 675887 729183
rect 675392 729088 675444 729094
rect 675392 729030 675444 729036
rect 675404 728484 675432 729030
rect 675300 726708 675352 726714
rect 675300 726650 675352 726656
rect 675220 726566 675432 726594
rect 675208 726504 675260 726510
rect 675208 726446 675260 726452
rect 675300 726504 675352 726510
rect 675300 726446 675352 726452
rect 674932 695982 674984 695988
rect 674944 695366 674972 695982
rect 675036 695978 675156 695994
rect 675024 695972 675156 695978
rect 675076 695966 675156 695972
rect 675024 695914 675076 695920
rect 674932 695360 674984 695366
rect 674932 695302 674984 695308
rect 674840 693252 674892 693258
rect 674840 693194 674892 693200
rect 674852 648038 674880 693194
rect 674944 650146 674972 695302
rect 675036 692102 675064 695914
rect 675220 693410 675248 726446
rect 675128 693382 675248 693410
rect 675024 692096 675076 692102
rect 675024 692038 675076 692044
rect 675036 683114 675064 692038
rect 675128 685234 675156 693382
rect 675208 691688 675260 691694
rect 675208 691630 675260 691636
rect 675116 685228 675168 685234
rect 675116 685170 675168 685176
rect 675128 683890 675156 685170
rect 675220 684078 675248 691630
rect 675312 691626 675340 726446
rect 675404 699038 675432 726566
rect 675392 699032 675444 699038
rect 675392 698974 675444 698980
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675404 695978 675432 696483
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675404 695366 675432 695844
rect 675392 695360 675444 695366
rect 675392 695302 675444 695308
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675392 693252 675444 693258
rect 675392 693194 675444 693200
rect 675404 692803 675432 693194
rect 675404 692102 675432 692172
rect 675392 692096 675444 692102
rect 675392 692038 675444 692044
rect 675392 691688 675444 691694
rect 675392 691630 675444 691636
rect 675300 691620 675352 691626
rect 675300 691562 675352 691568
rect 675404 691492 675432 691630
rect 675300 691416 675352 691422
rect 675300 691358 675352 691364
rect 675208 684072 675260 684078
rect 675208 684014 675260 684020
rect 675128 683862 675248 683890
rect 675036 683086 675156 683114
rect 675128 674218 675156 683086
rect 675116 674212 675168 674218
rect 675116 674154 675168 674160
rect 675116 674008 675168 674014
rect 675116 673950 675168 673956
rect 675024 671424 675076 671430
rect 675024 671366 675076 671372
rect 674932 650140 674984 650146
rect 674932 650082 674984 650088
rect 674840 648032 674892 648038
rect 674840 647974 674892 647980
rect 674852 602410 674880 647974
rect 674944 605538 674972 650082
rect 675036 639810 675064 671366
rect 675128 651438 675156 673950
rect 675220 671430 675248 683862
rect 675208 671424 675260 671430
rect 675208 671366 675260 671372
rect 675116 651432 675168 651438
rect 675116 651374 675168 651380
rect 675128 647494 675156 651374
rect 675116 647488 675168 647494
rect 675116 647430 675168 647436
rect 675024 639804 675076 639810
rect 675024 639746 675076 639752
rect 674932 605532 674984 605538
rect 674932 605474 674984 605480
rect 674840 602404 674892 602410
rect 674840 602346 674892 602352
rect 674944 602290 674972 605474
rect 674760 602262 674972 602290
rect 674760 602018 674788 602262
rect 674932 602132 674984 602138
rect 674932 602074 674984 602080
rect 674760 601990 674880 602018
rect 674852 560998 674880 601990
rect 674840 560992 674892 560998
rect 674840 560934 674892 560940
rect 674104 427848 674156 427854
rect 674104 427790 674156 427796
rect 42708 400444 42760 400450
rect 42708 400386 42760 400392
rect 674852 383790 674880 560934
rect 674944 557870 674972 602074
rect 675036 594726 675064 639746
rect 675128 605810 675156 647430
rect 675208 645788 675260 645794
rect 675208 645730 675260 645736
rect 675220 638858 675248 645730
rect 675208 638852 675260 638858
rect 675208 638794 675260 638800
rect 675116 605804 675168 605810
rect 675116 605746 675168 605752
rect 675128 601866 675156 605746
rect 675116 601860 675168 601866
rect 675116 601802 675168 601808
rect 675024 594720 675076 594726
rect 675024 594662 675076 594668
rect 674932 557864 674984 557870
rect 674932 557806 674984 557812
rect 675036 550526 675064 594662
rect 675128 561542 675156 601802
rect 675208 600840 675260 600846
rect 675208 600782 675260 600788
rect 675220 593842 675248 600782
rect 675208 593836 675260 593842
rect 675208 593778 675260 593784
rect 675116 561536 675168 561542
rect 675116 561478 675168 561484
rect 675128 557190 675156 561478
rect 675312 557534 675340 691358
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675404 685234 675432 685372
rect 675392 685228 675444 685234
rect 675392 685170 675444 685176
rect 675407 684127 675887 684183
rect 675392 684072 675444 684078
rect 675392 684014 675444 684020
rect 675404 683511 675432 684014
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675392 651432 675444 651438
rect 675392 651374 675444 651380
rect 675404 651283 675432 651374
rect 675404 650146 675432 650639
rect 675392 650140 675444 650146
rect 675392 650082 675444 650088
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675392 648032 675444 648038
rect 675392 647974 675444 647980
rect 675404 647603 675432 647974
rect 675392 647488 675444 647494
rect 675392 647430 675444 647436
rect 675404 646959 675432 647430
rect 675404 645794 675432 646340
rect 675392 645788 675444 645794
rect 675392 645730 675444 645736
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675404 639810 675432 640151
rect 675392 639804 675444 639810
rect 675392 639746 675444 639752
rect 675407 638927 675887 638983
rect 675392 638852 675444 638858
rect 675392 638794 675444 638800
rect 675404 638316 675432 638794
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675404 605834 675432 606283
rect 675404 605810 675616 605834
rect 675404 605806 675628 605810
rect 675576 605804 675628 605806
rect 675576 605746 675628 605752
rect 675404 605538 675432 605639
rect 675392 605532 675444 605538
rect 675392 605474 675444 605480
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675404 602138 675432 602603
rect 675392 602132 675444 602138
rect 675392 602074 675444 602080
rect 675404 601866 675432 601959
rect 675392 601860 675444 601866
rect 675392 601802 675444 601808
rect 675404 600846 675432 601324
rect 675392 600840 675444 600846
rect 675392 600782 675444 600788
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675404 594726 675432 595151
rect 675392 594720 675444 594726
rect 675392 594662 675444 594668
rect 675407 593927 675887 593983
rect 675392 593836 675444 593842
rect 675392 593778 675444 593784
rect 675404 593300 675432 593778
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675392 561536 675444 561542
rect 675392 561478 675444 561484
rect 675404 561068 675432 561478
rect 675392 560992 675444 560998
rect 675392 560934 675444 560940
rect 675404 560439 675432 560934
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675392 557864 675444 557870
rect 675392 557806 675444 557812
rect 675220 557506 675340 557534
rect 675116 557184 675168 557190
rect 675116 557126 675168 557132
rect 675220 555778 675248 557506
rect 675404 557396 675432 557806
rect 675392 557184 675444 557190
rect 675392 557126 675444 557132
rect 675404 556759 675432 557126
rect 675128 555750 675248 555778
rect 675024 550520 675076 550526
rect 675024 550462 675076 550468
rect 675128 547874 675156 555750
rect 675404 555626 675432 556115
rect 675208 555620 675260 555626
rect 675208 555562 675260 555568
rect 675392 555620 675444 555626
rect 675392 555562 675444 555568
rect 675220 548125 675248 555562
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675392 550520 675444 550526
rect 675392 550462 675444 550468
rect 675404 549951 675432 550462
rect 675407 548727 675887 548783
rect 675220 548097 675418 548125
rect 675128 547846 675340 547874
rect 675312 503946 675340 547846
rect 675300 503940 675352 503946
rect 675300 503882 675352 503888
rect 677428 503940 677480 503946
rect 677428 503882 677480 503888
rect 677440 503849 677468 503882
rect 677426 503840 677482 503849
rect 677426 503775 677482 503784
rect 677448 427848 677500 427854
rect 677448 427790 677500 427796
rect 677460 425629 677488 427790
rect 677446 425620 677502 425629
rect 677446 425555 677502 425564
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675220 383982 675432 384010
rect 674840 383784 674892 383790
rect 674840 383726 674892 383732
rect 674852 379514 674880 383726
rect 675024 379840 675076 379846
rect 675024 379782 675076 379788
rect 674852 379486 674972 379514
rect 674840 378412 674892 378418
rect 674840 378354 674892 378360
rect 674852 371482 674880 378354
rect 674840 371476 674892 371482
rect 674840 371418 674892 371424
rect 42616 368688 42668 368694
rect 42616 368630 42668 368636
rect 42524 360392 42576 360398
rect 42524 360334 42576 360340
rect 42432 357264 42484 357270
rect 42432 357206 42484 357212
rect 41722 357103 42380 357131
rect 42248 357060 42300 357066
rect 42248 357002 42300 357008
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 41722 326862 41828 326890
rect 41800 326398 41828 326862
rect 41788 326392 41840 326398
rect 41788 326334 41840 326340
rect 41713 326217 42193 326273
rect 41788 325168 41840 325174
rect 41788 325110 41840 325116
rect 41800 325063 41828 325110
rect 41722 325035 41828 325063
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41788 319456 41840 319462
rect 41788 319398 41840 319404
rect 41800 318899 41828 319398
rect 41722 318871 41828 318899
rect 41788 318776 41840 318782
rect 41788 318718 41840 318724
rect 41800 318255 41828 318718
rect 41722 318227 41828 318255
rect 41788 318164 41840 318170
rect 41788 318106 41840 318112
rect 41800 317611 41828 318106
rect 41722 317583 41828 317611
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41722 314547 41828 314575
rect 41800 314106 41828 314547
rect 42260 314106 42288 357002
rect 42352 318782 42380 357103
rect 42432 326392 42484 326398
rect 42432 326334 42484 326340
rect 42444 319462 42472 326334
rect 42628 325694 42656 368630
rect 42708 360392 42760 360398
rect 42708 360334 42760 360340
rect 42536 325666 42656 325694
rect 42536 325174 42564 325666
rect 42524 325168 42576 325174
rect 42524 325110 42576 325116
rect 42432 319456 42484 319462
rect 42432 319398 42484 319404
rect 42340 318776 42392 318782
rect 42340 318718 42392 318724
rect 41800 314078 42288 314106
rect 41722 313903 41828 313931
rect 41800 313546 41828 313903
rect 41788 313540 41840 313546
rect 41788 313482 41840 313488
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 41722 283675 41828 283703
rect 41800 283218 41828 283675
rect 41788 283212 41840 283218
rect 41788 283154 41840 283160
rect 41713 283017 42193 283073
rect 41788 282124 41840 282130
rect 41788 282066 41840 282072
rect 41800 281874 41828 282066
rect 41722 281846 41828 281874
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41788 276208 41840 276214
rect 41788 276150 41840 276156
rect 41800 275699 41828 276150
rect 41722 275671 41828 275699
rect 41722 275026 41828 275054
rect 41800 274582 41828 275026
rect 41788 274576 41840 274582
rect 41788 274518 41840 274524
rect 41722 274386 41828 274414
rect 41800 273970 41828 274386
rect 41788 273964 41840 273970
rect 41788 273906 41840 273912
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 42260 271538 42288 314078
rect 42352 313546 42380 318718
rect 42340 313540 42392 313546
rect 42340 313482 42392 313488
rect 42352 274582 42380 313482
rect 42432 283212 42484 283218
rect 42432 283154 42484 283160
rect 42444 276214 42472 283154
rect 42536 282130 42564 325110
rect 42720 318170 42748 360334
rect 674944 337550 674972 379486
rect 674932 337544 674984 337550
rect 674932 337486 674984 337492
rect 674840 328092 674892 328098
rect 674840 328034 674892 328040
rect 42708 318164 42760 318170
rect 42708 318106 42760 318112
rect 42720 316034 42748 318106
rect 42628 316006 42748 316034
rect 42524 282124 42576 282130
rect 42524 282066 42576 282072
rect 42432 276208 42484 276214
rect 42432 276150 42484 276156
rect 42340 274576 42392 274582
rect 42340 274518 42392 274524
rect 41800 271510 42288 271538
rect 41800 271382 41828 271510
rect 41722 271354 41828 271382
rect 41722 270694 41828 270722
rect 41800 270638 41828 270694
rect 41788 270632 41840 270638
rect 41788 270574 41840 270580
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 41722 240502 41828 240530
rect 41800 239970 41828 240502
rect 41788 239964 41840 239970
rect 41788 239906 41840 239912
rect 41713 239817 42193 239873
rect 41722 238635 41828 238663
rect 41800 238542 41828 238635
rect 41788 238536 41840 238542
rect 41788 238478 41840 238484
rect 41713 237977 42193 238033
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 41788 233028 41840 233034
rect 41788 232970 41840 232976
rect 41800 232506 41828 232970
rect 41722 232478 41828 232506
rect 41788 232416 41840 232422
rect 41788 232358 41840 232364
rect 41800 231855 41828 232358
rect 41722 231827 41828 231855
rect 41788 231736 41840 231742
rect 41788 231678 41840 231684
rect 41800 231211 41828 231678
rect 41722 231183 41828 231211
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41722 228146 41828 228174
rect 41800 227610 41828 228146
rect 42260 227610 42288 271510
rect 42352 270638 42380 274518
rect 42340 270632 42392 270638
rect 42340 270574 42392 270580
rect 42352 232422 42380 270574
rect 42432 239964 42484 239970
rect 42432 239906 42484 239912
rect 42444 233034 42472 239906
rect 42536 238542 42564 282066
rect 42628 273970 42656 316006
rect 674852 282334 674880 328034
rect 674944 293282 674972 337486
rect 675036 335442 675064 379782
rect 675220 379573 675248 383982
rect 675404 383860 675432 383982
rect 675392 383784 675444 383790
rect 675392 383726 675444 383732
rect 675404 383239 675432 383726
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675404 379846 675432 380188
rect 675392 379840 675444 379846
rect 675392 379782 675444 379788
rect 675220 379545 675418 379573
rect 675220 373994 675248 379545
rect 675404 378418 675432 378915
rect 675392 378412 675444 378418
rect 675392 378354 675444 378360
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675128 373966 675248 373994
rect 675128 338842 675156 373966
rect 675407 373367 675887 373423
rect 675220 372737 675418 372765
rect 675116 338836 675168 338842
rect 675116 338778 675168 338784
rect 675220 336002 675248 372737
rect 675407 371527 675887 371583
rect 675392 371476 675444 371482
rect 675392 371418 675444 371424
rect 675404 370911 675432 371418
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675392 338836 675444 338842
rect 675392 338778 675444 338784
rect 675404 338178 675432 338778
rect 675128 335974 675248 336002
rect 675312 338150 675432 338178
rect 675024 335436 675076 335442
rect 675024 335378 675076 335384
rect 675024 334280 675076 334286
rect 675024 334222 675076 334228
rect 675036 294166 675064 334222
rect 675128 328098 675156 335974
rect 675208 335436 675260 335442
rect 675208 335378 675260 335384
rect 675116 328092 675168 328098
rect 675116 328034 675168 328040
rect 675220 316034 675248 335378
rect 675312 334370 675340 338150
rect 675404 337550 675432 338028
rect 675392 337544 675444 337550
rect 675392 337486 675444 337492
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675392 335436 675444 335442
rect 675392 335378 675444 335384
rect 675404 335003 675432 335378
rect 675312 334356 675418 334370
rect 675312 334342 675432 334356
rect 675404 334286 675432 334342
rect 675392 334280 675444 334286
rect 675392 334222 675444 334228
rect 675312 333701 675418 333729
rect 675312 325725 675340 333701
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675392 328092 675444 328098
rect 675392 328034 675444 328040
rect 675404 327556 675432 328034
rect 675407 326327 675887 326383
rect 675312 325697 675418 325725
rect 675128 316006 675248 316034
rect 675128 306374 675156 316006
rect 675128 306346 675248 306374
rect 675220 302234 675248 306346
rect 675220 302206 675340 302234
rect 675024 294160 675076 294166
rect 675024 294102 675076 294108
rect 675312 293978 675340 302206
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675392 294160 675444 294166
rect 675392 294102 675444 294108
rect 675128 293950 675340 293978
rect 674932 293276 674984 293282
rect 674932 293218 674984 293224
rect 674944 289814 674972 293218
rect 674944 289786 675064 289814
rect 674932 289536 674984 289542
rect 674932 289478 674984 289484
rect 674840 282328 674892 282334
rect 674840 282270 674892 282276
rect 42616 273964 42668 273970
rect 42616 273906 42668 273912
rect 42524 238536 42576 238542
rect 42524 238478 42576 238484
rect 42432 233028 42484 233034
rect 42432 232970 42484 232976
rect 42340 232416 42392 232422
rect 42340 232358 42392 232364
rect 41800 227582 42288 227610
rect 41722 227503 41828 227531
rect 41800 227118 41828 227503
rect 41788 227112 41840 227118
rect 41788 227054 41840 227060
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41722 197274 41828 197302
rect 41800 196790 41828 197274
rect 41788 196784 41840 196790
rect 41788 196726 41840 196732
rect 41713 196617 42193 196673
rect 41722 195435 41828 195463
rect 41800 195362 41828 195435
rect 41788 195356 41840 195362
rect 41788 195298 41840 195304
rect 41713 194777 42193 194833
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41788 189848 41840 189854
rect 41788 189790 41840 189796
rect 41800 189299 41828 189790
rect 41722 189271 41828 189299
rect 41722 188627 41828 188655
rect 41800 188154 41828 188627
rect 41788 188148 41840 188154
rect 41788 188090 41840 188096
rect 41722 187986 41828 188014
rect 41800 187610 41828 187986
rect 41788 187604 41840 187610
rect 41788 187546 41840 187552
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 42260 184975 42288 227582
rect 42352 227118 42380 232358
rect 42340 227112 42392 227118
rect 42340 227054 42392 227060
rect 42352 188154 42380 227054
rect 42536 200114 42564 238478
rect 42628 231742 42656 273906
rect 674852 237726 674880 282270
rect 674944 244526 674972 289478
rect 675036 288658 675064 289786
rect 675128 289542 675156 293950
rect 675404 293706 675432 294102
rect 675312 293692 675432 293706
rect 675312 293678 675418 293692
rect 675116 289536 675168 289542
rect 675116 289478 675168 289484
rect 675312 289354 675340 293678
rect 675392 293276 675444 293282
rect 675392 293218 675444 293224
rect 675404 293012 675432 293218
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675404 289542 675432 290020
rect 675392 289536 675444 289542
rect 675392 289478 675444 289484
rect 675312 289340 675418 289354
rect 675312 289326 675432 289340
rect 675404 288810 675432 289326
rect 675128 288782 675432 288810
rect 675024 288652 675076 288658
rect 675024 288594 675076 288600
rect 675128 248810 675156 288782
rect 675220 288701 675418 288729
rect 675220 281246 675248 288701
rect 675300 288652 675352 288658
rect 675300 288594 675352 288600
rect 675208 281240 675260 281246
rect 675208 281182 675260 281188
rect 675116 248804 675168 248810
rect 675116 248746 675168 248752
rect 675128 248414 675156 248746
rect 675312 248554 675340 288594
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675404 282334 675432 282540
rect 675392 282328 675444 282334
rect 675392 282270 675444 282276
rect 675407 281327 675887 281383
rect 675392 281240 675444 281246
rect 675392 281182 675444 281188
rect 675404 280711 675432 281182
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675392 248804 675444 248810
rect 675392 248746 675444 248752
rect 675404 248676 675432 248746
rect 675312 248526 675432 248554
rect 675128 248386 675340 248414
rect 675024 247512 675076 247518
rect 675024 247454 675076 247460
rect 674932 244520 674984 244526
rect 674932 244462 674984 244468
rect 674840 237720 674892 237726
rect 674840 237662 674892 237668
rect 42616 231736 42668 231742
rect 42616 231678 42668 231684
rect 42444 200086 42564 200114
rect 42444 195362 42472 200086
rect 42432 195356 42484 195362
rect 42432 195298 42484 195304
rect 42340 188148 42392 188154
rect 42340 188090 42392 188096
rect 41722 184947 42288 184975
rect 41722 184303 41828 184331
rect 41800 184210 41828 184303
rect 41788 184204 41840 184210
rect 41788 184146 41840 184152
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 42062 113248 42118 113257
rect 42062 113183 42118 113192
rect 42076 42418 42104 113183
rect 42154 78296 42210 78305
rect 42154 78231 42210 78240
rect 42168 42486 42196 78231
rect 42156 42480 42208 42486
rect 42156 42422 42208 42428
rect 42064 42412 42116 42418
rect 42064 42354 42116 42360
rect 42260 42158 42288 184947
rect 42352 184210 42380 188090
rect 42340 184204 42392 184210
rect 42340 184146 42392 184152
rect 42248 42152 42300 42158
rect 42248 42094 42300 42100
rect 42352 42090 42380 184146
rect 42444 78305 42472 195298
rect 42628 190454 42656 231678
rect 674944 200258 674972 244462
rect 675036 202366 675064 247454
rect 675312 244373 675340 248386
rect 675404 247518 675432 248526
rect 675392 247512 675444 247518
rect 675392 247454 675444 247460
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675404 244526 675432 245004
rect 675392 244520 675444 244526
rect 675392 244462 675444 244468
rect 675312 244345 675418 244373
rect 675312 243794 675340 244345
rect 675128 243766 675340 243794
rect 675128 203522 675156 243766
rect 675220 243701 675418 243729
rect 675220 236298 675248 243701
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675392 237720 675444 237726
rect 675392 237662 675444 237668
rect 675404 237130 675432 237662
rect 675312 237102 675432 237130
rect 675208 236292 675260 236298
rect 675208 236234 675260 236240
rect 675312 205634 675340 237102
rect 675407 236327 675887 236383
rect 675392 236292 675444 236298
rect 675392 236234 675444 236240
rect 675404 235711 675432 236234
rect 675220 205606 675340 205634
rect 675116 203516 675168 203522
rect 675116 203458 675168 203464
rect 675024 202360 675076 202366
rect 675024 202302 675076 202308
rect 674932 200252 674984 200258
rect 674932 200194 674984 200200
rect 42708 196784 42760 196790
rect 42708 196726 42760 196732
rect 42536 190426 42656 190454
rect 42536 187610 42564 190426
rect 42720 189854 42748 196726
rect 42708 189848 42760 189854
rect 42708 189790 42760 189796
rect 42524 187604 42576 187610
rect 42524 187546 42576 187552
rect 42536 113257 42564 187546
rect 674840 157344 674892 157350
rect 674840 157286 674892 157292
rect 42522 113248 42578 113257
rect 42522 113183 42578 113192
rect 674852 112538 674880 157286
rect 674944 155242 674972 200194
rect 675036 157350 675064 202302
rect 675220 199306 675248 205606
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675312 203522 675340 203580
rect 675300 203516 675352 203522
rect 675352 203469 675418 203497
rect 675300 203458 675352 203464
rect 675208 199300 675260 199306
rect 675208 199242 675260 199248
rect 675312 199186 675340 203458
rect 675404 202366 675432 202844
rect 675392 202360 675444 202366
rect 675392 202302 675444 202308
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675392 200252 675444 200258
rect 675392 200194 675444 200200
rect 675404 199803 675432 200194
rect 675128 199158 675418 199186
rect 675128 158658 675156 199158
rect 675208 199096 675260 199102
rect 675208 199038 675260 199044
rect 675220 191962 675248 199038
rect 675312 198614 675432 198642
rect 675208 191956 675260 191962
rect 675208 191898 675260 191904
rect 675220 171134 675248 191898
rect 675312 190525 675340 198614
rect 675404 198492 675432 198614
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675404 191962 675432 192372
rect 675392 191956 675444 191962
rect 675392 191898 675444 191904
rect 675407 191127 675887 191183
rect 675312 190497 675418 190525
rect 675220 171106 675340 171134
rect 675312 158778 675340 171106
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675300 158772 675352 158778
rect 675300 158714 675352 158720
rect 675128 158630 675340 158658
rect 675116 158568 675168 158574
rect 675116 158510 675168 158516
rect 675024 157344 675076 157350
rect 675024 157286 675076 157292
rect 675128 156618 675156 158510
rect 675036 156590 675156 156618
rect 675312 158386 675340 158630
rect 675404 158386 675432 158508
rect 675312 158358 675432 158386
rect 674932 155236 674984 155242
rect 674932 155178 674984 155184
rect 674840 112532 674892 112538
rect 674840 112474 674892 112480
rect 42430 78296 42486 78305
rect 42430 78231 42486 78240
rect 527456 43208 527508 43214
rect 527456 43150 527508 43156
rect 523776 43140 523828 43146
rect 523776 43082 523828 43088
rect 516140 43072 516192 43078
rect 516140 43014 516192 43020
rect 459652 43004 459704 43010
rect 459652 42946 459704 42952
rect 467656 43004 467708 43010
rect 467656 42946 467708 42952
rect 415308 42936 415360 42942
rect 415308 42878 415360 42884
rect 411076 42868 411128 42874
rect 411076 42810 411128 42816
rect 295248 42800 295300 42806
rect 195980 42772 196032 42778
rect 295248 42742 295300 42748
rect 303252 42800 303304 42806
rect 303252 42742 303304 42748
rect 350080 42800 350132 42806
rect 350080 42742 350132 42748
rect 358084 42800 358136 42806
rect 358084 42742 358136 42748
rect 360568 42800 360620 42806
rect 360568 42742 360620 42748
rect 406752 42800 406804 42806
rect 406752 42742 406804 42748
rect 195980 42714 196032 42720
rect 188528 42596 188580 42602
rect 188528 42538 188580 42544
rect 192852 42596 192904 42602
rect 192852 42538 192904 42544
rect 147680 42480 147732 42486
rect 188540 42466 188568 42538
rect 147680 42422 147732 42428
rect 188528 42460 188580 42466
rect 88800 42304 88852 42310
rect 88800 42246 88852 42252
rect 42340 42084 42392 42090
rect 42340 42026 42392 42032
rect 88812 39953 88840 42246
rect 140964 42152 141016 42158
rect 147692 42106 147720 42422
rect 188528 42402 188580 42408
rect 186688 42392 186740 42398
rect 186688 42334 186740 42340
rect 140964 42094 141016 42100
rect 147680 42100 147732 42106
rect 140976 40202 141004 42094
rect 145104 42084 145156 42090
rect 147680 42042 147732 42048
rect 145104 42026 145156 42032
rect 145116 41478 145144 42026
rect 143080 41472 143132 41478
rect 143080 41414 143132 41420
rect 145104 41472 145156 41478
rect 145104 41414 145156 41420
rect 143092 40361 143120 41414
rect 144644 41404 144696 41410
rect 144644 41346 144696 41352
rect 143078 40352 143134 40361
rect 143078 40287 143134 40296
rect 140976 40174 141036 40202
rect 141008 40118 141036 40174
rect 143092 40118 143120 40287
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143080 40112 143132 40118
rect 143080 40054 143132 40060
rect 141008 39984 141036 40054
rect 143092 39982 143120 40054
rect 144656 39982 144684 41346
rect 145116 40202 145144 41414
rect 145103 40174 145144 40202
rect 145103 40000 145131 40174
rect 145091 39986 145143 40000
rect 147692 39953 147720 42042
rect 186136 41880 186188 41886
rect 186136 41822 186188 41828
rect 186148 41478 186176 41822
rect 186700 41820 186728 42334
rect 187327 41713 187383 42193
rect 188540 41820 188568 42402
rect 189198 41818 189304 41834
rect 191038 41818 191144 41834
rect 192234 41818 192340 41834
rect 192864 41820 192892 42538
rect 195992 42466 196020 42714
rect 199016 42664 199068 42670
rect 199016 42606 199068 42612
rect 200856 42664 200908 42670
rect 200856 42606 200908 42612
rect 241336 42664 241388 42670
rect 241336 42606 241388 42612
rect 195980 42460 196032 42466
rect 195980 42402 196032 42408
rect 194692 42392 194744 42398
rect 194692 42334 194744 42340
rect 193522 41818 193628 41834
rect 189198 41812 189316 41818
rect 189198 41806 189264 41812
rect 191038 41812 191156 41818
rect 191038 41806 191104 41812
rect 189264 41754 189316 41760
rect 192234 41812 192352 41818
rect 192234 41806 192300 41812
rect 191104 41754 191156 41760
rect 193522 41812 193640 41818
rect 193522 41806 193588 41812
rect 192300 41754 192352 41760
rect 193588 41754 193640 41760
rect 194043 41713 194099 42193
rect 194704 41820 194732 42334
rect 195244 41880 195296 41886
rect 195296 41828 195362 41834
rect 195244 41822 195362 41828
rect 195256 41806 195362 41822
rect 195992 41820 196020 42402
rect 198464 41948 198516 41954
rect 198464 41890 198516 41896
rect 198476 41834 198504 41890
rect 196452 41818 198504 41834
rect 199028 41820 199056 42606
rect 199660 42528 199712 42534
rect 199660 42470 199712 42476
rect 199568 41880 199620 41886
rect 199672 41834 199700 42470
rect 200120 41948 200172 41954
rect 200120 41890 200172 41896
rect 199620 41828 199700 41834
rect 199568 41822 199700 41828
rect 199580 41820 199700 41822
rect 200132 41834 200160 41890
rect 200868 41834 200896 42606
rect 201500 42596 201552 42602
rect 201500 42538 201552 42544
rect 200132 41820 200896 41834
rect 201512 41820 201540 42538
rect 196440 41812 198504 41818
rect 196492 41806 198504 41812
rect 199580 41806 199686 41820
rect 200132 41806 200882 41820
rect 196440 41754 196492 41760
rect 186136 41472 186188 41478
rect 186136 41414 186188 41420
rect 88798 39944 88854 39953
rect 88798 39879 88854 39888
rect 147678 39944 147734 39953
rect 147678 39879 147734 39888
rect 241348 39817 241376 42606
rect 295260 41834 295288 42742
rect 297732 42664 297784 42670
rect 297732 42606 297784 42612
rect 300768 42664 300820 42670
rect 300768 42606 300820 42612
rect 297088 42596 297140 42602
rect 297088 42538 297140 42544
rect 297100 41834 297128 42538
rect 297744 41834 297772 42606
rect 299572 42596 299624 42602
rect 299572 42538 299624 42544
rect 299584 41834 299612 42538
rect 300780 41834 300808 42606
rect 295260 41806 295311 41834
rect 297100 41806 297151 41834
rect 297744 41806 297795 41834
rect 299584 41806 299635 41834
rect 300780 41806 302119 41834
rect 302643 41713 302699 42193
rect 303264 41834 303292 42742
rect 307576 42732 307628 42738
rect 307576 42674 307628 42680
rect 305092 42664 305144 42670
rect 305092 42606 305144 42612
rect 303896 42528 303948 42534
rect 303896 42470 303948 42476
rect 303908 41834 303936 42470
rect 304540 42460 304592 42466
rect 304540 42402 304592 42408
rect 304552 41834 304580 42402
rect 305104 41834 305132 42606
rect 305736 42596 305788 42602
rect 305736 42538 305788 42544
rect 305276 41948 305328 41954
rect 305276 41890 305328 41896
rect 305288 41834 305316 41890
rect 303264 41806 303315 41834
rect 303908 41806 303959 41834
rect 304552 41806 304603 41834
rect 305104 41806 305316 41834
rect 305748 41834 305776 42538
rect 306300 41954 306420 41967
rect 306288 41948 306420 41954
rect 306340 41939 306420 41948
rect 306288 41890 306340 41896
rect 306392 41834 306420 41939
rect 305748 41806 305799 41834
rect 306392 41806 306443 41834
rect 306967 41713 307023 42193
rect 307588 41834 307616 42674
rect 309416 42664 309468 42670
rect 309416 42606 309468 42612
rect 308220 42528 308272 42534
rect 308220 42470 308272 42476
rect 308232 41834 308260 42470
rect 308680 41948 308732 41954
rect 308680 41890 308732 41896
rect 308692 41834 308720 41890
rect 309428 41834 309456 42606
rect 307588 41806 307639 41834
rect 308232 41806 308283 41834
rect 308692 41806 309479 41834
rect 310095 41713 310151 42193
rect 350092 41820 350120 42742
rect 352564 42664 352616 42670
rect 352564 42606 352616 42612
rect 355600 42664 355652 42670
rect 355600 42606 355652 42612
rect 351920 42596 351972 42602
rect 351920 42538 351972 42544
rect 351932 41820 351960 42538
rect 352576 41820 352604 42606
rect 354404 42596 354456 42602
rect 354404 42538 354456 42544
rect 354416 41820 354444 42538
rect 355612 41834 355640 42606
rect 355612 41820 356914 41834
rect 355626 41806 356914 41820
rect 357443 41713 357499 42193
rect 358096 41820 358124 42742
rect 359924 42664 359976 42670
rect 359924 42606 359976 42612
rect 358728 42528 358780 42534
rect 358728 42470 358780 42476
rect 358740 41820 358768 42470
rect 359372 42460 359424 42466
rect 359372 42402 359424 42408
rect 359384 41820 359412 42402
rect 359936 41834 359964 42606
rect 360580 42602 360608 42742
rect 362408 42732 362460 42738
rect 362408 42674 362460 42680
rect 360568 42596 360620 42602
rect 360568 42538 360620 42544
rect 359936 41820 360056 41834
rect 360580 41820 360608 42538
rect 359950 41818 360056 41820
rect 361132 41818 361238 41834
rect 359950 41812 360068 41818
rect 359950 41806 360016 41812
rect 360016 41754 360068 41760
rect 361120 41812 361238 41818
rect 361172 41806 361238 41812
rect 361120 41754 361172 41760
rect 361767 41713 361823 42193
rect 362420 41820 362448 42674
rect 364248 42664 364300 42670
rect 364248 42606 364300 42612
rect 363052 42528 363104 42534
rect 363052 42470 363104 42476
rect 363064 41820 363092 42470
rect 364260 41834 364288 42606
rect 404912 42596 404964 42602
rect 404912 42538 404964 42544
rect 363524 41820 364288 41834
rect 363524 41818 364274 41820
rect 363512 41812 364274 41818
rect 363564 41806 364274 41812
rect 363512 41754 363564 41760
rect 364895 41713 364951 42193
rect 404924 41820 404952 42538
rect 405527 41713 405583 42193
rect 406764 41820 406792 42742
rect 407396 42664 407448 42670
rect 407396 42606 407448 42612
rect 410432 42664 410484 42670
rect 410432 42606 410484 42612
rect 407408 41820 407436 42606
rect 409236 42392 409288 42398
rect 409236 42334 409288 42340
rect 409248 41820 409276 42334
rect 410444 41834 410472 42606
rect 410444 41820 410564 41834
rect 411088 41820 411116 42810
rect 412916 42596 412968 42602
rect 412916 42538 412968 42544
rect 413560 42596 413612 42602
rect 413560 42538 413612 42544
rect 412272 42392 412324 42398
rect 412272 42334 412324 42340
rect 412284 42193 412312 42334
rect 410458 41818 410564 41820
rect 411548 41818 411746 41834
rect 410458 41812 410576 41818
rect 410458 41806 410524 41812
rect 410524 41754 410576 41760
rect 411536 41812 411746 41818
rect 411588 41806 411746 41812
rect 412243 41820 412312 42193
rect 412928 41820 412956 42538
rect 413572 41820 413600 42538
rect 415320 42466 415348 42878
rect 419724 42868 419776 42874
rect 419724 42810 419776 42816
rect 417240 42732 417292 42738
rect 417240 42674 417292 42680
rect 416044 42664 416096 42670
rect 416044 42606 416096 42612
rect 414204 42460 414256 42466
rect 414204 42402 414256 42408
rect 415308 42460 415360 42466
rect 415308 42402 415360 42408
rect 414216 41820 414244 42402
rect 415400 42392 415452 42398
rect 415400 42334 415452 42340
rect 411536 41754 411588 41760
rect 412243 41713 412299 41820
rect 414782 41818 414888 41834
rect 415412 41820 415440 42334
rect 416056 41834 416084 42606
rect 415872 41820 416084 41834
rect 415872 41818 416070 41820
rect 414782 41812 414900 41818
rect 414782 41806 414848 41812
rect 414848 41754 414900 41760
rect 415860 41812 416070 41818
rect 415912 41806 416070 41812
rect 415860 41754 415912 41760
rect 416567 41713 416623 42193
rect 417252 41820 417280 42674
rect 419080 42664 419132 42670
rect 419080 42606 419132 42612
rect 417884 42596 417936 42602
rect 417884 42538 417936 42544
rect 417896 41820 417924 42538
rect 419092 41834 419120 42606
rect 419736 42193 419764 42810
rect 418462 41820 419120 41834
rect 419695 41820 419764 42193
rect 459664 41834 459692 42946
rect 461492 42868 461544 42874
rect 461492 42810 461544 42816
rect 418462 41806 419106 41820
rect 419695 41713 419751 41820
rect 459664 41806 459711 41834
rect 460327 41713 460383 42193
rect 461504 41834 461532 42810
rect 462136 42664 462188 42670
rect 462136 42606 462188 42612
rect 465172 42664 465224 42670
rect 465172 42606 465224 42612
rect 462148 41834 462176 42606
rect 464160 41880 464212 41886
rect 461504 41806 461551 41834
rect 462148 41806 462195 41834
rect 464035 41828 464160 41834
rect 464035 41822 464212 41828
rect 465184 41834 465212 42606
rect 465816 42528 465868 42534
rect 465816 42470 465868 42476
rect 465828 41834 465856 42470
rect 467043 41834 467099 42193
rect 467196 41880 467248 41886
rect 464035 41806 464200 41822
rect 465184 41818 465396 41834
rect 465184 41812 465408 41818
rect 465184 41806 465356 41812
rect 465828 41806 465875 41834
rect 466380 41818 466519 41834
rect 466368 41812 466519 41818
rect 465356 41754 465408 41760
rect 466420 41806 466519 41812
rect 467043 41828 467196 41834
rect 467043 41822 467248 41828
rect 467668 41834 467696 42946
rect 467840 42936 467892 42942
rect 467840 42878 467892 42884
rect 473268 42936 473320 42942
rect 473268 42878 473320 42884
rect 467852 42806 467880 42878
rect 467840 42800 467892 42806
rect 467840 42742 467892 42748
rect 468944 42800 468996 42806
rect 468944 42742 468996 42748
rect 468300 42596 468352 42602
rect 468300 42538 468352 42544
rect 468312 41834 468340 42538
rect 468956 41834 468984 42742
rect 473280 42738 473308 42878
rect 516152 42874 516180 43014
rect 516140 42868 516192 42874
rect 516140 42810 516192 42816
rect 471980 42732 472032 42738
rect 471980 42674 472032 42680
rect 473268 42732 473320 42738
rect 473268 42674 473320 42680
rect 514484 42732 514536 42738
rect 514484 42674 514536 42680
rect 470784 42664 470836 42670
rect 470784 42606 470836 42612
rect 469680 42016 469732 42022
rect 469680 41958 469732 41964
rect 470692 42016 470744 42022
rect 470796 41970 470824 42606
rect 470744 41964 470824 41970
rect 470692 41958 470824 41964
rect 469692 41834 469720 41958
rect 470704 41942 470824 41958
rect 467043 41806 467236 41822
rect 467668 41806 467715 41834
rect 468312 41806 468359 41834
rect 468956 41806 469003 41834
rect 469416 41818 469720 41834
rect 470048 41880 470100 41886
rect 470796 41834 470824 41942
rect 470100 41828 470199 41834
rect 470048 41822 470199 41828
rect 469404 41812 469720 41818
rect 466368 41754 466420 41760
rect 467043 41713 467099 41806
rect 469456 41806 469720 41812
rect 470060 41806 470199 41822
rect 470796 41806 470843 41834
rect 469404 41754 469456 41760
rect 471367 41713 471423 42193
rect 471992 41834 472020 42674
rect 473820 42664 473872 42670
rect 473820 42606 473872 42612
rect 472624 42596 472676 42602
rect 472624 42538 472676 42544
rect 472636 41834 472664 42538
rect 473832 41834 473860 42606
rect 474464 42528 474516 42534
rect 474464 42470 474516 42476
rect 474476 42193 474504 42470
rect 471992 41806 472039 41834
rect 472636 41806 472683 41834
rect 473235 41806 473879 41834
rect 474476 41806 474551 42193
rect 514496 41820 514524 42674
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 516152 41834 516180 42810
rect 523788 42806 523816 43082
rect 526812 42936 526864 42942
rect 526812 42878 526864 42884
rect 523776 42800 523828 42806
rect 523776 42742 523828 42748
rect 522488 42732 522540 42738
rect 522488 42674 522540 42680
rect 516968 42664 517020 42670
rect 516968 42606 517020 42612
rect 520004 42664 520056 42670
rect 520004 42606 520056 42612
rect 516152 41806 516350 41834
rect 516980 41820 517008 42606
rect 518808 42392 518860 42398
rect 518808 42334 518860 42340
rect 518820 41820 518848 42334
rect 520016 41834 520044 42606
rect 520016 41820 520136 41834
rect 520030 41818 520136 41820
rect 520030 41812 520148 41818
rect 520030 41806 520096 41812
rect 520096 41754 520148 41760
rect 520647 41713 520703 42193
rect 521212 41818 521318 41834
rect 521200 41812 521318 41818
rect 521252 41806 521318 41812
rect 521200 41754 521252 41760
rect 521843 41713 521899 42193
rect 522500 41820 522528 42674
rect 523132 42596 523184 42602
rect 523132 42538 523184 42544
rect 523144 41820 523172 42538
rect 523788 41820 523816 42742
rect 524972 42392 525024 42398
rect 524972 42334 525024 42340
rect 524984 42193 525012 42334
rect 524248 41818 524354 41834
rect 524236 41812 524354 41818
rect 524288 41806 524354 41812
rect 524236 41754 524288 41760
rect 524971 41713 525027 42193
rect 525536 41818 525642 41834
rect 525524 41812 525642 41818
rect 525576 41806 525642 41812
rect 525524 41754 525576 41760
rect 526167 41713 526223 42193
rect 526824 41820 526852 42878
rect 527468 42602 527496 43150
rect 527456 42596 527508 42602
rect 527456 42538 527508 42544
rect 527468 41820 527496 42538
rect 528480 41939 528692 41967
rect 528480 41834 528508 41939
rect 527928 41818 528508 41834
rect 528664 41820 528692 41939
rect 527916 41812 528508 41818
rect 527968 41806 528508 41812
rect 527916 41754 527968 41760
rect 529295 41713 529351 42193
rect 572720 40904 572772 40910
rect 572720 40846 572772 40852
rect 572732 40730 572760 40846
rect 674852 40730 674880 112474
rect 674944 109138 674972 155178
rect 675036 147150 675064 156590
rect 675312 154170 675340 158358
rect 675404 157350 675432 157828
rect 675392 157344 675444 157350
rect 675392 157286 675444 157292
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675392 155236 675444 155242
rect 675392 155178 675444 155184
rect 675404 154803 675432 155178
rect 675128 154142 675418 154170
rect 675024 147144 675076 147150
rect 675024 147086 675076 147092
rect 675128 142154 675156 154142
rect 675312 153501 675418 153529
rect 675208 147144 675260 147150
rect 675208 147086 675260 147092
rect 675036 142126 675156 142154
rect 675220 142154 675248 147086
rect 675312 145525 675340 153501
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675404 147150 675432 147356
rect 675392 147144 675444 147150
rect 675392 147086 675444 147092
rect 675407 146127 675887 146183
rect 675312 145497 675418 145525
rect 675220 142126 675340 142154
rect 675036 113150 675064 142126
rect 675024 113144 675076 113150
rect 675024 113086 675076 113092
rect 674932 109132 674984 109138
rect 674932 109074 674984 109080
rect 674944 41046 674972 109074
rect 675036 108866 675064 113086
rect 675024 108860 675076 108866
rect 675024 108802 675076 108808
rect 675036 41114 675064 108802
rect 675208 107840 675260 107846
rect 675208 107782 675260 107788
rect 675220 102066 675248 107782
rect 675208 102060 675260 102066
rect 675208 102002 675260 102008
rect 675312 101946 675340 142126
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675404 113150 675432 113283
rect 675392 113144 675444 113150
rect 675392 113086 675444 113092
rect 675404 112538 675432 112639
rect 675392 112532 675444 112538
rect 675392 112474 675444 112480
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675404 109138 675432 109603
rect 675392 109132 675444 109138
rect 675392 109074 675444 109080
rect 675404 108866 675432 108959
rect 675392 108860 675444 108866
rect 675392 108802 675444 108808
rect 675404 107846 675432 108324
rect 675392 107840 675444 107846
rect 675392 107782 675444 107788
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675404 101946 675432 102151
rect 675128 101918 675432 101946
rect 675024 41108 675076 41114
rect 675024 41050 675076 41056
rect 674932 41040 674984 41046
rect 674932 40982 674984 40988
rect 675128 40978 675156 101918
rect 675300 101856 675352 101862
rect 675300 101798 675352 101804
rect 675312 100314 675340 101798
rect 675407 100927 675887 100983
rect 675312 100286 675418 100314
rect 675116 40972 675168 40978
rect 675116 40914 675168 40920
rect 572720 40724 572772 40730
rect 572720 40666 572772 40672
rect 674840 40724 674892 40730
rect 674840 40666 674892 40672
rect 572732 40225 572760 40666
rect 572718 40216 572774 40225
rect 572718 40151 572774 40160
rect 241334 39808 241390 39817
rect 241334 39743 241390 39752
<< via2 >>
rect 333242 997872 333298 997928
rect 41418 881864 41474 881920
rect 41418 879960 41474 880016
rect 42246 879960 42302 880016
rect 580630 997802 580686 997858
rect 42614 881864 42670 881920
rect 677506 818372 677562 818408
rect 677506 818352 677508 818372
rect 677508 818352 677560 818372
rect 677560 818352 677562 818372
rect 677426 503784 677482 503840
rect 677446 425564 677502 425620
rect 42062 113192 42118 113248
rect 42154 78240 42210 78296
rect 42522 113192 42578 113248
rect 42430 78240 42486 78296
rect 143078 40296 143134 40352
rect 88798 39888 88854 39944
rect 147678 39888 147734 39944
rect 572718 40160 572774 40216
rect 241334 39752 241390 39808
<< metal3 >>
rect 333237 997930 333303 997933
rect 333237 997928 333530 997930
rect 333237 997872 333242 997928
rect 333298 997872 333530 997928
rect 333237 997870 333530 997872
rect 333237 997867 333303 997870
rect 333470 997628 333530 997870
rect 580625 997860 580691 997863
rect 576902 997858 580691 997860
rect 576902 997802 580630 997858
rect 580686 997802 580691 997858
rect 576902 997800 580691 997802
rect 576902 997628 576962 997800
rect 580625 997797 580691 997800
rect 40854 926876 46818 926940
rect 40854 922268 44294 926876
rect 46702 922268 46818 926876
rect 40854 922151 46818 922268
rect 670772 922374 676724 922500
rect 40854 921736 46818 921852
rect 40854 917280 41096 921736
rect 43504 917280 46818 921736
rect 670772 917822 674136 922374
rect 676496 917822 676724 922374
rect 670772 917700 676724 917822
rect 40854 917190 46818 917280
rect 670772 917268 676724 917410
rect 40854 916770 46818 916900
rect 40854 912162 44274 916770
rect 46682 912162 46818 916770
rect 670772 912862 670974 917268
rect 673314 912862 676724 917268
rect 670772 912748 676724 912862
rect 40854 912100 46818 912162
rect 670772 912322 676724 912449
rect 670772 907790 674170 912322
rect 676504 907790 676724 912322
rect 670772 907660 676724 907790
rect 41413 881922 41479 881925
rect 42609 881922 42675 881925
rect 41413 881920 42675 881922
rect 41413 881864 41418 881920
rect 41474 881864 42614 881920
rect 42670 881864 42675 881920
rect 41413 881862 42675 881864
rect 41413 881859 41479 881862
rect 42609 881859 42675 881862
rect 41413 880018 41479 880021
rect 42241 880018 42307 880021
rect 39652 880016 42307 880018
rect 39652 879960 41418 880016
rect 41474 879960 42246 880016
rect 42302 879960 42307 880016
rect 39652 879958 42307 879960
rect 41413 879955 41479 879958
rect 42241 879955 42307 879958
rect 677501 818410 677567 818413
rect 677734 818410 677794 818652
rect 677501 818408 677794 818410
rect 677501 818352 677506 818408
rect 677562 818352 677794 818408
rect 677501 818350 677794 818352
rect 677501 818347 677567 818350
rect 677421 503842 677487 503845
rect 677734 503842 677794 503948
rect 677421 503840 677794 503842
rect 677421 503784 677426 503840
rect 677482 503784 677794 503840
rect 677421 503782 677794 503784
rect 677421 503779 677487 503782
rect 670794 474564 676878 474700
rect 670794 470046 670926 474564
rect 673294 470046 676878 474564
rect 670794 469900 676878 470046
rect 670794 469480 676878 469600
rect 670794 465058 674144 469480
rect 676512 465058 676878 469480
rect 670794 464949 676878 465058
rect 670794 464548 676878 464649
rect 670794 460030 670932 464548
rect 673300 460030 676878 464548
rect 670794 459860 676878 460030
rect 41220 455654 46828 455740
rect 43508 451042 46828 455654
rect 41220 450951 46828 451042
rect 41220 450528 46828 450651
rect 41220 446104 44290 450528
rect 46690 446104 46828 450528
rect 41220 446000 46828 446104
rect 41220 445596 46828 445700
rect 43488 440984 46828 445596
rect 41220 440900 46828 440984
rect 677600 425625 677794 425748
rect 677441 425620 677794 425625
rect 677441 425564 677446 425620
rect 677502 425564 677794 425620
rect 677441 425562 677794 425564
rect 677441 425559 677507 425562
rect 42057 113250 42123 113253
rect 42517 113250 42583 113253
rect 39652 113248 42583 113250
rect 39652 113192 42062 113248
rect 42118 113192 42522 113248
rect 42578 113192 42583 113248
rect 39652 113190 42583 113192
rect 42057 113187 42123 113190
rect 42517 113187 42583 113190
rect 42149 78298 42215 78301
rect 42425 78298 42491 78301
rect 39468 78296 42491 78298
rect 39468 78240 42154 78296
rect 42210 78240 42430 78296
rect 42486 78240 42491 78296
rect 39468 78238 42491 78240
rect 42149 78235 42215 78238
rect 42425 78235 42491 78238
rect 142110 40430 144010 40490
rect 142110 40218 142170 40430
rect 143073 40354 143139 40357
rect 143073 40352 143458 40354
rect 143073 40296 143078 40352
rect 143134 40296 143458 40352
rect 143073 40294 143458 40296
rect 143073 40291 143139 40294
rect 133094 40158 142170 40218
rect 133094 39984 133154 40158
rect 143398 39984 143458 40294
rect 143950 39984 144010 40430
rect 572713 40218 572779 40221
rect 572670 40216 572779 40218
rect 572670 40160 572718 40216
rect 572774 40160 572779 40216
rect 572670 40155 572779 40160
rect 145816 40022 147690 40082
rect 145816 39996 145920 40022
rect 147630 39949 147690 40022
rect 88793 39944 88994 39949
rect 88793 39888 88798 39944
rect 88854 39888 88994 39944
rect 88793 39883 88994 39888
rect 147630 39944 147739 39949
rect 147630 39888 147678 39944
rect 147734 39888 147739 39944
rect 147630 39886 147739 39888
rect 147673 39883 147739 39886
rect 88934 39644 88994 39883
rect 241329 39810 241395 39813
rect 241286 39808 241395 39810
rect 241286 39752 241334 39808
rect 241390 39752 241395 39808
rect 241286 39747 241395 39752
rect 241286 39372 241346 39747
rect 572670 39644 572730 40155
<< via3 >>
rect 44294 922268 46702 926876
rect 41096 917280 43504 921736
rect 674136 917822 676496 922374
rect 44274 912162 46682 916770
rect 670974 912862 673314 917268
rect 674170 907790 676504 912322
rect 670926 470046 673294 474564
rect 674144 465058 676512 469480
rect 670932 460030 673300 464548
rect 41142 451042 43508 455654
rect 44290 446104 46690 450528
rect 41122 440984 43488 445596
<< metal4 >>
rect 44198 926876 46800 926958
rect 44198 922268 44294 926876
rect 46702 922268 46800 926876
rect 44198 922154 46800 922268
rect 674010 922374 676616 922486
rect 40982 921736 43584 921844
rect 40982 917280 41096 921736
rect 43504 917280 43584 921736
rect 674010 917822 674136 922374
rect 676496 917822 676616 922374
rect 674010 917716 676616 917822
rect 40982 917186 43584 917280
rect 670826 917268 673434 917414
rect 44194 916770 46796 916898
rect 44194 912162 44274 916770
rect 46682 912162 46796 916770
rect 670826 912862 670974 917268
rect 673314 912862 673434 917268
rect 670826 912756 673434 912862
rect 44194 912094 46796 912162
rect 674016 912322 676622 912440
rect 674016 907790 674170 912322
rect 676504 907790 676622 912322
rect 674016 907670 676622 907790
rect 670824 474564 673424 474684
rect 670824 470046 670926 474564
rect 673294 470046 673424 474564
rect 670824 469900 673424 470046
rect 674024 469480 676618 469590
rect 674024 465058 674144 469480
rect 676512 465058 676618 469480
rect 674024 464954 676618 465058
rect 670826 464548 673426 464648
rect 670826 460030 670932 464548
rect 673300 460030 673426 464548
rect 670826 459864 673426 460030
rect 680587 459800 681277 459992
rect 688881 459800 688947 474800
rect 7 455645 4843 456093
rect 28653 440800 28719 455800
rect 32933 455546 33623 455800
rect 36323 455607 37013 455799
rect 38503 455546 39593 455800
rect 41008 455654 43618 455758
rect 41008 451042 41142 455654
rect 43508 451042 43618 455654
rect 41008 450950 43618 451042
rect 44202 450528 46812 450636
rect 44202 446104 44290 450528
rect 46690 446104 46812 450528
rect 44202 446016 46812 446104
rect 40994 445596 43604 445704
rect 40994 440984 41122 445596
rect 43488 440984 43604 445596
rect 40994 440896 43604 440984
rect 132600 36323 132792 37013
rect 132580 30762 132848 31674
rect 132600 28653 147600 28719
<< via4 >>
rect 44294 922268 46702 926876
rect 41096 917280 43504 921736
rect 674136 917822 676496 922374
rect 44274 912162 46682 916770
rect 670974 912862 673314 917268
rect 674170 907790 676504 912322
rect 670926 470046 673294 474564
rect 674144 465058 676512 469480
rect 670932 460030 673300 464548
rect 41142 451042 43508 455654
rect 44290 446104 46690 450528
rect 41122 440984 43488 445596
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628240 1018512 640760 1031002
rect 348400 1007147 348466 1008947
rect 348400 1004968 348466 1005617
rect 348400 1000607 348527 1001257
rect 6598 956440 19088 968960
rect 6167 914054 19619 924934
rect 40998 921736 43598 995004
rect 40998 917280 41096 921736
rect 43504 917280 43598 921736
rect 6811 871210 18975 883378
rect 6811 829010 18975 841178
rect 6598 786640 19088 799160
rect 6598 743440 19088 755960
rect 6598 700240 19088 712760
rect 6598 657040 19088 669560
rect 6598 613840 19088 626360
rect 6598 570640 19088 583160
rect 6598 527440 19088 539960
rect 6811 484410 18975 496578
rect 40998 455654 43598 917280
rect 6167 442854 19619 453734
rect 40998 451042 41142 455654
rect 43508 451042 43598 455654
rect 40998 445596 43598 451042
rect 40998 440984 41122 445596
rect 43488 440984 43598 445596
rect 6598 399840 19088 412360
rect 6598 356640 19088 369160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 6598 227040 19088 239560
rect 6598 183840 19088 196360
rect 40998 179300 43598 440984
rect 44198 926876 46798 995004
rect 44198 922268 44294 926876
rect 46702 922268 46798 926876
rect 44198 916770 46798 922268
rect 44198 912162 44274 916770
rect 46682 912162 46798 916770
rect 44198 450528 46798 912162
rect 44198 446104 44290 450528
rect 46690 446104 46798 450528
rect 44198 179300 46798 446104
rect 670820 917268 673420 992714
rect 670820 912862 670974 917268
rect 673314 912862 673420 917268
rect 670820 474564 673420 912862
rect 670820 470046 670926 474564
rect 673294 470046 673420 474564
rect 670820 464548 673420 470046
rect 670820 460030 670932 464548
rect 673300 460030 673420 464548
rect 6811 111610 18975 123778
rect 670820 95156 673420 460030
rect 674020 922374 676620 992714
rect 698512 952840 711002 965360
rect 674020 917822 674136 922374
rect 676496 917822 676620 922374
rect 674020 912322 676620 917822
rect 674020 907790 674170 912322
rect 676504 907790 676620 912322
rect 697980 909666 711432 920546
rect 674020 469480 676620 907790
rect 698512 863640 711002 876160
rect 698624 819822 710788 831990
rect 698512 774440 711002 786960
rect 698512 729440 711002 741960
rect 698512 684440 711002 696960
rect 698512 639240 711002 651760
rect 698512 594240 711002 606760
rect 698512 549040 711002 561560
rect 698624 505222 710788 517390
rect 674020 465058 674144 469480
rect 676512 465058 676620 469480
rect 674020 95156 676620 465058
rect 697980 461866 711432 472746
rect 698624 417022 710788 429190
rect 698512 371840 711002 384360
rect 698512 326640 711002 339160
rect 698512 281640 711002 294160
rect 698512 236640 711002 249160
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use sky130_ef_io__corner_pad  mgmt_corner\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_170 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_374
timestamp 1636986397
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1636986397
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1
timestamp 1636986397
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_174 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_173
timestamp 1636986397
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_172 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_171 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_181
timestamp 1636986397
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1636986397
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1636986397
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1636986397
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1636986397
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_184
timestamp 1636986397
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_183
timestamp 1636986397
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_182
timestamp 1636986397
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_187
timestamp 1636986397
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_189
timestamp 1636986397
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_188
timestamp 1636986397
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1636986397
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1636986397
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_190
timestamp 1636986397
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1636986397
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1636986397
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1636986397
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1636986397
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1636986397
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_198
timestamp 1636986397
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1636986397
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_201
timestamp 1636986397
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_200
timestamp 1636986397
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_199
timestamp 1636986397
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__com_bus_slice_20um  FILLER_204
timestamp 1636986397
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1636986397
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1636986397
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_207
timestamp 1636986397
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_206
timestamp 1636986397
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_205
timestamp 1636986397
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1636986397
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1636986397
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1636986397
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_215
timestamp 1636986397
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1636986397
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1636986397
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_216
timestamp 1636986397
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1636986397
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_218
timestamp 1636986397
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_217
timestamp 1636986397
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 202400 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_221
timestamp 1636986397
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1636986397
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1636986397
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_224
timestamp 1636986397
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_223
timestamp 1636986397
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_222
timestamp 1636986397
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1636986397
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1636986397
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1636986397
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1636986397
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_232
timestamp 1636986397
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1636986397
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1636986397
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_235
timestamp 1636986397
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_234
timestamp 1636986397
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_233
timestamp 1636986397
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 256200 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_238
timestamp 1636986397
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1636986397
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1636986397
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1636986397
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_241
timestamp 1636986397
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_240
timestamp 1636986397
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_239
timestamp 1636986397
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1636986397
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1636986397
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1636986397
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1636986397
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_249
timestamp 1636986397
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1636986397
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_252
timestamp 1636986397
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_251
timestamp 1636986397
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_250
timestamp 1636986397
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1636986397
transform -1 0 311000 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_255
timestamp 1636986397
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_256
timestamp 1636986397
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1636986397
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1636986397
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_258
timestamp 1636986397
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_257
timestamp 1636986397
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1636986397
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1636986397
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1636986397
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1636986397
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_266
timestamp 1636986397
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1636986397
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1636986397
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_269
timestamp 1636986397
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_268
timestamp 1636986397
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_267
timestamp 1636986397
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1636986397
transform -1 0 365800 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_272
timestamp 1636986397
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1636986397
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1636986397
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1636986397
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_275
timestamp 1636986397
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_274
timestamp 1636986397
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_273
timestamp 1636986397
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1636986397
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1636986397
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1636986397
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1636986397
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_283
timestamp 1636986397
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1636986397
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_286
timestamp 1636986397
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_285
timestamp 1636986397
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_284
timestamp 1636986397
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1636986397
transform -1 0 420600 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_289
timestamp 1636986397
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1636986397
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1636986397
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1636986397
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1636986397
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_292
timestamp 1636986397
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_291
timestamp 1636986397
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_290
timestamp 1636986397
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_300
timestamp 1636986397
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1636986397
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1636986397
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1636986397
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1636986397
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_303
timestamp 1636986397
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_302
timestamp 1636986397
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_301
timestamp 1636986397
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1636986397
transform -1 0 475400 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_306
timestamp 1636986397
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_307
timestamp 1636986397
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1636986397
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1636986397
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_309
timestamp 1636986397
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_308
timestamp 1636986397
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1636986397
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1636986397
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1636986397
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1636986397
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1636986397
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_317
timestamp 1636986397
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1636986397
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_320
timestamp 1636986397
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_319
timestamp 1636986397
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_318
timestamp 1636986397
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1636986397
transform -1 0 530200 0 -1 42193
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_323
timestamp 1636986397
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1636986397
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1636986397
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_326
timestamp 1636986397
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_325
timestamp 1636986397
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_324
timestamp 1636986397
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1636986397
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1636986397
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_334
timestamp 1636986397
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1636986397
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1636986397
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1636986397
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1636986397
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_337
timestamp 1636986397
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_336
timestamp 1636986397
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_335
timestamp 1636986397
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_340
timestamp 1636986397
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_342
timestamp 1636986397
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_341
timestamp 1636986397
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1636986397
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1636986397
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1636986397
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1636986397
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1636986397
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_343
timestamp 1636986397
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_351
timestamp 1636986397
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1636986397
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1636986397
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_352
timestamp 1636986397
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_355
timestamp 1636986397
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_354
timestamp 1636986397
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_353
timestamp 1636986397
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1636986397
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1636986397
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_359
timestamp 1636986397
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_358
timestamp 1636986397
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1636986397
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1636986397
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1636986397
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1636986397
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1636986397
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1636986397
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1636986397
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_368
timestamp 1636986397
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_369
timestamp 1636986397
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1636986397
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1636986397
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_371
timestamp 1636986397
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_372
timestamp 1636986397
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_373
timestamp 1636986397
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_370
timestamp 1636986397
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1636986397
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1636986397
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_376
timestamp 1636986397
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1636986397
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1636986397
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_382
timestamp 1636986397
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_381
timestamp 1636986397
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_380
timestamp 1636986397
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform 0 -1 39593 1 0 68000
box 0 -2107 17239 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1636986397
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1636986397
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1636986397
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_608
timestamp 1636986397
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1636986397
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_610
timestamp 1636986397
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_611
timestamp 1636986397
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_612
timestamp 1636986397
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB1
timestamp 1636986397
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1 $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1636986397
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1636986397
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1636986397
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1636986397
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_388
timestamp 1636986397
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_387
timestamp 1636986397
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1636986397
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1636986397
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_389
timestamp 1636986397
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_392
timestamp 1636986397
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_391
timestamp 1636986397
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_390
timestamp 1636986397
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1636986397
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_619
timestamp 1636986397
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_620
timestamp 1636986397
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_621
timestamp 1636986397
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1636986397
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1636986397
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1636986397
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_622
timestamp 1636986397
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1636986397
transform 0 1 675407 -1 0 116000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1636986397
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1636986397
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_397
timestamp 1636986397
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_398
timestamp 1636986397
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_399
timestamp 1636986397
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_400
timestamp 1636986397
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1636986397
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_402
timestamp 1636986397
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_401
timestamp 1636986397
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB2
timestamp 1636986397
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1636986397
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1636986397
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_407
timestamp 1636986397
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_408
timestamp 1636986397
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1636986397
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1636986397
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_629
timestamp 1636986397
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_630
timestamp 1636986397
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1636986397
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1636986397
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_632
timestamp 1636986397
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_631
timestamp 1636986397
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1636986397
transform 0 1 675407 -1 0 161200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_410
timestamp 1636986397
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_409
timestamp 1636986397
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_413
timestamp 1636986397
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_412
timestamp 1636986397
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_411
timestamp 1636986397
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[18\]
timestamp 1636986397
transform 0 -1 42193 1 0 181600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1636986397
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_418
timestamp 1636986397
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_417
timestamp 1636986397
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1636986397
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1636986397
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1636986397
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_638
timestamp 1636986397
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1636986397
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1636986397
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1636986397
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1636986397
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_641
timestamp 1636986397
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1636986397
transform 0 1 675407 -1 0 206200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_420
timestamp 1636986397
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_419
timestamp 1636986397
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_423
timestamp 1636986397
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_422
timestamp 1636986397
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_421
timestamp 1636986397
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[17\]
timestamp 1636986397
transform 0 -1 42193 1 0 224800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1636986397
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_428
timestamp 1636986397
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1636986397
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1636986397
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1636986397
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1636986397
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1636986397
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_648
timestamp 1636986397
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_649
timestamp 1636986397
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1636986397
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_651
timestamp 1636986397
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_650
timestamp 1636986397
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1636986397
transform 0 1 675407 -1 0 251400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_429
timestamp 1636986397
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_430
timestamp 1636986397
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1636986397
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1636986397
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1636986397
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_433
timestamp 1636986397
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_432
timestamp 1636986397
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_431
timestamp 1636986397
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[16\]
timestamp 1636986397
transform 0 -1 42193 1 0 268000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1636986397
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1636986397
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1636986397
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_657
timestamp 1636986397
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_658
timestamp 1636986397
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_659
timestamp 1636986397
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_660
timestamp 1636986397
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1636986397
transform 0 1 675407 -1 0 296400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_440
timestamp 1636986397
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_439
timestamp 1636986397
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_438
timestamp 1636986397
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_443
timestamp 1636986397
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_442
timestamp 1636986397
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_441
timestamp 1636986397
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[15\]
timestamp 1636986397
transform 0 -1 42193 1 0 311200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1636986397
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1636986397
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1636986397
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1636986397
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1636986397
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1636986397
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1636986397
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1636986397
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1636986397
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1636986397
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_669
timestamp 1636986397
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1636986397
transform 0 1 675407 -1 0 341400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_450
timestamp 1636986397
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_449
timestamp 1636986397
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_448
timestamp 1636986397
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_452
timestamp 1636986397
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_451
timestamp 1636986397
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_453
timestamp 1636986397
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[14\]
timestamp 1636986397
transform 0 -1 42193 1 0 354400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1636986397
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1636986397
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1636986397
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1636986397
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1636986397
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1636986397
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1636986397
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1636986397
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1636986397
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1636986397
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_678
timestamp 1636986397
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_679
timestamp 1636986397
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1636986397
transform 0 1 675407 -1 0 386600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_460
timestamp 1636986397
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_459
timestamp 1636986397
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_458
timestamp 1636986397
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_461
timestamp 1636986397
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_463
timestamp 1636986397
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_462
timestamp 1636986397
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[13\]
timestamp 1636986397
transform 0 -1 42193 1 0 397600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1636986397
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1636986397
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1636986397
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1636986397
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1636986397
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1636986397
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1636986397
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_685
timestamp 1636986397
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_686
timestamp 1636986397
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1636986397
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_688
timestamp 1636986397
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1636986397
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_470
timestamp 1636986397
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_469
timestamp 1636986397
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_468
timestamp 1636986397
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_471
timestamp 1636986397
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1636986397
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_473
timestamp 1636986397
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_472
timestamp 1636986397
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user2_vssd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform 0 -1 39593 1 0 440800
box 0 -2177 17187 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1636986397
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1636986397
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1636986397
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1636986397
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1636986397
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_696
timestamp 1636986397
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_695
timestamp 1636986397
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1636986397
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1636986397
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_698
timestamp 1636986397
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_697
timestamp 1636986397
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user1_vssd_lvclamp_pad
timestamp 1636986397
transform 0 1 678007 -1 0 474800
box 0 -2177 17187 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_480
timestamp 1636986397
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_479
timestamp 1636986397
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_478
timestamp 1636986397
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_483
timestamp 1636986397
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_482
timestamp 1636986397
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_481
timestamp 1636986397
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1636986397
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1636986397
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1636986397
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1636986397
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1636986397
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1636986397
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1636986397
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1636986397
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1636986397
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_705
timestamp 1636986397
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1636986397
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_707
timestamp 1636986397
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1636986397
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_488
timestamp 1636986397
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_489
timestamp 1636986397
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_490
timestamp 1636986397
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1636986397
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1636986397
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_493
timestamp 1636986397
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_492
timestamp 1636986397
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_491
timestamp 1636986397
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1636986397
transform 0 -1 42193 1 0 525200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1636986397
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1636986397
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1636986397
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1636986397
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1636986397
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1636986397
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1636986397
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_716
timestamp 1636986397
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1636986397
transform 0 1 675407 -1 0 563800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_500
timestamp 1636986397
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_499
timestamp 1636986397
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_498
timestamp 1636986397
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1636986397
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_503
timestamp 1636986397
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_502
timestamp 1636986397
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_501
timestamp 1636986397
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1636986397
transform 0 -1 42193 1 0 568400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1636986397
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1636986397
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1636986397
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1636986397
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1636986397
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1636986397
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1636986397
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_723
timestamp 1636986397
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_724
timestamp 1636986397
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_510
timestamp 1636986397
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_509
timestamp 1636986397
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_508
timestamp 1636986397
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1636986397
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_513
timestamp 1636986397
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_512
timestamp 1636986397
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_511
timestamp 1636986397
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1636986397
transform 0 -1 42193 1 0 611600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1636986397
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1636986397
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1636986397
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1636986397
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1636986397
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1636986397
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_732
timestamp 1636986397
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1636986397
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_726
timestamp 1636986397
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_725
timestamp 1636986397
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1636986397
transform 0 1 675407 -1 0 609000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_520
timestamp 1636986397
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_519
timestamp 1636986397
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_518
timestamp 1636986397
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1636986397
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_523
timestamp 1636986397
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_522
timestamp 1636986397
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_521
timestamp 1636986397
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1636986397
transform 0 -1 42193 1 0 654800
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1636986397
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1636986397
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1636986397
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1636986397
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1636986397
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1636986397
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1636986397
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1636986397
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_742
timestamp 1636986397
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_735
timestamp 1636986397
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1636986397
transform 0 1 675407 -1 0 654000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1636986397
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_528
timestamp 1636986397
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_529
timestamp 1636986397
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_530
timestamp 1636986397
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1636986397
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_533
timestamp 1636986397
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_532
timestamp 1636986397
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_531
timestamp 1636986397
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1636986397
transform 0 -1 42193 1 0 698000
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1636986397
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1636986397
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1636986397
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1636986397
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1636986397
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_751
timestamp 1636986397
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_745
timestamp 1636986397
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_744
timestamp 1636986397
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1636986397
transform 0 1 675407 -1 0 699200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_539
timestamp 1636986397
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_538
timestamp 1636986397
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1636986397
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1636986397
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_540
timestamp 1636986397
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_543
timestamp 1636986397
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_542
timestamp 1636986397
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_541
timestamp 1636986397
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1636986397
transform 0 -1 42193 1 0 741200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1636986397
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_752
timestamp 1636986397
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1636986397
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1636986397
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1636986397
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1636986397
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1636986397
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_754
timestamp 1636986397
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1636986397
transform 0 1 675407 -1 0 744200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_549
timestamp 1636986397
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_548
timestamp 1636986397
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1636986397
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1636986397
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_550
timestamp 1636986397
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_553
timestamp 1636986397
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_552
timestamp 1636986397
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_551
timestamp 1636986397
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1636986397
transform 0 -1 42193 1 0 784400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1636986397
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1636986397
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_761
timestamp 1636986397
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1636986397
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1636986397
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1636986397
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1636986397
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1636986397
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_763
timestamp 1636986397
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1636986397
transform 0 1 675407 -1 0 789200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_559
timestamp 1636986397
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_558
timestamp 1636986397
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1636986397
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1636986397
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_560
timestamp 1636986397
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_563
timestamp 1636986397
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_562
timestamp 1636986397
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_561
timestamp 1636986397
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1636986397
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1636986397
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1636986397
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1636986397
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1636986397
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1636986397
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1636986397
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1636986397
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_773
timestamp 1636986397
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_772
timestamp 1636986397
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1636986397
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_569
timestamp 1636986397
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_568
timestamp 1636986397
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1636986397
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1636986397
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1636986397
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_573
timestamp 1636986397
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_572
timestamp 1636986397
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_571
timestamp 1636986397
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1636986397
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1636986397
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_778
timestamp 1636986397
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_779
timestamp 1636986397
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_780
timestamp 1636986397
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1636986397
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1636986397
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1636986397
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_782
timestamp 1636986397
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1636986397
transform 0 1 675407 -1 0 878400
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_579
timestamp 1636986397
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_578
timestamp 1636986397
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1636986397
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1636986397
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_580
timestamp 1636986397
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_583
timestamp 1636986397
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_582
timestamp 1636986397
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_581
timestamp 1636986397
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__vccd_lvc_clamped3_pad  user2_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/maglef
timestamp 1636986397
transform 0 -1 39593 1 0 912000
box 0 -2177 17187 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1636986397
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_790
timestamp 1636986397
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_789
timestamp 1636986397
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_788
timestamp 1636986397
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1636986397
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1636986397
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_792
timestamp 1636986397
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_791
timestamp 1636986397
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__vccd_lvc_clamped3_pad  user1_vccd_lvclamp_pad
timestamp 1636986397
transform 0 1 678007 -1 0 922600
box 0 -2177 17187 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1636986397
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1636986397
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_589
timestamp 1636986397
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_588
timestamp 1636986397
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1636986397
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1636986397
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_590
timestamp 1636986397
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_593
timestamp 1636986397
transform 0 -1 39593 1 0 954000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_592
timestamp 1636986397
transform 0 -1 39593 1 0 953000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_591
timestamp 1636986397
transform 0 -1 39593 1 0 951000
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1636986397
transform 0 -1 42193 1 0 954200
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1636986397
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1636986397
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1636986397
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_798
timestamp 1636986397
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_799
timestamp 1636986397
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_800
timestamp 1636986397
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_803
timestamp 1636986397
transform 0 1 678007 -1 0 971600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_801
timestamp 1636986397
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[14\]
timestamp 1636986397
transform 0 1 675407 -1 0 967600
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_600
timestamp 1636986397
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1636986397
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_598
timestamp 1636986397
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1636986397
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1636986397
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_604
timestamp 1636986397
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_603
timestamp 1636986397
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_602
timestamp 1636986397
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_601
timestamp 1636986397
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1636986397
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1636986397
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1636986397
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1636986397
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1636986397
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1636986397
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1636986397
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1636986397
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1636986397
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13
timestamp 1636986397
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1636986397
transform 1 0 76000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1636986397
transform 1 0 75800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_14
timestamp 1636986397
transform 1 0 74800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1636986397
transform 1 0 76200 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1636986397
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1636986397
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1636986397
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1636986397
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1636986397
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1636986397
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1636986397
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1636986397
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_27
timestamp 1636986397
transform 1 0 126200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_26
timestamp 1636986397
transform 1 0 124200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1636986397
transform 1 0 127400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1636986397
transform 1 0 127200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1636986397
transform 1 0 127600 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1636986397
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1636986397
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1636986397
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1636986397
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1636986397
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1636986397
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1636986397
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1636986397
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1636986397
transform 1 0 178800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1636986397
transform 1 0 178600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_40
timestamp 1636986397
transform 1 0 177600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_39
timestamp 1636986397
transform 1 0 175600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1636986397
transform 1 0 179000 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1636986397
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1636986397
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1636986397
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1636986397
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1636986397
transform 1 0 223000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1636986397
transform 1 0 219000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1636986397
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1636986397
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_52
timestamp 1636986397
transform 1 0 227000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1636986397
transform 1 0 230200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1636986397
transform 1 0 230000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1636986397
transform 1 0 229000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1636986397
transform 1 0 230400 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1636986397
transform 1 0 250400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1636986397
transform 1 0 246400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1636986397
transform 1 0 266400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1636986397
transform 1 0 262400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1636986397
transform 1 0 258400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1636986397
transform 1 0 254400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1636986397
transform 1 0 274400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1636986397
transform 1 0 270400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1636986397
transform 1 0 281800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1636986397
transform 1 0 281600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1636986397
transform 1 0 281400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1636986397
transform 1 0 280400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1636986397
transform 1 0 278400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1636986397
transform 1 0 282000 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1636986397
transform 1 0 310000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1636986397
transform 1 0 306000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1636986397
transform 1 0 302000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1636986397
transform 1 0 298000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1636986397
transform 1 0 322000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1636986397
transform 1 0 318000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1636986397
transform 1 0 314000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1636986397
transform 1 0 326000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1636986397
transform 1 0 333200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1636986397
transform 1 0 333000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_80
timestamp 1636986397
transform 1 0 332000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_79
timestamp 1636986397
transform 1 0 330000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1636986397
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB3
timestamp 1636986397
transform 1 0 349400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1636986397
transform 1 0 348400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1636986397
transform 1 0 354400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1636986397
transform 1 0 350400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1636986397
transform 1 0 358400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1636986397
transform 1 0 362400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1636986397
transform 1 0 366400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1636986397
transform 1 0 370400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1636986397
transform 1 0 374400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_93
timestamp 1636986397
transform 1 0 378400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_96
timestamp 1636986397
transform 1 0 383600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1636986397
transform 1 0 383400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_94
timestamp 1636986397
transform 1 0 382400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[18\]
timestamp 1636986397
transform 1 0 383800 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1636986397
transform 1 0 411800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1636986397
transform 1 0 407800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1636986397
transform 1 0 403800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1636986397
transform 1 0 399800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1636986397
transform 1 0 419800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1636986397
transform 1 0 415800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1636986397
transform 1 0 423800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1636986397
transform 1 0 427800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1636986397
transform 1 0 431800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_107
timestamp 1636986397
transform 1 0 435800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_108
timestamp 1636986397
transform 1 0 439800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_109
timestamp 1636986397
transform 1 0 443800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_110
timestamp 1636986397
transform 1 0 447800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1636986397
transform 1 0 451800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1636986397
transform 1 0 455800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1636986397
transform 1 0 459800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1636986397
transform 1 0 463800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1636986397
transform 1 0 467800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1636986397
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_119
timestamp 1636986397
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_120
timestamp 1636986397
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_121
timestamp 1636986397
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_122
timestamp 1636986397
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_116
timestamp 1636986397
transform 1 0 471800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[17\]
timestamp 1636986397
transform 1 0 472800 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1636986397
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_124
timestamp 1636986397
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1636986397
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_126
timestamp 1636986397
transform 1 0 520800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_129
timestamp 1636986397
transform 1 0 524000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_128
timestamp 1636986397
transform 1 0 523800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_127
timestamp 1636986397
transform 1 0 522800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[16\]
timestamp 1636986397
transform 1 0 524200 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_133
timestamp 1636986397
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1636986397
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1636986397
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1636986397
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1636986397
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_134
timestamp 1636986397
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1636986397
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_137
timestamp 1636986397
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_142
timestamp 1636986397
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_141
timestamp 1636986397
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_140
timestamp 1636986397
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_139
timestamp 1636986397
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1636986397
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1636986397
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_148
timestamp 1636986397
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_147
timestamp 1636986397
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_146
timestamp 1636986397
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1636986397
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1636986397
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_150
timestamp 1636986397
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_149
timestamp 1636986397
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_152
timestamp 1636986397
transform 1 0 622600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_155
timestamp 1636986397
transform 1 0 625800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_154
timestamp 1636986397
transform 1 0 625600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_153
timestamp 1636986397
transform 1 0 624600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[15\]
timestamp 1636986397
transform 1 0 626000 0 1 995407
box -32 0 16032 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1636986397
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1636986397
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_159
timestamp 1636986397
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_160
timestamp 1636986397
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_161
timestamp 1636986397
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_162
timestamp 1636986397
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_163
timestamp 1636986397
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1636986397
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_165
timestamp 1636986397
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_808
timestamp 1636986397
transform 0 1 678007 -1 0 991600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1636986397
transform 0 1 678007 -1 0 987600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1636986397
transform 0 1 678007 -1 0 983600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1636986397
transform 0 1 678007 -1 0 979600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1636986397
transform 0 1 678007 -1 0 975600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_809
timestamp 1636986397
transform 0 1 678007 -1 0 995600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_811
timestamp 1636986397
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_810
timestamp 1636986397
transform 0 1 678007 -1 0 996600
box 0 0 1000 39593
use sky130_ef_io__corner_pad  user1_corner
timestamp 1636986397
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1636986397
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1636986397
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_167
timestamp 1636986397
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_166
timestamp 1636986397
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 0 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 1 nsew signal tristate
rlabel metal2 s 194043 41713 194099 42193 6 por
port 2 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 3 nsew signal tristate
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 4 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 5 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 6 nsew signal input
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 7 nsew signal tristate
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 8 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 9 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 10 nsew signal input
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 11 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 12 nsew signal tristate
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 13 nsew signal input
rlabel metal2 s 412243 41713 412299 42193 6 flash_io0_ieb_core
port 14 nsew signal input
rlabel metal2 s 419695 41713 419751 42193 6 flash_io0_oeb_core
port 15 nsew signal input
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 16 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 17 nsew signal tristate
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 18 nsew signal input
rlabel metal2 s 467043 41713 467099 42193 6 flash_io1_ieb_core
port 19 nsew signal input
rlabel metal2 s 474495 41713 474551 42193 6 flash_io1_oeb_core
port 20 nsew signal input
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 21 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 22 nsew signal tristate
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 23 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 24 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 25 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 26 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 27 nsew signal input
rlabel metal5 s 6167 70054 19619 80934 6 vccd_pad
port 28 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18975 6 vdda_pad
port 29 nsew signal bidirectional
rlabel metal5 s 6811 111610 18975 123778 6 vddio_pad
port 30 nsew signal bidirectional
rlabel metal5 s 6811 871210 18975 883378 6 vddio_pad2
port 31 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18975 6 vssa_pad
port 32 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19619 6 vssd_pad
port 33 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18975 6 vssio_pad
port 34 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030788 6 vssio_pad2
port 35 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113780 6 mprj_io[0]
port 36 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 37 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 38 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 39 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 40 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 41 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 42 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 43 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 44 nsew signal input
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 45 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 46 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 47 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 48 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 49 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 50 nsew signal tristate
rlabel metal2 s 675407 686611 675887 686667 6 mprj_analog_io[3]
port 51 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696980 6 mprj_io[10]
port 52 nsew signal bidirectional
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 53 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 54 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 55 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 56 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 57 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 58 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 59 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 60 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 61 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 62 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 63 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 64 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 65 nsew signal input
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 66 nsew signal tristate
rlabel metal2 s 675407 731611 675887 731667 6 mprj_analog_io[4]
port 67 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741980 6 mprj_io[11]
port 68 nsew signal bidirectional
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 69 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 70 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 71 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 72 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 73 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 74 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 75 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 76 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 77 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 78 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 79 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 80 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 81 nsew signal input
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 82 nsew signal tristate
rlabel metal2 s 675407 776611 675887 776667 6 mprj_analog_io[5]
port 83 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786980 6 mprj_io[12]
port 84 nsew signal bidirectional
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 85 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 86 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 87 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 88 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 89 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 90 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 91 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 92 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 93 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 94 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 95 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 96 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 97 nsew signal input
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 98 nsew signal tristate
rlabel metal2 s 675407 865811 675887 865867 6 mprj_analog_io[6]
port 99 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876180 6 mprj_io[13]
port 100 nsew signal bidirectional
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 101 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 102 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 103 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 104 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 105 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 106 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 107 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 108 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 109 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 110 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 111 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 112 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 113 nsew signal input
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 114 nsew signal tristate
rlabel metal2 s 675407 955011 675887 955067 6 mprj_analog_io[7]
port 115 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965380 6 mprj_io[14]
port 116 nsew signal bidirectional
rlabel metal2 s 675407 957403 675887 957459 6 mprj_io_analog_en[14]
port 117 nsew signal input
rlabel metal2 s 675407 958691 675887 958747 6 mprj_io_analog_pol[14]
port 118 nsew signal input
rlabel metal2 s 675407 961727 675887 961783 6 mprj_io_analog_sel[14]
port 119 nsew signal input
rlabel metal2 s 675407 958047 675887 958103 6 mprj_io_dm[42]
port 120 nsew signal input
rlabel metal2 s 675407 956207 675887 956263 6 mprj_io_dm[43]
port 121 nsew signal input
rlabel metal2 s 675407 962371 675887 962427 6 mprj_io_dm[44]
port 122 nsew signal input
rlabel metal2 s 675407 963015 675887 963071 6 mprj_io_holdover[14]
port 123 nsew signal input
rlabel metal2 s 675407 966051 675887 966107 6 mprj_io_ib_mode_sel[14]
port 124 nsew signal input
rlabel metal2 s 675407 959243 675887 959299 6 mprj_io_inp_dis[14]
port 125 nsew signal input
rlabel metal2 s 675407 966695 675887 966751 6 mprj_io_oeb[14]
port 126 nsew signal input
rlabel metal2 s 675407 963567 675887 963623 6 mprj_io_out[14]
port 127 nsew signal input
rlabel metal2 s 675407 954367 675887 954423 6 mprj_io_slow_sel[14]
port 128 nsew signal input
rlabel metal2 s 675407 965407 675887 965463 6 mprj_io_vtrip_sel[14]
port 129 nsew signal input
rlabel metal2 s 675407 952527 675887 952583 6 mprj_io_in[14]
port 130 nsew signal tristate
rlabel metal2 s 638533 995407 638589 995887 6 mprj_analog_io[8]
port 131 nsew signal bidirectional
rlabel metal5 s 628220 1018512 640760 1031002 6 mprj_io[15]
port 132 nsew signal bidirectional
rlabel metal2 s 636141 995407 636197 995887 6 mprj_io_analog_en[15]
port 133 nsew signal input
rlabel metal2 s 634853 995407 634909 995887 6 mprj_io_analog_pol[15]
port 134 nsew signal input
rlabel metal2 s 631817 995407 631873 995887 6 mprj_io_analog_sel[15]
port 135 nsew signal input
rlabel metal2 s 635497 995407 635553 995887 6 mprj_io_dm[45]
port 136 nsew signal input
rlabel metal2 s 637337 995407 637393 995887 6 mprj_io_dm[46]
port 137 nsew signal input
rlabel metal2 s 631173 995407 631229 995887 6 mprj_io_dm[47]
port 138 nsew signal input
rlabel metal2 s 630529 995407 630585 995887 6 mprj_io_holdover[15]
port 139 nsew signal input
rlabel metal2 s 627493 995407 627549 995887 6 mprj_io_ib_mode_sel[15]
port 140 nsew signal input
rlabel metal2 s 634301 995407 634357 995887 6 mprj_io_inp_dis[15]
port 141 nsew signal input
rlabel metal2 s 626849 995407 626905 995887 6 mprj_io_oeb[15]
port 142 nsew signal input
rlabel metal2 s 629977 995407 630033 995887 6 mprj_io_out[15]
port 143 nsew signal input
rlabel metal2 s 639177 995407 639233 995887 6 mprj_io_slow_sel[15]
port 144 nsew signal input
rlabel metal2 s 628137 995407 628193 995887 6 mprj_io_vtrip_sel[15]
port 145 nsew signal input
rlabel metal2 s 641017 995407 641073 995887 6 mprj_io_in[15]
port 146 nsew signal tristate
rlabel metal2 s 536733 995407 536789 995887 6 mprj_analog_io[9]
port 147 nsew signal bidirectional
rlabel metal5 s 526420 1018512 538960 1031002 6 mprj_io[16]
port 148 nsew signal bidirectional
rlabel metal2 s 534341 995407 534397 995887 6 mprj_io_analog_en[16]
port 149 nsew signal input
rlabel metal2 s 533053 995407 533109 995887 6 mprj_io_analog_pol[16]
port 150 nsew signal input
rlabel metal2 s 530017 995407 530073 995887 6 mprj_io_analog_sel[16]
port 151 nsew signal input
rlabel metal2 s 533697 995407 533753 995887 6 mprj_io_dm[48]
port 152 nsew signal input
rlabel metal2 s 535537 995407 535593 995887 6 mprj_io_dm[49]
port 153 nsew signal input
rlabel metal2 s 529373 995407 529429 995887 6 mprj_io_dm[50]
port 154 nsew signal input
rlabel metal2 s 528729 995407 528785 995887 6 mprj_io_holdover[16]
port 155 nsew signal input
rlabel metal2 s 525693 995407 525749 995887 6 mprj_io_ib_mode_sel[16]
port 156 nsew signal input
rlabel metal2 s 532501 995407 532557 995887 6 mprj_io_inp_dis[16]
port 157 nsew signal input
rlabel metal2 s 525049 995407 525105 995887 6 mprj_io_oeb[16]
port 158 nsew signal input
rlabel metal2 s 528177 995407 528233 995887 6 mprj_io_out[16]
port 159 nsew signal input
rlabel metal2 s 537377 995407 537433 995887 6 mprj_io_slow_sel[16]
port 160 nsew signal input
rlabel metal2 s 526337 995407 526393 995887 6 mprj_io_vtrip_sel[16]
port 161 nsew signal input
rlabel metal2 s 539217 995407 539273 995887 6 mprj_io_in[16]
port 162 nsew signal tristate
rlabel metal2 s 485333 995407 485389 995887 6 mprj_analog_io[10]
port 163 nsew signal bidirectional
rlabel metal5 s 475020 1018512 487560 1031002 6 mprj_io[17]
port 164 nsew signal bidirectional
rlabel metal2 s 482941 995407 482997 995887 6 mprj_io_analog_en[17]
port 165 nsew signal input
rlabel metal2 s 481653 995407 481709 995887 6 mprj_io_analog_pol[17]
port 166 nsew signal input
rlabel metal2 s 478617 995407 478673 995887 6 mprj_io_analog_sel[17]
port 167 nsew signal input
rlabel metal2 s 482297 995407 482353 995887 6 mprj_io_dm[51]
port 168 nsew signal input
rlabel metal2 s 484137 995407 484193 995887 6 mprj_io_dm[52]
port 169 nsew signal input
rlabel metal2 s 477973 995407 478029 995887 6 mprj_io_dm[53]
port 170 nsew signal input
rlabel metal2 s 477329 995407 477385 995887 6 mprj_io_holdover[17]
port 171 nsew signal input
rlabel metal2 s 474293 995407 474349 995887 6 mprj_io_ib_mode_sel[17]
port 172 nsew signal input
rlabel metal2 s 481101 995407 481157 995887 6 mprj_io_inp_dis[17]
port 173 nsew signal input
rlabel metal2 s 473649 995407 473705 995887 6 mprj_io_oeb[17]
port 174 nsew signal input
rlabel metal2 s 476777 995407 476833 995887 6 mprj_io_out[17]
port 175 nsew signal input
rlabel metal2 s 485977 995407 486033 995887 6 mprj_io_slow_sel[17]
port 176 nsew signal input
rlabel metal2 s 474937 995407 474993 995887 6 mprj_io_vtrip_sel[17]
port 177 nsew signal input
rlabel metal2 s 487817 995407 487873 995887 6 mprj_io_in[17]
port 178 nsew signal tristate
rlabel metal2 s 396333 995407 396389 995887 6 mprj_analog_io[11]
port 179 nsew signal bidirectional
rlabel metal5 s 386020 1018512 398560 1031002 6 mprj_io[18]
port 180 nsew signal bidirectional
rlabel metal2 s 393941 995407 393997 995887 6 mprj_io_analog_en[18]
port 181 nsew signal input
rlabel metal2 s 392653 995407 392709 995887 6 mprj_io_analog_pol[18]
port 182 nsew signal input
rlabel metal2 s 389617 995407 389673 995887 6 mprj_io_analog_sel[18]
port 183 nsew signal input
rlabel metal2 s 393297 995407 393353 995887 6 mprj_io_dm[54]
port 184 nsew signal input
rlabel metal2 s 395137 995407 395193 995887 6 mprj_io_dm[55]
port 185 nsew signal input
rlabel metal2 s 388973 995407 389029 995887 6 mprj_io_dm[56]
port 186 nsew signal input
rlabel metal2 s 388329 995407 388385 995887 6 mprj_io_holdover[18]
port 187 nsew signal input
rlabel metal2 s 385293 995407 385349 995887 6 mprj_io_ib_mode_sel[18]
port 188 nsew signal input
rlabel metal2 s 392101 995407 392157 995887 6 mprj_io_inp_dis[18]
port 189 nsew signal input
rlabel metal2 s 384649 995407 384705 995887 6 mprj_io_oeb[18]
port 190 nsew signal input
rlabel metal2 s 387777 995407 387833 995887 6 mprj_io_out[18]
port 191 nsew signal input
rlabel metal2 s 396977 995407 397033 995887 6 mprj_io_slow_sel[18]
port 192 nsew signal input
rlabel metal2 s 385937 995407 385993 995887 6 mprj_io_vtrip_sel[18]
port 193 nsew signal input
rlabel metal2 s 398817 995407 398873 995887 6 mprj_io_in[18]
port 194 nsew signal tristate
rlabel metal5 s 698512 146440 711002 158980 6 mprj_io[1]
port 195 nsew signal bidirectional
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 196 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 197 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 198 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 199 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 200 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 201 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 202 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 203 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 204 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 205 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 206 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 207 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 208 nsew signal input
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 209 nsew signal tristate
rlabel metal5 s 698512 191440 711002 203980 6 mprj_io[2]
port 210 nsew signal bidirectional
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 211 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 212 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 213 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 214 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 215 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 216 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 217 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 218 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 219 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 220 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 221 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 222 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 223 nsew signal input
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 224 nsew signal tristate
rlabel metal5 s 698512 236640 711002 249180 6 mprj_io[3]
port 225 nsew signal bidirectional
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 226 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 227 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 228 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 229 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 230 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 231 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 232 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 233 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 234 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 235 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 236 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 237 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 238 nsew signal input
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 239 nsew signal tristate
rlabel metal5 s 698512 281640 711002 294180 6 mprj_io[4]
port 240 nsew signal bidirectional
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 241 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 242 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 243 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 244 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 245 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 246 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 247 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 248 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 249 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 250 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 251 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 252 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 253 nsew signal input
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 254 nsew signal tristate
rlabel metal5 s 698512 326640 711002 339180 6 mprj_io[5]
port 255 nsew signal bidirectional
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 256 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 257 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 258 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 259 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 260 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 261 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 262 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 263 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 264 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 265 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 266 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 267 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 268 nsew signal input
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 269 nsew signal tristate
rlabel metal5 s 698512 371840 711002 384380 6 mprj_io[6]
port 270 nsew signal bidirectional
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 271 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 272 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 273 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 274 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 275 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 276 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 277 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 278 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 279 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 280 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 281 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 282 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 283 nsew signal input
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 284 nsew signal tristate
rlabel metal2 s 675407 551211 675887 551267 6 mprj_analog_io[0]
port 285 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561580 6 mprj_io[7]
port 286 nsew signal bidirectional
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 287 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 288 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 289 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 290 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 291 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 292 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 293 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 294 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 295 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 296 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 297 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 298 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 299 nsew signal input
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 300 nsew signal tristate
rlabel metal2 s 675407 596411 675887 596467 6 mprj_analog_io[1]
port 301 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606780 6 mprj_io[8]
port 302 nsew signal bidirectional
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 303 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 304 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 305 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 306 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 307 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 308 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 309 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 310 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 311 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 312 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 313 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 314 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 315 nsew signal input
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 316 nsew signal tristate
rlabel metal2 s 675407 641411 675887 641467 6 mprj_analog_io[2]
port 317 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651780 6 mprj_io[9]
port 318 nsew signal bidirectional
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 319 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 320 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 321 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 322 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 323 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 324 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 325 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 326 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 327 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 328 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 329 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 330 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 331 nsew signal input
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 332 nsew signal tristate
rlabel metal2 s 294533 995407 294589 995887 6 mprj_analog_io[12]
port 333 nsew signal bidirectional
rlabel metal5 s 284220 1018512 296760 1031002 6 mprj_io[19]
port 334 nsew signal bidirectional
rlabel metal2 s 292141 995407 292197 995887 6 mprj_io_analog_en[19]
port 335 nsew signal input
rlabel metal2 s 290853 995407 290909 995887 6 mprj_io_analog_pol[19]
port 336 nsew signal input
rlabel metal2 s 287817 995407 287873 995887 6 mprj_io_analog_sel[19]
port 337 nsew signal input
rlabel metal2 s 291497 995407 291553 995887 6 mprj_io_dm[57]
port 338 nsew signal input
rlabel metal2 s 293337 995407 293393 995887 6 mprj_io_dm[58]
port 339 nsew signal input
rlabel metal2 s 287173 995407 287229 995887 6 mprj_io_dm[59]
port 340 nsew signal input
rlabel metal2 s 286529 995407 286585 995887 6 mprj_io_holdover[19]
port 341 nsew signal input
rlabel metal2 s 283493 995407 283549 995887 6 mprj_io_ib_mode_sel[19]
port 342 nsew signal input
rlabel metal2 s 290301 995407 290357 995887 6 mprj_io_inp_dis[19]
port 343 nsew signal input
rlabel metal2 s 282849 995407 282905 995887 6 mprj_io_oeb[19]
port 344 nsew signal input
rlabel metal2 s 285977 995407 286033 995887 6 mprj_io_out[19]
port 345 nsew signal input
rlabel metal2 s 295177 995407 295233 995887 6 mprj_io_slow_sel[19]
port 346 nsew signal input
rlabel metal2 s 284137 995407 284193 995887 6 mprj_io_vtrip_sel[19]
port 347 nsew signal input
rlabel metal2 s 297017 995407 297073 995887 6 mprj_io_in[19]
port 348 nsew signal tristate
rlabel metal2 s 41713 624133 42193 624189 6 mprj_analog_io[22]
port 349 nsew signal bidirectional
rlabel metal5 s 6598 613820 19088 626360 6 mprj_io[29]
port 350 nsew signal bidirectional
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[29]
port 351 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[29]
port 352 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[29]
port 353 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[87]
port 354 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[88]
port 355 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[89]
port 356 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[29]
port 357 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[29]
port 358 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[29]
port 359 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[29]
port 360 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[29]
port 361 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[29]
port 362 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[29]
port 363 nsew signal input
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[29]
port 364 nsew signal tristate
rlabel metal2 s 41713 580933 42193 580989 6 mprj_analog_io[23]
port 365 nsew signal bidirectional
rlabel metal5 s 6598 570620 19088 583160 6 mprj_io[30]
port 366 nsew signal bidirectional
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[30]
port 367 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[30]
port 368 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[30]
port 369 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[90]
port 370 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[91]
port 371 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[92]
port 372 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[30]
port 373 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[30]
port 374 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[30]
port 375 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[30]
port 376 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[30]
port 377 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[30]
port 378 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[30]
port 379 nsew signal input
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[30]
port 380 nsew signal tristate
rlabel metal2 s 41713 537733 42193 537789 6 mprj_analog_io[24]
port 381 nsew signal bidirectional
rlabel metal5 s 6598 527420 19088 539960 6 mprj_io[31]
port 382 nsew signal bidirectional
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[31]
port 383 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[31]
port 384 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[31]
port 385 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[93]
port 386 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[94]
port 387 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[95]
port 388 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[31]
port 389 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[31]
port 390 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[31]
port 391 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[31]
port 392 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[31]
port 393 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[31]
port 394 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[31]
port 395 nsew signal input
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[31]
port 396 nsew signal tristate
rlabel metal2 s 41713 410133 42193 410189 6 mprj_analog_io[25]
port 397 nsew signal bidirectional
rlabel metal5 s 6598 399820 19088 412360 6 mprj_io[32]
port 398 nsew signal bidirectional
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[32]
port 399 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[32]
port 400 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[32]
port 401 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[96]
port 402 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[97]
port 403 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[98]
port 404 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[32]
port 405 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[32]
port 406 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[32]
port 407 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[32]
port 408 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[32]
port 409 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[32]
port 410 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[32]
port 411 nsew signal input
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[32]
port 412 nsew signal tristate
rlabel metal2 s 41713 366933 42193 366989 6 mprj_analog_io[26]
port 413 nsew signal bidirectional
rlabel metal5 s 6598 356620 19088 369160 6 mprj_io[33]
port 414 nsew signal bidirectional
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[33]
port 415 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[33]
port 416 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[33]
port 417 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[100]
port 418 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[101]
port 419 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[99]
port 420 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[33]
port 421 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[33]
port 422 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[33]
port 423 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[33]
port 424 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[33]
port 425 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[33]
port 426 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[33]
port 427 nsew signal input
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[33]
port 428 nsew signal tristate
rlabel metal2 s 41713 323733 42193 323789 6 mprj_analog_io[27]
port 429 nsew signal bidirectional
rlabel metal5 s 6598 313420 19088 325960 6 mprj_io[34]
port 430 nsew signal bidirectional
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[34]
port 431 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[34]
port 432 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[34]
port 433 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[102]
port 434 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[103]
port 435 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[104]
port 436 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[34]
port 437 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[34]
port 438 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[34]
port 439 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[34]
port 440 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[34]
port 441 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[34]
port 442 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[34]
port 443 nsew signal input
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[34]
port 444 nsew signal tristate
rlabel metal2 s 41713 280533 42193 280589 6 mprj_analog_io[28]
port 445 nsew signal bidirectional
rlabel metal5 s 6598 270220 19088 282760 6 mprj_io[35]
port 446 nsew signal bidirectional
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[35]
port 447 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[35]
port 448 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[35]
port 449 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[105]
port 450 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[106]
port 451 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[107]
port 452 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[35]
port 453 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[35]
port 454 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[35]
port 455 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[35]
port 456 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[35]
port 457 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[35]
port 458 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[35]
port 459 nsew signal input
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[35]
port 460 nsew signal tristate
rlabel metal5 s 6598 227020 19088 239560 6 mprj_io[36]
port 461 nsew signal bidirectional
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[36]
port 462 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[36]
port 463 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[36]
port 464 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[108]
port 465 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[109]
port 466 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[110]
port 467 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[36]
port 468 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[36]
port 469 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[36]
port 470 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[36]
port 471 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[36]
port 472 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[36]
port 473 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[36]
port 474 nsew signal input
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[36]
port 475 nsew signal tristate
rlabel metal5 s 6598 183820 19088 196360 6 mprj_io[37]
port 476 nsew signal bidirectional
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[37]
port 477 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[37]
port 478 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[37]
port 479 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[111]
port 480 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[112]
port 481 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[113]
port 482 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[37]
port 483 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[37]
port 484 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[37]
port 485 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[37]
port 486 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[37]
port 487 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[37]
port 488 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[37]
port 489 nsew signal input
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[37]
port 490 nsew signal tristate
rlabel metal2 s 242933 995407 242989 995887 6 mprj_analog_io[13]
port 491 nsew signal bidirectional
rlabel metal5 s 232620 1018512 245160 1031002 6 mprj_io[20]
port 492 nsew signal bidirectional
rlabel metal2 s 240541 995407 240597 995887 6 mprj_io_analog_en[20]
port 493 nsew signal input
rlabel metal2 s 239253 995407 239309 995887 6 mprj_io_analog_pol[20]
port 494 nsew signal input
rlabel metal2 s 236217 995407 236273 995887 6 mprj_io_analog_sel[20]
port 495 nsew signal input
rlabel metal2 s 239897 995407 239953 995887 6 mprj_io_dm[60]
port 496 nsew signal input
rlabel metal2 s 241737 995407 241793 995887 6 mprj_io_dm[61]
port 497 nsew signal input
rlabel metal2 s 235573 995407 235629 995887 6 mprj_io_dm[62]
port 498 nsew signal input
rlabel metal2 s 234929 995407 234985 995887 6 mprj_io_holdover[20]
port 499 nsew signal input
rlabel metal2 s 231893 995407 231949 995887 6 mprj_io_ib_mode_sel[20]
port 500 nsew signal input
rlabel metal2 s 238701 995407 238757 995887 6 mprj_io_inp_dis[20]
port 501 nsew signal input
rlabel metal2 s 231249 995407 231305 995887 6 mprj_io_oeb[20]
port 502 nsew signal input
rlabel metal2 s 234377 995407 234433 995887 6 mprj_io_out[20]
port 503 nsew signal input
rlabel metal2 s 243577 995407 243633 995887 6 mprj_io_slow_sel[20]
port 504 nsew signal input
rlabel metal2 s 232537 995407 232593 995887 6 mprj_io_vtrip_sel[20]
port 505 nsew signal input
rlabel metal2 s 245417 995407 245473 995887 6 mprj_io_in[20]
port 506 nsew signal tristate
rlabel metal2 s 191533 995407 191589 995887 6 mprj_analog_io[14]
port 507 nsew signal bidirectional
rlabel metal5 s 181220 1018512 193760 1031002 6 mprj_io[21]
port 508 nsew signal bidirectional
rlabel metal2 s 189141 995407 189197 995887 6 mprj_io_analog_en[21]
port 509 nsew signal input
rlabel metal2 s 187853 995407 187909 995887 6 mprj_io_analog_pol[21]
port 510 nsew signal input
rlabel metal2 s 184817 995407 184873 995887 6 mprj_io_analog_sel[21]
port 511 nsew signal input
rlabel metal2 s 188497 995407 188553 995887 6 mprj_io_dm[63]
port 512 nsew signal input
rlabel metal2 s 190337 995407 190393 995887 6 mprj_io_dm[64]
port 513 nsew signal input
rlabel metal2 s 184173 995407 184229 995887 6 mprj_io_dm[65]
port 514 nsew signal input
rlabel metal2 s 183529 995407 183585 995887 6 mprj_io_holdover[21]
port 515 nsew signal input
rlabel metal2 s 180493 995407 180549 995887 6 mprj_io_ib_mode_sel[21]
port 516 nsew signal input
rlabel metal2 s 187301 995407 187357 995887 6 mprj_io_inp_dis[21]
port 517 nsew signal input
rlabel metal2 s 179849 995407 179905 995887 6 mprj_io_oeb[21]
port 518 nsew signal input
rlabel metal2 s 182977 995407 183033 995887 6 mprj_io_out[21]
port 519 nsew signal input
rlabel metal2 s 192177 995407 192233 995887 6 mprj_io_slow_sel[21]
port 520 nsew signal input
rlabel metal2 s 181137 995407 181193 995887 6 mprj_io_vtrip_sel[21]
port 521 nsew signal input
rlabel metal2 s 194017 995407 194073 995887 6 mprj_io_in[21]
port 522 nsew signal tristate
rlabel metal2 s 140133 995407 140189 995887 6 mprj_analog_io[15]
port 523 nsew signal bidirectional
rlabel metal5 s 129820 1018512 142360 1031002 6 mprj_io[22]
port 524 nsew signal bidirectional
rlabel metal2 s 137741 995407 137797 995887 6 mprj_io_analog_en[22]
port 525 nsew signal input
rlabel metal2 s 136453 995407 136509 995887 6 mprj_io_analog_pol[22]
port 526 nsew signal input
rlabel metal2 s 133417 995407 133473 995887 6 mprj_io_analog_sel[22]
port 527 nsew signal input
rlabel metal2 s 137097 995407 137153 995887 6 mprj_io_dm[66]
port 528 nsew signal input
rlabel metal2 s 138937 995407 138993 995887 6 mprj_io_dm[67]
port 529 nsew signal input
rlabel metal2 s 132773 995407 132829 995887 6 mprj_io_dm[68]
port 530 nsew signal input
rlabel metal2 s 132129 995407 132185 995887 6 mprj_io_holdover[22]
port 531 nsew signal input
rlabel metal2 s 129093 995407 129149 995887 6 mprj_io_ib_mode_sel[22]
port 532 nsew signal input
rlabel metal2 s 135901 995407 135957 995887 6 mprj_io_inp_dis[22]
port 533 nsew signal input
rlabel metal2 s 128449 995407 128505 995887 6 mprj_io_oeb[22]
port 534 nsew signal input
rlabel metal2 s 131577 995407 131633 995887 6 mprj_io_out[22]
port 535 nsew signal input
rlabel metal2 s 140777 995407 140833 995887 6 mprj_io_slow_sel[22]
port 536 nsew signal input
rlabel metal2 s 129737 995407 129793 995887 6 mprj_io_vtrip_sel[22]
port 537 nsew signal input
rlabel metal2 s 142617 995407 142673 995887 6 mprj_io_in[22]
port 538 nsew signal tristate
rlabel metal2 s 88733 995407 88789 995887 6 mprj_analog_io[16]
port 539 nsew signal bidirectional
rlabel metal5 s 78420 1018512 90960 1031002 6 mprj_io[23]
port 540 nsew signal bidirectional
rlabel metal2 s 86341 995407 86397 995887 6 mprj_io_analog_en[23]
port 541 nsew signal input
rlabel metal2 s 85053 995407 85109 995887 6 mprj_io_analog_pol[23]
port 542 nsew signal input
rlabel metal2 s 82017 995407 82073 995887 6 mprj_io_analog_sel[23]
port 543 nsew signal input
rlabel metal2 s 85697 995407 85753 995887 6 mprj_io_dm[69]
port 544 nsew signal input
rlabel metal2 s 87537 995407 87593 995887 6 mprj_io_dm[70]
port 545 nsew signal input
rlabel metal2 s 81373 995407 81429 995887 6 mprj_io_dm[71]
port 546 nsew signal input
rlabel metal2 s 80729 995407 80785 995887 6 mprj_io_holdover[23]
port 547 nsew signal input
rlabel metal2 s 77693 995407 77749 995887 6 mprj_io_ib_mode_sel[23]
port 548 nsew signal input
rlabel metal2 s 84501 995407 84557 995887 6 mprj_io_inp_dis[23]
port 549 nsew signal input
rlabel metal2 s 77049 995407 77105 995887 6 mprj_io_oeb[23]
port 550 nsew signal input
rlabel metal2 s 80177 995407 80233 995887 6 mprj_io_out[23]
port 551 nsew signal input
rlabel metal2 s 89377 995407 89433 995887 6 mprj_io_slow_sel[23]
port 552 nsew signal input
rlabel metal2 s 78337 995407 78393 995887 6 mprj_io_vtrip_sel[23]
port 553 nsew signal input
rlabel metal2 s 91217 995407 91273 995887 6 mprj_io_in[23]
port 554 nsew signal tristate
rlabel metal2 s 41713 966733 42193 966789 6 mprj_analog_io[17]
port 555 nsew signal bidirectional
rlabel metal5 s 6598 956420 19088 968960 6 mprj_io[24]
port 556 nsew signal bidirectional
rlabel metal2 s 41713 964341 42193 964397 6 mprj_io_analog_en[24]
port 557 nsew signal input
rlabel metal2 s 41713 963053 42193 963109 6 mprj_io_analog_pol[24]
port 558 nsew signal input
rlabel metal2 s 41713 960017 42193 960073 6 mprj_io_analog_sel[24]
port 559 nsew signal input
rlabel metal2 s 41713 963697 42193 963753 6 mprj_io_dm[72]
port 560 nsew signal input
rlabel metal2 s 41713 965537 42193 965593 6 mprj_io_dm[73]
port 561 nsew signal input
rlabel metal2 s 41713 959373 42193 959429 6 mprj_io_dm[74]
port 562 nsew signal input
rlabel metal2 s 41713 958729 42193 958785 6 mprj_io_holdover[24]
port 563 nsew signal input
rlabel metal2 s 41713 955693 42193 955749 6 mprj_io_ib_mode_sel[24]
port 564 nsew signal input
rlabel metal2 s 41713 962501 42193 962557 6 mprj_io_inp_dis[24]
port 565 nsew signal input
rlabel metal2 s 41713 955049 42193 955105 6 mprj_io_oeb[24]
port 566 nsew signal input
rlabel metal2 s 41713 958177 42193 958233 6 mprj_io_out[24]
port 567 nsew signal input
rlabel metal2 s 41713 967377 42193 967433 6 mprj_io_slow_sel[24]
port 568 nsew signal input
rlabel metal2 s 41713 956337 42193 956393 6 mprj_io_vtrip_sel[24]
port 569 nsew signal input
rlabel metal2 s 41713 969217 42193 969273 6 mprj_io_in[24]
port 570 nsew signal tristate
rlabel metal2 s 41713 796933 42193 796989 6 mprj_analog_io[18]
port 571 nsew signal bidirectional
rlabel metal5 s 6598 786620 19088 799160 6 mprj_io[25]
port 572 nsew signal bidirectional
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[25]
port 573 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[25]
port 574 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[25]
port 575 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[75]
port 576 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[76]
port 577 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[77]
port 578 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[25]
port 579 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[25]
port 580 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[25]
port 581 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[25]
port 582 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[25]
port 583 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[25]
port 584 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[25]
port 585 nsew signal input
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[25]
port 586 nsew signal tristate
rlabel metal2 s 41713 753733 42193 753789 6 mprj_analog_io[19]
port 587 nsew signal bidirectional
rlabel metal5 s 6598 743420 19088 755960 6 mprj_io[26]
port 588 nsew signal bidirectional
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[26]
port 589 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[26]
port 590 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[26]
port 591 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[78]
port 592 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[79]
port 593 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[80]
port 594 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[26]
port 595 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[26]
port 596 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[26]
port 597 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[26]
port 598 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[26]
port 599 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[26]
port 600 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[26]
port 601 nsew signal input
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[26]
port 602 nsew signal tristate
rlabel metal2 s 41713 710533 42193 710589 6 mprj_analog_io[20]
port 603 nsew signal bidirectional
rlabel metal5 s 6598 700220 19088 712760 6 mprj_io[27]
port 604 nsew signal bidirectional
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[27]
port 605 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[27]
port 606 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[27]
port 607 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[81]
port 608 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[82]
port 609 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[83]
port 610 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[27]
port 611 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[27]
port 612 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[27]
port 613 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[27]
port 614 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[27]
port 615 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[27]
port 616 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[27]
port 617 nsew signal input
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[27]
port 618 nsew signal tristate
rlabel metal2 s 41713 667333 42193 667389 6 mprj_analog_io[21]
port 619 nsew signal bidirectional
rlabel metal5 s 6598 657020 19088 669560 6 mprj_io[28]
port 620 nsew signal bidirectional
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[28]
port 621 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[28]
port 622 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[28]
port 623 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[84]
port 624 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[85]
port 625 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[86]
port 626 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[28]
port 627 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[28]
port 628 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[28]
port 629 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[28]
port 630 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[28]
port 631 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[28]
port 632 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[28]
port 633 nsew signal input
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[28]
port 634 nsew signal tristate
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 635 nsew signal input
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 636 nsew signal input
rlabel metal4 s 132600 36323 132792 37013 6 vdda
port 638 nsew signal bidirectional
rlabel metal4 s 132600 28653 147600 28719 6 vssa
port 639 nsew signal bidirectional
rlabel metal5 s 697980 909666 711432 920546 6 vccd1_pad
port 641 nsew signal bidirectional
rlabel metal5 s 698624 819822 710788 831990 6 vdda1_pad
port 642 nsew signal bidirectional
rlabel metal5 s 698624 505222 710788 517390 6 vdda1_pad2
port 643 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030788 6 vssa1_pad
port 644 nsew signal bidirectional
rlabel metal5 s 698624 417022 710788 429190 6 vssa1_pad2
port 645 nsew signal bidirectional
rlabel metal4 s 680587 459800 681277 459992 6 vdda1
port 647 nsew signal bidirectional
rlabel metal4 s 688881 459800 688947 474800 6 vssa1
port 648 nsew signal bidirectional
rlabel metal5 s 697980 461866 711432 472746 6 vssd1_pad
port 650 nsew signal bidirectional
rlabel metal5 s 6167 914054 19619 924934 6 vccd2_pad
port 651 nsew signal bidirectional
rlabel metal5 s 6811 484410 18975 496578 6 vdda2_pad
port 652 nsew signal bidirectional
rlabel metal5 s 6811 829010 18975 841178 6 vssa2_pad
port 653 nsew signal bidirectional
rlabel metal4 s 38503 455546 39593 455800 6 vccd
port 654 nsew signal bidirectional
rlabel metal4 s 36323 455607 37013 455799 6 vdda2
port 656 nsew signal bidirectional
rlabel metal4 s 32933 455546 33623 455800 6 vddio
port 657 nsew signal bidirectional
rlabel metal4 s 28653 440800 28719 455800 6 vssa2
port 658 nsew signal bidirectional
rlabel metal5 s 6167 442854 19619 453734 6 vssd2_pad
port 660 nsew signal bidirectional
rlabel metal4 s 7 455645 4843 456093 6 vssio
port 661 nsew signal bidirectional
flabel metal5 41130 179416 43498 180132 0 FreeSans 3200 0 0 0 vssd2
port 659 nsew
flabel metal5 44242 179326 46748 180098 0 FreeSans 3200 0 0 0 vccd2
port 655 nsew
flabel metal5 670926 95262 673290 96090 0 FreeSans 3200 180 0 0 vssd1
port 649 nsew
flabel metal5 674122 95266 676502 96062 0 FreeSans 3200 180 0 0 vccd1
port 646 nsew
rlabel metal4 s 132580 30762 132848 31674 6 vssd
port 640 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
