VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO xres_buf
  CLASS BLOCK ;
  FOREIGN xres_buf ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.000 BY 17.000 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.420 13.000 16.700 19.000 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 2.980 -2.000 3.260 4.000 ;
    END
  END X
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3.950 3.815 4.850 16.535 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 10.450 3.815 11.350 16.535 ;
    END
  END VGND
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.350 4.070 9.250 16.280 ;
    END
  END LVPWR
  PIN LVGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.850 4.070 15.750 16.280 ;
    END
  END LVGND
  OBS
      LAYER nwell ;
        RECT 2.070 10.025 10.170 14.395 ;
        RECT 2.070 3.655 17.610 6.255 ;
      LAYER li1 ;
        RECT 2.400 3.985 17.280 16.365 ;
      LAYER met1 ;
        RECT 2.400 3.815 17.280 16.535 ;
      LAYER met2 ;
        RECT 2.990 12.720 16.140 16.535 ;
        RECT 2.990 4.280 16.630 12.720 ;
        RECT 3.540 3.815 16.630 4.280 ;
      LAYER met3 ;
        RECT 3.950 3.905 11.350 16.445 ;
  END
END xres_buf
END LIBRARY

