module open_source ();
endmodule
