magic
tech sky130A
magscale 1 2
timestamp 1695745122
<< metal1 >>
rect 675768 115799 675774 116011
rect 675826 115799 675832 116011
rect 675682 113371 675734 115709
rect 675586 112665 675638 112671
rect 675586 112487 675638 112493
rect 675588 108330 675636 112487
rect 675682 108990 675734 113199
rect 675586 108324 675638 108330
rect 675586 108146 675638 108152
rect 675588 100462 675636 108146
rect 675586 100456 675638 100462
rect 675586 100278 675638 100284
rect 675588 100265 675636 100278
rect 675682 99896 675734 108806
rect 675776 102383 675824 115799
rect 675878 109636 675930 109642
rect 675878 109452 675930 109458
rect 675774 102377 675826 102383
rect 675774 102119 675826 102125
rect 675880 101831 675928 109452
rect 677392 103462 677399 103674
rect 677451 103514 677458 103674
rect 677451 103462 677652 103514
rect 675878 101825 675930 101831
rect 675878 101567 675930 101573
<< via1 >>
rect 675774 115799 675826 116011
rect 675682 113199 675734 113371
rect 675586 112493 675638 112665
rect 675682 108806 675734 108990
rect 675586 108152 675638 108324
rect 675586 100284 675638 100456
rect 675878 109458 675930 109636
rect 675774 102125 675826 102377
rect 677399 103462 677451 103674
rect 675878 101573 675930 101825
<< metal2 >>
rect 675774 116011 675826 116017
rect 676698 116015 676758 116024
rect 675826 115961 676698 116009
rect 675826 115801 675836 115961
rect 676685 115801 676698 115961
rect 675774 115793 675826 115799
rect 676698 115786 676758 115795
rect 677000 115915 677278 115920
rect 677000 115801 677159 115915
rect 677273 115801 677282 115915
rect 677000 115796 677278 115801
rect 677000 115703 677085 115796
rect 675831 115647 677085 115703
rect 677025 115279 677614 115325
rect 677025 115151 677071 115279
rect 675874 115095 677071 115151
rect 676855 114870 677614 114916
rect 676855 114507 676901 114870
rect 675874 114451 676901 114507
rect 677017 114722 677614 114774
rect 677017 113863 677069 114722
rect 675874 113807 677069 113863
rect 676969 113397 677614 113449
rect 675676 113199 675682 113371
rect 675734 113311 675740 113371
rect 676969 113311 677021 113397
rect 675734 113255 677021 113311
rect 675734 113199 675740 113255
rect 677022 112686 677614 112738
rect 677022 112667 677074 112686
rect 675580 112665 677074 112667
rect 675580 112493 675586 112665
rect 675638 112611 677074 112665
rect 675638 112493 675644 112611
rect 675874 111967 677216 112023
rect 677164 111529 677216 111967
rect 677164 111477 677614 111529
rect 675874 111415 677044 111471
rect 675874 110771 676892 110827
rect 676836 110302 676892 110771
rect 676992 110680 677044 111415
rect 676992 110628 677614 110680
rect 676836 110250 677614 110302
rect 675874 110127 676727 110183
rect 676671 109850 676727 110127
rect 676671 109798 677614 109850
rect 675872 109637 675936 109643
rect 675872 109636 677614 109637
rect 675872 109458 675878 109636
rect 675930 109585 677614 109636
rect 675930 109581 676776 109585
rect 675930 109458 675936 109581
rect 675872 109451 675936 109458
rect 675676 108990 675740 108997
rect 675676 108806 675682 108990
rect 675734 108908 675740 108990
rect 675734 108856 677614 108908
rect 675734 108806 675740 108856
rect 675676 108799 675740 108806
rect 675580 108326 675644 108331
rect 675580 108324 677230 108326
rect 675580 108152 675586 108324
rect 675638 108322 677230 108324
rect 675638 108270 677614 108322
rect 675638 108152 675644 108270
rect 675580 108145 675644 108152
rect 675874 107643 677216 107699
rect 675874 107091 677086 107147
rect 677020 106982 677086 107091
rect 677016 106766 677025 106982
rect 677081 106766 677090 106982
rect 677164 106951 677216 107643
rect 677164 106899 677614 106951
rect 677020 106761 677086 106766
rect 675874 106447 677230 106503
rect 677174 106029 677230 106447
rect 677174 105977 677614 106029
rect 675874 105803 677451 105859
rect 676806 105386 677010 105390
rect 675407 105381 677015 105386
rect 675407 105172 676806 105381
rect 676801 104977 676806 105172
rect 677010 104977 677015 105381
rect 676801 104972 677015 104977
rect 676806 104968 677010 104972
rect 675874 104607 676520 104663
rect 675407 103375 676368 103503
rect 676240 103038 676368 103375
rect 676466 103185 676518 104607
rect 677399 103674 677451 105803
rect 677399 103456 677451 103462
rect 676466 103133 677240 103185
rect 676240 102910 677133 103038
rect 675874 102767 676909 102823
rect 675769 102377 675832 102383
rect 675769 102125 675774 102377
rect 675826 102179 675832 102377
rect 675826 102125 676776 102179
rect 675769 102123 676776 102125
rect 675769 102116 675832 102123
rect 675871 101825 675936 101834
rect 675871 101573 675878 101825
rect 675930 101627 675936 101825
rect 675930 101573 676610 101627
rect 675871 101571 676610 101573
rect 675871 101564 675936 101571
rect 675874 100927 676467 100983
rect 675580 100456 675644 100463
rect 675580 100284 675586 100456
rect 675638 100339 675644 100456
rect 675638 100284 676255 100339
rect 676401 100307 676467 100927
rect 675580 100283 676255 100284
rect 675580 100276 675644 100283
rect 676214 100057 676254 100283
rect 676397 100091 676406 100307
rect 676462 100091 676471 100307
rect 676570 100259 676610 101571
rect 676710 100595 676776 102123
rect 676710 100379 676715 100595
rect 676771 100379 676776 100595
rect 676857 100478 676909 102767
rect 677005 100744 677133 102910
rect 677188 102633 677240 103133
rect 677188 102581 677614 102633
rect 677005 100616 677614 100744
rect 676857 100426 677614 100478
rect 676710 100374 676776 100379
rect 676715 100370 676771 100374
rect 676570 100219 677614 100259
rect 676401 100086 676467 100091
rect 676214 100017 677614 100057
<< via2 >>
rect 676698 115795 676758 116015
rect 677159 115801 677273 115915
rect 677025 106766 677081 106982
rect 676806 104977 677010 105381
rect 676406 100091 676462 100307
rect 676715 100379 676771 100595
<< metal3 >>
rect 676696 116020 676756 117658
rect 676693 116015 676763 116020
rect 676693 115795 676698 116015
rect 676758 115795 676763 116015
rect 677154 115915 677614 115920
rect 677154 115801 677159 115915
rect 677273 115801 677614 115915
rect 677154 115796 677614 115801
rect 676693 115790 676763 115795
rect 676696 115783 676756 115790
rect 677020 106982 677095 106987
rect 677020 106766 677025 106982
rect 677081 106827 677095 106982
rect 677081 106766 677614 106827
rect 677020 106761 677614 106766
rect 676801 105381 677015 105386
rect 676801 104977 676806 105381
rect 677010 104977 677015 105381
rect 676801 103436 677015 104977
rect 676801 103222 677614 103436
rect 676710 100595 676776 100600
rect 676710 100379 676715 100595
rect 676771 100379 676776 100595
rect 676401 100307 676472 100312
rect 676401 100091 676406 100307
rect 676462 100152 676472 100307
rect 676710 100284 676776 100379
rect 676710 100218 677614 100284
rect 676462 100091 677614 100152
rect 676401 100086 677614 100091
<< properties >>
string flatten true
<< end >>
