magic
tech sky130A
magscale 1 2
timestamp 1513420866
<< checkpaint >>
rect -4476 -9457 636864 957006
<< metal3 >>
tri 39202 941418 39844 942060 se
rect 39844 941960 44844 955662
rect 39844 941418 44302 941960
tri 44302 941418 44844 941960 nw
rect 91244 941418 96244 955672
rect 39202 940618 44202 941418
tri 44202 941318 44302 941418 nw
rect 91202 941282 96244 941418
rect 142644 941418 147644 955636
rect 178700 953492 192979 955636
rect 178700 951748 179127 953492
rect 192551 951748 192979 953492
rect 178700 951320 192979 951748
tri 178700 942060 187960 951320 ne
rect 187960 942060 192979 951320
tri 187960 941960 188060 942060 ne
rect 188060 941960 192979 942060
tri 188060 941418 188602 941960 ne
rect 188602 941418 192979 941960
rect 193279 942041 195479 955636
rect 195678 942142 197878 955636
tri 195678 942041 195779 942142 ne
rect 195779 942041 197878 942142
tri 193279 941418 193902 942041 ne
rect 193902 941418 195479 942041
tri 195779 941768 196052 942041 ne
rect 196052 941768 197878 942041
rect 198178 953492 212500 955636
rect 198178 951748 198605 953492
rect 212029 951748 212500 953492
rect 198178 950016 212500 951748
rect 231300 953492 245579 955654
rect 231300 951748 231727 953492
rect 245151 951748 245579 953492
rect 231300 950420 245579 951748
tri 231300 950016 231704 950420 ne
rect 231704 950016 245579 950420
rect 198178 942142 204626 950016
tri 204626 942142 212500 950016 nw
tri 231704 942142 239578 950016 ne
rect 239578 942142 245579 950016
tri 198178 941768 198552 942142 ne
rect 198552 941768 204252 942142
tri 204252 941768 204626 942142 nw
tri 239578 941768 239952 942142 ne
rect 239952 941768 245579 942142
tri 195479 941418 195829 941768 sw
tri 196052 941418 196402 941768 ne
rect 196402 941418 197878 941768
tri 197878 941418 198228 941768 sw
tri 198552 941418 198902 941768 ne
rect 142644 941352 148202 941418
rect 91202 940618 96202 941282
rect 143202 940618 148202 941352
rect 188602 940618 193602 941418
rect 193902 940618 196102 941418
rect 196402 940618 198602 941418
rect 198902 940618 203902 941768
tri 203902 941418 204252 941768 nw
tri 239952 941418 240302 941768 ne
rect 240302 941695 245579 941768
rect 240302 940618 245302 941695
tri 245302 941418 245579 941695 nw
rect 245879 941695 248079 955654
rect 245879 941618 248002 941695
tri 248002 941618 248079 941695 nw
tri 245679 941418 245879 941618 se
rect 245879 941418 247802 941618
tri 247802 941418 248002 941618 nw
rect 248278 941594 250478 955654
tri 248102 941418 248278 941594 se
rect 248278 941418 250302 941594
tri 250302 941418 250478 941594 nw
rect 250778 953492 265100 955654
rect 250778 951748 251205 953492
rect 264629 951748 265100 953492
rect 250778 950916 265100 951748
rect 250778 950420 264604 950916
tri 264604 950420 265100 950916 nw
rect 333100 953492 347379 955622
rect 333100 951748 333527 953492
rect 346951 951748 347379 953492
rect 250778 941695 255879 950420
tri 255879 941695 264604 950420 nw
rect 333100 950320 347379 951748
tri 333100 941695 341725 950320 ne
rect 341725 941795 347379 950320
rect 341725 941695 347002 941795
rect 250778 941618 255802 941695
tri 255802 941618 255879 941695 nw
tri 341725 941618 341802 941695 ne
rect 341802 941618 347002 941695
rect 250778 941594 255778 941618
tri 255778 941594 255802 941618 nw
tri 341802 941594 341826 941618 ne
rect 341826 941594 347002 941618
rect 250778 941418 255602 941594
tri 255602 941418 255778 941594 nw
tri 341826 941418 342002 941594 ne
rect 245602 940618 247802 941418
rect 248102 940618 250302 941418
rect 250602 940618 255602 941418
rect 342002 940618 347002 941594
tri 347002 941418 347379 941795 nw
rect 347679 941795 349879 955622
rect 347679 941698 349782 941795
tri 349782 941698 349879 941795 nw
tri 347399 941418 347679 941698 se
rect 347679 941694 349778 941698
tri 349778 941694 349782 941698 nw
rect 350078 941694 352278 955622
rect 347679 941418 349502 941694
tri 349502 941418 349778 941694 nw
tri 349802 941418 350078 941694 se
rect 350078 941418 352002 941694
tri 352002 941418 352278 941694 nw
rect 352578 953492 366900 955622
rect 352578 951748 353005 953492
rect 366429 951748 366900 953492
rect 352578 951016 366900 951748
rect 352578 950916 366800 951016
tri 366800 950916 366900 951016 nw
rect 352578 950420 366304 950916
tri 366304 950420 366800 950916 nw
rect 352578 950320 366204 950420
tri 366204 950320 366304 950420 nw
rect 352578 941795 357679 950320
tri 357679 941795 366204 950320 nw
rect 352578 941698 357582 941795
tri 357582 941698 357679 941795 nw
rect 352578 941694 357578 941698
tri 357578 941694 357582 941698 nw
rect 352578 941418 357302 941694
tri 357302 941418 357578 941694 nw
rect 436444 941418 441444 955604
rect 487844 941964 492844 955692
rect 533400 946135 538179 955592
rect 533400 942391 533585 946135
rect 537969 942391 538179 946135
tri 492844 941964 492856 941976 sw
tri 487844 941795 488013 941964 ne
rect 488013 941795 492856 941964
tri 488013 941698 488110 941795 ne
rect 488110 941698 492856 941795
tri 488110 941694 488114 941698 ne
rect 488114 941694 492856 941698
tri 488114 941418 488390 941694 ne
rect 488390 941418 492856 941694
tri 492856 941418 493402 941964 sw
rect 533400 941578 538179 942391
rect 543378 946135 548158 955592
rect 543378 942391 543585 946135
rect 547969 942391 548158 946135
rect 543378 941641 548158 942391
tri 548158 941641 548179 941662 sw
tri 538179 941578 538242 941641 sw
rect 543378 941600 548179 941641
tri 548179 941600 548220 941641 sw
tri 543378 941578 543400 941600 ne
rect 543400 941578 548220 941600
tri 533400 941418 533560 941578 ne
rect 533560 941418 538242 941578
tri 538242 941418 538402 941578 sw
tri 543400 941418 543560 941578 ne
rect 543560 941418 548220 941578
tri 548220 941418 548402 941600 sw
rect 589644 941418 594644 955746
rect 347302 940618 349502 941418
rect 349802 940618 352002 941418
rect 352302 940618 357302 941418
rect 436402 941284 441444 941418
tri 488390 941406 488402 941418 ne
rect 436402 940618 441402 941284
rect 488402 940618 493402 941418
tri 533560 941406 533572 941418 ne
rect 533572 941406 538402 941418
tri 533572 941376 533602 941406 ne
rect 533602 940618 538402 941406
tri 543560 941376 543602 941418 ne
rect 543602 940618 548402 941418
rect 589602 941274 594644 941418
rect 589602 940618 594602 941274
rect -2536 921860 21164 923044
tri 21164 921860 22348 923044 sw
rect -2536 918044 23008 921860
tri 21025 916861 22208 918044 ne
rect 22208 916860 23008 918044
rect 607008 919556 607808 919602
rect 607008 914602 635506 919556
rect 607716 914556 635506 914602
rect 22208 884840 23008 885260
rect -3216 884758 23008 884840
rect -3216 880134 -1777 884758
rect 1087 880460 23008 884758
rect 1087 880134 22252 880460
rect -3216 880051 22252 880134
rect 607008 880402 607808 881202
tri 607808 880402 608608 881202 sw
rect 607008 880400 634180 880402
rect 607008 880318 635604 880400
rect -2200 879648 1182 879730
rect -2200 875184 -1777 879648
rect 1087 875184 1182 879648
rect 607008 876402 631301 880318
tri 607626 875600 608428 876402 ne
rect 608428 875694 631301 876402
rect 634165 875694 635604 880318
rect 608428 875611 635604 875694
rect 608428 875600 634180 875611
rect -2200 875120 1182 875184
rect 22208 874800 23008 875261
rect -3216 874718 23008 874800
rect -3216 870094 -1777 874718
rect 1087 870460 23008 874718
rect 631206 875208 635204 875290
rect 1087 870094 22260 870460
rect -3216 870011 22260 870094
rect -1244 870000 22260 870011
rect 607008 870349 607808 871202
tri 607808 870349 608661 871202 sw
rect 631206 870744 631301 875208
rect 634165 870744 635204 875208
rect 631206 870669 635204 870744
rect 607008 870267 635604 870349
rect 607008 866402 631301 870267
tri 607634 865560 608476 866402 ne
rect 608476 865643 631301 866402
rect 634165 865643 635604 870267
rect 608476 865560 635604 865643
tri 21706 800358 22208 800860 se
rect 22208 800358 23008 800860
rect -2400 800174 23008 800358
rect -2400 795790 17500 800174
rect 21244 796060 23008 800174
rect 21244 795790 21852 796060
rect -2400 795578 21852 795790
tri 21852 795578 22334 796060 nw
rect 607008 791201 607808 791980
rect 607008 791015 635332 791201
tri 21727 790379 22208 790860 se
rect 22208 790379 23008 790860
rect -2400 790174 23008 790379
rect -2400 786060 17500 790174
rect 7592 786059 17500 786060
rect -2400 785790 17500 786059
rect 21244 786060 23008 790174
rect 607008 787180 613569 791015
rect 607558 786631 613569 787180
rect 617313 786631 635332 791015
rect 607558 786421 635332 786631
rect 21244 786059 22334 786060
rect 21244 785790 21874 786059
rect -2400 785599 21874 785790
tri 21874 785599 22334 786059 nw
rect 607008 781222 607808 781980
rect 607008 781015 635332 781222
rect 607008 777180 613569 781015
rect 607558 776631 613569 777180
rect 617313 776631 635332 781015
rect 607558 776442 635332 776631
rect 607008 476601 607808 476648
rect 607008 476415 635332 476601
rect 607008 472031 613569 476415
rect 617313 472031 635332 476415
rect 607008 471848 635332 472031
rect 607758 471821 624816 471848
rect 607008 466622 607808 466648
rect 607008 466415 635332 466622
rect 607008 462031 613569 466415
rect 617313 462031 635332 466415
rect 607008 461848 635332 462031
rect 607766 461842 624824 461848
tri 21660 455758 22208 456306 se
rect 22208 455758 23008 456306
rect -2400 455574 23008 455758
rect -2400 451190 13000 455574
rect 16744 451506 23008 455574
rect 16744 451190 21712 451506
rect -2400 450978 21712 451190
tri 21712 450978 22240 451506 nw
tri 21682 445779 22208 446305 se
rect 22208 445779 23008 446306
rect -2400 445574 23008 445779
rect -2400 441190 13000 445574
rect 16744 441506 23008 445574
rect 16744 441190 21741 441506
rect -2400 440999 21741 441190
tri 21741 440999 22248 441506 nw
rect 607008 432600 607808 432848
rect 607008 432518 635604 432600
rect 607008 428048 631301 432518
rect 607742 427894 631301 428048
rect 634165 427894 635604 432518
rect 607742 427811 635604 427894
rect 607742 427800 633878 427811
rect 631206 427408 635204 427490
rect 631206 422944 631301 427408
rect 634165 422944 635204 427408
rect 631206 422869 635204 422944
rect 607008 422549 607808 422848
rect 607008 422467 635604 422549
rect 607008 418048 631301 422467
rect 607742 417843 631301 418048
rect 634165 417843 635604 422467
rect 607742 417760 635604 417843
tri 21542 413640 22208 414306 se
rect 22208 413640 23008 414306
rect -3216 413558 23008 413640
rect -3216 408934 -1777 413558
rect 1087 409506 23008 413558
rect 1087 408934 21627 409506
rect -3216 408851 21627 408934
tri 21627 408851 22282 409506 nw
rect -2216 408448 1182 408530
rect -2216 403984 -1777 408448
rect 1087 403984 1182 408448
rect -2216 403920 1182 403984
tri 21822 403920 22208 404306 se
rect 22208 403920 23008 404306
tri 21502 403600 21822 403920 se
rect 21822 403600 23008 403920
rect -3216 403518 23008 403600
rect -3216 398894 -1777 403518
rect 1087 399506 23008 403518
rect 1087 398894 21558 399506
rect -3216 398811 21558 398894
rect -900 398800 21558 398811
tri 21558 398800 22264 399506 nw
rect 607768 388248 635376 388401
rect 607008 388215 635376 388248
rect 607008 383831 608769 388215
rect 612513 383831 635376 388215
rect 607008 383621 635376 383831
rect 607008 383462 634724 383621
rect 607008 383448 607808 383462
rect 607758 378248 635376 378422
rect 607008 378215 635376 378248
rect 607008 373831 608769 378215
rect 612513 373831 635376 378215
rect 607008 373642 635376 373831
rect 607008 373448 607808 373642
rect -3216 40758 1182 40840
rect -3216 36134 -1777 40758
rect 1087 36134 1182 40758
rect -3216 36051 1182 36134
rect -3216 30718 1182 30800
rect -3216 26094 -1777 30718
rect 1087 26094 1182 30718
rect 208144 27328 212703 27373
rect 208144 27104 208191 27328
rect 209055 27104 212703 27328
rect 208144 27054 212703 27104
rect 226824 26900 227464 26936
rect 223584 26888 227464 26900
rect 223584 26664 226871 26888
rect 227415 26664 227464 26888
rect 223584 26653 227464 26664
rect 226824 26619 227464 26653
rect -3216 26011 1182 26094
rect 130944 7832 139976 7881
rect 130944 7608 130995 7832
rect 131859 7733 139976 7832
rect 131859 7608 139772 7733
rect 130944 7589 139772 7608
rect 139916 7589 139976 7733
rect 130944 7560 139976 7589
rect 132304 7169 138678 7214
rect 132304 7168 138472 7169
rect 132304 6944 132347 7168
rect 133211 7025 138472 7168
rect 138616 7025 138678 7169
rect 133211 6944 138678 7025
rect 132304 6894 138678 6944
rect 198943 -112 203749 -22
rect 171700 -225 175302 -135
rect 171700 -1809 171798 -225
rect 175222 -1809 175302 -225
rect 171700 -6251 175302 -1809
rect 193205 -225 195949 -135
rect 193205 -1809 193303 -225
rect 195847 -1809 195949 -225
rect 193205 -7342 195949 -1809
rect 198943 -1696 199023 -112
rect 203647 -1696 203749 -112
rect 198943 -2938 203749 -1696
rect 208994 -112 213800 -22
rect 208994 -1696 209074 -112
rect 213698 -1696 213800 -112
rect 208994 -2938 213800 -1696
rect 193205 -8126 193308 -7342
rect 195772 -8126 195949 -7342
rect 193205 -8197 195949 -8126
<< via3 >>
rect 179127 951748 192551 953492
rect 198605 951748 212029 953492
rect 231727 951748 245151 953492
rect 251205 951748 264629 953492
rect 333527 951748 346951 953492
rect 353005 951748 366429 953492
rect 533585 942391 537969 946135
rect 543585 942391 547969 946135
rect -1777 880134 1087 884758
rect -1777 875184 1087 879648
rect 631301 875694 634165 880318
rect -1777 870094 1087 874718
rect 631301 870744 634165 875208
rect 631301 865643 634165 870267
rect 17500 795790 21244 800174
rect 17500 785790 21244 790174
rect 613569 786631 617313 791015
rect 613569 776631 617313 781015
rect 613569 472031 617313 476415
rect 613569 462031 617313 466415
rect 13000 451190 16744 455574
rect 13000 441190 16744 445574
rect 631301 427894 634165 432518
rect 631301 422944 634165 427408
rect 631301 417843 634165 422467
rect -1777 408934 1087 413558
rect -1777 403984 1087 408448
rect -1777 398894 1087 403518
rect 608769 383831 612513 388215
rect 608769 373831 612513 378215
rect -1777 36134 1087 40758
rect -1777 26094 1087 30718
rect 208191 27104 209055 27328
rect 226871 26664 227415 26888
rect 130995 7608 131859 7832
rect 139772 7589 139916 7733
rect 132347 6944 133211 7168
rect 138472 7025 138616 7169
rect 171798 -1809 175222 -225
rect 193303 -1809 195847 -225
rect 199023 -1696 203647 -112
rect 209074 -1696 213698 -112
rect 193308 -8126 195772 -7342
<< metal4 >>
rect 178700 953492 192979 953920
rect 178700 951748 179127 953492
rect 192551 951748 192979 953492
rect 178700 951320 192979 951748
tri 178700 946135 183885 951320 ne
rect 183885 946135 192979 951320
tri 183885 942391 187629 946135 ne
rect 187629 942391 192979 946135
tri 187629 941418 188602 942391 ne
rect 188602 941418 192979 942391
rect 198178 953492 212457 953920
rect 198178 951748 198605 953492
rect 212029 951748 212457 953492
rect 198178 951720 212457 951748
rect 231300 953492 245579 953920
rect 231300 951748 231727 953492
rect 245151 951748 245579 953492
rect 198178 950016 212500 951720
rect 231300 950420 245579 951748
tri 231300 950016 231704 950420 ne
rect 231704 950016 245579 950420
rect 198178 946135 208619 950016
tri 208619 946135 212500 950016 nw
tri 231704 946135 235585 950016 ne
rect 235585 946135 245579 950016
rect 198178 942391 204875 946135
tri 204875 942391 208619 946135 nw
tri 235585 942391 239329 946135 ne
rect 239329 942391 245579 946135
rect 198178 942142 204626 942391
tri 204626 942142 204875 942391 nw
tri 239329 942142 239578 942391 ne
rect 239578 942142 245579 942391
tri 198178 941418 198902 942142 ne
rect 188602 940618 193602 941418
rect 198902 940618 203902 942142
tri 203902 941418 204626 942142 nw
tri 239578 941418 240302 942142 ne
rect 240302 941695 245579 942142
rect 240302 940618 245302 941695
tri 245302 941418 245579 941695 nw
rect 250778 953492 265057 953920
rect 250778 951748 251205 953492
rect 264629 951748 265057 953492
rect 250778 951720 265057 951748
rect 333100 953492 347379 953920
rect 333100 951748 333527 953492
rect 346951 951748 347379 953492
rect 250778 950916 265100 951720
rect 250778 950420 264604 950916
tri 264604 950420 265100 950916 nw
rect 250778 946135 260319 950420
tri 260319 946135 264604 950420 nw
rect 333100 950320 347379 951748
tri 333100 946135 337285 950320 ne
rect 337285 946135 347379 950320
rect 250778 942391 256575 946135
tri 256575 942391 260319 946135 nw
tri 337285 942391 341029 946135 ne
rect 341029 942391 347379 946135
rect 250778 941695 255879 942391
tri 255879 941695 256575 942391 nw
tri 341029 941695 341725 942391 ne
rect 341725 941795 347379 942391
rect 341725 941695 347002 941795
rect 250778 941418 255602 941695
tri 255602 941418 255879 941695 nw
tri 341725 941418 342002 941695 ne
rect 250602 940618 255602 941418
rect 342002 940618 347002 941695
tri 347002 941418 347379 941795 nw
rect 352578 953492 366857 953920
rect 352578 951748 353005 953492
rect 366429 951748 366857 953492
rect 352578 951720 366857 951748
rect 352578 951016 366900 951720
rect 352578 950916 366800 951016
tri 366800 950916 366900 951016 nw
rect 352578 950420 366304 950916
tri 366304 950420 366800 950916 nw
rect 352578 950320 366204 950420
tri 366204 950320 366304 950420 nw
rect 352578 946135 362019 950320
tri 362019 946135 366204 950320 nw
rect 533401 946135 538179 946282
rect 352578 942391 358275 946135
tri 358275 942391 362019 946135 nw
rect 533401 942391 533585 946135
rect 537969 942391 538179 946135
rect 352578 941795 357679 942391
tri 357679 941795 358275 942391 nw
rect 533401 942282 538179 942391
rect 543378 946135 548158 946282
rect 543378 942391 543585 946135
rect 547969 942391 548158 946135
rect 543378 942282 548158 942391
rect 352578 941418 357302 941795
tri 357302 941418 357679 941795 nw
rect 352302 940618 357302 941418
rect -1858 884758 1182 884840
rect -1858 880134 -1777 884758
rect 1087 880134 1182 884758
rect -1858 880051 1182 880134
rect -1858 879648 1182 879730
rect -1858 875184 -1777 879648
rect 1087 875184 1182 879648
rect -1858 875120 1182 875184
rect 6984 879608 7984 884840
rect 6984 875212 7046 879608
rect 7922 875212 7984 879608
rect -1858 874718 1182 874800
rect -1858 870094 -1777 874718
rect 1087 870094 1182 874718
rect -1858 870011 1182 870094
rect 6984 808000 7984 875212
rect 8184 884718 9184 884840
rect 8184 880322 8246 884718
rect 9122 880322 9184 884718
rect 8184 874678 9184 880322
rect 8184 870282 8246 874678
rect 9122 870282 9184 874678
rect 8184 808000 9184 870282
rect 625836 875168 626836 880402
rect 625836 870772 625898 875168
rect 626774 870772 626836 875168
rect 17391 800174 21391 800358
rect 17391 795790 17500 800174
rect 21244 795790 21391 800174
rect 17391 795580 21391 795790
rect 613460 791015 617460 791199
rect 17391 790174 21391 790381
rect 17391 785790 17500 790174
rect 21244 785790 21391 790174
rect 613460 786631 613569 791015
rect 617313 786631 617460 791015
rect 625836 788000 626836 870772
rect 627036 880278 628036 880402
rect 627036 875882 627098 880278
rect 627974 875882 628036 880278
rect 627036 870227 628036 875882
rect 631206 880318 634246 880400
rect 631206 875694 631301 880318
rect 634165 875694 634246 880318
rect 631206 875611 634246 875694
rect 631206 875208 634246 875290
rect 631206 870744 631301 875208
rect 634165 870744 634246 875208
rect 631206 870669 634246 870744
rect 627036 865831 627098 870227
rect 627974 865831 628036 870227
rect 627036 788000 628036 865831
rect 631206 870267 634246 870349
rect 631206 865643 631301 870267
rect 634165 865643 634246 870267
rect 631206 865560 634246 865643
rect 613460 786421 617460 786631
rect 17391 785601 21391 785790
rect 613460 781015 617460 781222
rect 613460 776631 613569 781015
rect 617313 776631 617460 781015
rect 613460 776442 617460 776631
rect 613460 476415 617460 476599
rect 613460 472031 613569 476415
rect 617313 472031 617460 476415
rect 613460 471821 617460 472031
rect 613460 466415 617460 466622
rect 613460 462031 613569 466415
rect 617313 462031 617460 466415
rect 613460 461842 617460 462031
rect 12891 455574 16891 455758
rect 12891 451190 13000 455574
rect 16744 451190 16891 455574
rect 12891 450980 16891 451190
rect 12891 445574 16891 445781
rect 12891 441190 13000 445574
rect 16744 441190 16891 445574
rect 12891 441001 16891 441190
rect 631206 432518 634246 432600
rect 631206 427894 631301 432518
rect 634165 427894 634246 432518
rect 631206 427811 634246 427894
rect 631206 427408 634246 427490
rect 631206 422944 631301 427408
rect 634165 422944 634246 427408
rect 631206 422869 634246 422944
rect 631206 422467 634246 422549
rect 631206 417843 631301 422467
rect 634165 417843 634246 422467
rect 631206 417760 634246 417843
rect -1858 413558 1182 413640
rect -1858 408934 -1777 413558
rect 1087 408934 1182 413558
rect -1858 408851 1182 408934
rect -1858 408448 1182 408530
rect -1858 403984 -1777 408448
rect 1087 403984 1182 408448
rect -1858 403920 1182 403984
rect -1858 403518 1182 403600
rect -1858 398894 -1777 403518
rect 1087 398894 1182 403518
rect -1858 398811 1182 398894
rect 608660 388215 612660 388399
rect 608660 383831 608769 388215
rect 612513 383831 612660 388215
rect 608660 383462 612660 383831
rect 608660 378215 612660 378422
rect 608660 373831 608769 378215
rect 612513 373831 612660 378215
rect 608660 373642 612660 373831
rect 12891 243281 16891 243658
rect 12891 239205 13130 243281
rect 16566 239205 16891 243281
rect 12891 230754 16891 239205
rect 12891 228918 13130 230754
rect 16566 228918 16891 230754
rect 12891 228836 16891 228918
rect 608660 243281 612660 243658
rect 608660 239205 608899 243281
rect 612335 239205 612660 243281
rect 608660 228434 612660 239205
rect 608660 226598 608899 228434
rect 612335 226598 612660 228434
rect 608660 226516 612660 226598
rect 613460 243281 617460 243658
rect 613460 239205 613699 243281
rect 617135 239205 617460 243281
rect 613460 226114 617460 239205
rect 613460 224278 613699 226114
rect 617135 224278 617460 226114
rect 613460 224196 617460 224278
rect -1858 40758 1182 40840
rect -1858 36134 -1777 40758
rect 1087 36134 1182 40758
rect -1858 36051 1182 36134
rect 193205 34214 195949 34276
rect 193205 33338 193351 34214
rect 195827 33338 195949 34214
rect 171700 32814 175302 32876
rect 171700 31938 171946 32814
rect 175062 31938 175302 32814
rect -1858 30718 1182 30800
rect -1858 26094 -1777 30718
rect 1087 26094 1182 30718
rect 171700 30014 175302 31938
rect 171700 29138 171946 30014
rect 175062 29138 175302 30014
rect -1858 26011 1182 26094
rect 137400 6414 137791 6496
rect 137400 6178 137476 6414
rect 137712 6178 137791 6414
rect 137400 6094 137791 6178
rect 137400 5858 137476 6094
rect 137712 5858 137791 6094
rect 137400 5774 137791 5858
rect 137400 5538 137476 5774
rect 137712 5538 137791 5774
rect 137400 5454 137791 5538
rect 137400 5218 137476 5454
rect 137712 5218 137791 5454
rect 137400 5134 137791 5218
rect 137400 4898 137476 5134
rect 137712 4898 137791 5134
rect 137400 4814 137791 4898
rect 137400 4578 137476 4814
rect 137712 4578 137791 4814
rect 137400 4497 137791 4578
rect 138800 4094 139282 6496
rect 138800 3858 138932 4094
rect 139168 3858 139282 4094
rect 138800 3774 139282 3858
rect 138800 3538 138932 3774
rect 139168 3538 139282 3774
rect 138800 3454 139282 3538
rect 138800 3218 138932 3454
rect 139168 3218 139282 3454
rect 138800 3134 139282 3218
rect 138800 2898 138932 3134
rect 139168 2898 139282 3134
rect 138800 2814 139282 2898
rect 138800 2578 138932 2814
rect 139168 2578 139282 2814
rect 138800 2494 139282 2578
rect 138800 2258 138932 2494
rect 139168 2258 139282 2494
rect 138800 2176 139282 2258
rect 171700 -225 175302 29138
rect 171700 -1809 171798 -225
rect 175222 -1809 175302 -225
rect 171700 -1937 175302 -1809
rect 193205 31414 195949 33338
rect 193205 30538 193351 31414
rect 195827 30538 195949 31414
rect 193205 -225 195949 30538
rect 209504 27682 212862 28083
rect 223604 27047 226064 27376
rect 193205 -1809 193303 -225
rect 195847 -1809 195949 -225
rect 193205 -1937 195949 -1809
rect 198943 6414 203749 6496
rect 198943 4578 199106 6414
rect 203502 4578 203749 6414
rect 198943 -112 203749 4578
rect 198943 -1696 199023 -112
rect 203647 -1696 203749 -112
rect 198943 -1824 203749 -1696
rect 208994 6414 213800 6496
rect 208994 4578 209157 6414
rect 213553 4578 213800 6414
rect 208994 -112 213800 4578
rect 208994 -1696 209074 -112
rect 213698 -1696 213800 -112
rect 208994 -1824 213800 -1696
<< via4 >>
rect 179161 951862 192517 953378
rect 198639 951862 211995 953378
rect 231761 951862 245117 953378
rect 251239 951862 264595 953378
rect 333561 951862 346917 953378
rect 353039 951862 366395 953378
rect 533739 942465 537815 945901
rect 543739 942465 547815 945901
rect -1736 880322 1060 884718
rect -1736 875212 1060 879608
rect 7046 875212 7922 879608
rect -1736 870282 1060 874678
rect 8246 880322 9122 884718
rect 8246 870282 9122 874678
rect 625898 870772 626774 875168
rect 17574 795944 21010 800020
rect 17574 785944 21010 790020
rect 613643 786785 617079 790861
rect 627098 875882 627974 880278
rect 631328 875882 634124 880278
rect 631328 870772 634124 875168
rect 627098 865831 627974 870227
rect 631328 865831 634124 870227
rect 613643 776785 617079 780861
rect 613643 472185 617079 476261
rect 613643 462185 617079 466261
rect 13074 451344 16510 455420
rect 13074 441344 16510 445420
rect 625898 428082 626774 432478
rect 631328 428082 634124 432478
rect 627098 422972 627974 427368
rect 631328 422972 634124 427368
rect 625898 418031 626774 422427
rect 631328 418031 634124 422427
rect -1736 409122 1060 413518
rect 7046 409122 7922 413518
rect -1736 404012 1060 408408
rect 8246 404012 9122 408408
rect -1736 399082 1060 403478
rect 7046 399082 7922 403478
rect 608843 383985 612279 388061
rect 608843 373985 612279 378061
rect 13130 239205 16566 243281
rect 13130 228918 16566 230754
rect 608899 239205 612335 243281
rect 608899 226598 612335 228434
rect 613699 239205 617135 243281
rect 613699 224278 617135 226114
rect -1736 36322 1060 40718
rect 2246 36322 3122 40718
rect 193351 33338 195827 34214
rect 171946 31938 175062 32814
rect -1736 26282 1060 30678
rect 2246 26282 3122 30678
rect 171946 29138 175062 30014
rect 137476 6178 137712 6414
rect 137476 5858 137712 6094
rect 137476 5538 137712 5774
rect 137476 5218 137712 5454
rect 137476 4898 137712 5134
rect 137476 4578 137712 4814
rect 138932 3858 139168 4094
rect 138932 3538 139168 3774
rect 138932 3218 139168 3454
rect 138932 2898 139168 3134
rect 138932 2578 139168 2814
rect 138932 2258 139168 2494
rect 193351 30538 195827 31414
rect 199106 4578 203502 6414
rect 209157 4578 213553 6414
<< metal5 >>
rect 178700 953378 192979 953920
rect 178700 951862 179161 953378
rect 192517 951862 192979 953378
rect 178700 951320 192979 951862
tri 178700 941418 188602 951320 ne
rect 188602 941418 192979 951320
rect 198178 953378 212457 953920
rect 198178 951862 198639 953378
rect 211995 951862 212457 953378
rect 198178 951720 212457 951862
rect 231300 953378 245579 953920
rect 231300 951862 231761 953378
rect 245117 951862 245579 953378
rect 198178 950016 212500 951720
rect 231300 950420 245579 951862
tri 231300 950016 231704 950420 ne
rect 231704 950016 245579 950420
rect 198178 942142 204626 950016
tri 204626 942142 212500 950016 nw
tri 231704 942142 239578 950016 ne
rect 239578 942142 245579 950016
tri 198178 941418 198902 942142 ne
rect 188602 940618 193602 941418
rect 198902 940618 203902 942142
tri 203902 941418 204626 942142 nw
tri 239578 941418 240302 942142 ne
rect 240302 941695 245579 942142
rect 240302 940618 245302 941695
tri 245302 941418 245579 941695 nw
rect 250778 953378 265057 953920
rect 250778 951862 251239 953378
rect 264595 951862 265057 953378
rect 250778 951720 265057 951862
rect 333100 953378 347379 953920
rect 333100 951862 333561 953378
rect 346917 951862 347379 953378
rect 250778 950916 265100 951720
rect 250778 950420 264604 950916
tri 264604 950420 265100 950916 nw
rect 250778 941695 255879 950420
tri 255879 941695 264604 950420 nw
rect 333100 950320 347379 951862
tri 333100 941695 341725 950320 ne
rect 341725 941795 347379 950320
rect 341725 941695 347002 941795
rect 250778 941418 255602 941695
tri 255602 941418 255879 941695 nw
tri 341725 941418 342002 941695 ne
rect 250602 940618 255602 941418
rect 342002 940618 347002 941695
tri 347002 941418 347379 941795 nw
rect 352578 953378 366857 953920
rect 352578 951862 353039 953378
rect 366395 951862 366857 953378
rect 352578 951720 366857 951862
rect 352578 951016 366900 951720
rect 352578 950916 366800 951016
tri 366800 950916 366900 951016 nw
rect 352578 950420 366304 950916
tri 366304 950420 366800 950916 nw
rect 352578 950320 366204 950420
tri 366204 950320 366304 950420 nw
rect 352578 941795 357679 950320
tri 357679 941795 366204 950320 nw
rect 533400 945901 612660 946282
rect 533400 942465 533739 945901
rect 537815 942465 543739 945901
rect 547815 942465 612660 945901
rect 533400 942282 612660 942465
rect 352578 941418 357302 941795
tri 357302 941418 357679 941795 nw
rect 352302 940618 357302 941418
rect -1858 884718 9184 884840
rect -1858 880322 -1736 884718
rect 1060 880322 8246 884718
rect 9122 880322 9184 884718
rect -1858 880050 9184 880322
rect -1858 879608 7984 879730
rect -1858 875212 -1736 879608
rect 1060 875212 7046 879608
rect 7922 875212 7984 879608
rect -1858 875120 7984 875212
rect -1858 874678 9184 874800
rect -1858 870282 -1736 874678
rect 1060 870282 8246 874678
rect 9122 870282 9184 874678
rect -1858 870010 9184 870282
rect 17391 800020 21391 800358
rect 17391 795944 17574 800020
rect 21010 795944 21391 800020
rect 17391 790020 21391 795944
rect 17391 785944 17574 790020
rect 21010 785944 21391 790020
rect 12891 455420 16891 455758
rect 12891 451344 13074 455420
rect 16510 451344 16891 455420
rect 12891 445420 16891 451344
rect 12891 441344 13074 445420
rect 16510 441344 16891 445420
rect -1858 413518 8184 413640
rect -1858 409122 -1736 413518
rect 1060 409122 7046 413518
rect 7922 409122 8184 413518
rect -1858 408850 8184 409122
rect -1858 408408 9184 408530
rect -1858 404012 -1736 408408
rect 1060 404012 8246 408408
rect 9122 404012 9184 408408
rect -1858 403920 9184 404012
rect -1858 403478 8184 403600
rect -1858 399082 -1736 403478
rect 1060 399082 7046 403478
rect 7922 399082 8184 403478
rect -1858 398810 8184 399082
rect 12891 243281 16891 441344
rect 12891 239205 13130 243281
rect 16566 239205 16891 243281
rect 12891 239000 16891 239205
rect 17391 231156 21391 785944
rect 608660 388061 612660 942282
rect 627036 880278 634246 880400
rect 627036 875882 627098 880278
rect 627974 875882 631328 880278
rect 634124 875882 634246 880278
rect 627036 875610 634246 875882
rect 625836 875168 634246 875290
rect 625836 870772 625898 875168
rect 626774 870772 631328 875168
rect 634124 870772 634246 875168
rect 625836 870669 634246 870772
rect 627036 870227 634246 870349
rect 627036 865831 627098 870227
rect 627974 865831 631328 870227
rect 634124 865831 634246 870227
rect 627036 865559 634246 865831
rect 608660 383985 608843 388061
rect 612279 383985 612660 388061
rect 608660 378061 612660 383985
rect 608660 373985 608843 378061
rect 612279 373985 612660 378061
rect 608660 243281 612660 373985
rect 608660 239205 608899 243281
rect 612335 239205 612660 243281
rect 608660 239000 612660 239205
rect 613460 790861 617460 791201
rect 613460 786785 613643 790861
rect 617079 786785 617460 790861
rect 613460 780861 617460 786785
rect 613460 776785 613643 780861
rect 617079 776785 617460 780861
rect 613460 476261 617460 776785
rect 613460 472185 613643 476261
rect 617079 472185 617460 476261
rect 613460 466261 617460 472185
rect 613460 462185 613643 466261
rect 617079 462185 617460 466261
rect 613460 243281 617460 462185
rect 625836 432478 634246 432600
rect 625836 428082 625898 432478
rect 626774 428082 631328 432478
rect 634124 428082 634246 432478
rect 625836 427810 634246 428082
rect 627036 427368 634246 427490
rect 627036 422972 627098 427368
rect 627974 422972 631328 427368
rect 634124 422972 634246 427368
rect 627036 422869 634246 422972
rect 625836 422427 634246 422549
rect 625836 418031 625898 422427
rect 626774 418031 631328 422427
rect 634124 418031 634246 422427
rect 625836 417759 634246 418031
rect 613460 239205 613699 243281
rect 617135 239205 617460 243281
rect 613460 239000 617460 239205
rect -1858 40718 3184 40840
rect -1858 36322 -1736 40718
rect 1060 36322 2246 40718
rect 3122 36322 3184 40718
rect -1858 36050 3184 36322
rect -1858 30678 3184 30800
rect -1858 26282 -1736 30678
rect 1060 26282 2246 30678
rect 3122 26282 3184 30678
rect -1858 26010 3184 26282
<< properties >>
string FIXED_BBOX 0 0 633000 953400
<< end >>
