VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO manual_power_connections
  CLASS BLOCK ;
  FOREIGN manual_power_connections ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.100 BY 0.100 ;
END manual_power_connections
END LIBRARY

